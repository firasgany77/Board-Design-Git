-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     May 24 2022 18:35:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : in std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : in std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__39256\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39246\ : std_logic;
signal \N__39245\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39229\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39227\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39218\ : std_logic;
signal \N__39211\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39202\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39200\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39191\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39182\ : std_logic;
signal \N__39175\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39173\ : std_logic;
signal \N__39166\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39164\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39155\ : std_logic;
signal \N__39148\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39139\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39130\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39121\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39112\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39103\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39101\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39092\ : std_logic;
signal \N__39085\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39083\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39074\ : std_logic;
signal \N__39067\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39065\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39056\ : std_logic;
signal \N__39049\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39038\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39021\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39003\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38993\ : std_logic;
signal \N__38986\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38977\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38975\ : std_logic;
signal \N__38968\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38966\ : std_logic;
signal \N__38959\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38950\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38948\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38939\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38930\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38921\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38896\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38887\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38876\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38841\ : std_logic;
signal \N__38840\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38831\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38813\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38797\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38795\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38786\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38777\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38769\ : std_logic;
signal \N__38768\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38752\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38711\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38702\ : std_logic;
signal \N__38701\ : std_logic;
signal \N__38698\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38692\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38636\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38628\ : std_logic;
signal \N__38625\ : std_logic;
signal \N__38624\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38615\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38611\ : std_logic;
signal \N__38610\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38595\ : std_logic;
signal \N__38594\ : std_logic;
signal \N__38591\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38589\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38585\ : std_logic;
signal \N__38582\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38578\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38575\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38564\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38549\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38522\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38514\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38506\ : std_logic;
signal \N__38503\ : std_logic;
signal \N__38500\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38488\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38477\ : std_logic;
signal \N__38474\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38453\ : std_logic;
signal \N__38450\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38441\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38423\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38421\ : std_logic;
signal \N__38420\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38412\ : std_logic;
signal \N__38409\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38396\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38386\ : std_logic;
signal \N__38383\ : std_logic;
signal \N__38380\ : std_logic;
signal \N__38377\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38371\ : std_logic;
signal \N__38368\ : std_logic;
signal \N__38367\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38355\ : std_logic;
signal \N__38354\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38345\ : std_logic;
signal \N__38342\ : std_logic;
signal \N__38341\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38314\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38309\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38299\ : std_logic;
signal \N__38296\ : std_logic;
signal \N__38293\ : std_logic;
signal \N__38290\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38267\ : std_logic;
signal \N__38264\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38262\ : std_logic;
signal \N__38261\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38232\ : std_logic;
signal \N__38229\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38210\ : std_logic;
signal \N__38207\ : std_logic;
signal \N__38206\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38195\ : std_logic;
signal \N__38192\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38186\ : std_logic;
signal \N__38183\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38173\ : std_logic;
signal \N__38170\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38155\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38149\ : std_logic;
signal \N__38146\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38123\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38117\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38075\ : std_logic;
signal \N__38072\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38020\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38008\ : std_logic;
signal \N__37999\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37955\ : std_logic;
signal \N__37952\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37913\ : std_logic;
signal \N__37910\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37883\ : std_logic;
signal \N__37882\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37862\ : std_logic;
signal \N__37855\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37813\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37796\ : std_logic;
signal \N__37793\ : std_logic;
signal \N__37790\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37777\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37775\ : std_logic;
signal \N__37774\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37772\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37769\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37763\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37760\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37734\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37697\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37677\ : std_logic;
signal \N__37674\ : std_logic;
signal \N__37671\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37563\ : std_logic;
signal \N__37562\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37532\ : std_logic;
signal \N__37529\ : std_logic;
signal \N__37526\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37484\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37480\ : std_logic;
signal \N__37477\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37475\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37462\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37438\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37408\ : std_logic;
signal \N__37405\ : std_logic;
signal \N__37400\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37385\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37367\ : std_logic;
signal \N__37364\ : std_logic;
signal \N__37361\ : std_logic;
signal \N__37358\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37340\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37316\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37304\ : std_logic;
signal \N__37301\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37283\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37271\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37265\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37250\ : std_logic;
signal \N__37247\ : std_logic;
signal \N__37244\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37158\ : std_logic;
signal \N__37155\ : std_logic;
signal \N__37152\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37088\ : std_logic;
signal \N__37087\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37076\ : std_logic;
signal \N__37075\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37069\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36986\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36976\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36966\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36899\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36890\ : std_logic;
signal \N__36889\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36879\ : std_logic;
signal \N__36878\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36876\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36867\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36863\ : std_logic;
signal \N__36860\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36854\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36842\ : std_logic;
signal \N__36833\ : std_logic;
signal \N__36830\ : std_logic;
signal \N__36827\ : std_logic;
signal \N__36824\ : std_logic;
signal \N__36821\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36815\ : std_logic;
signal \N__36812\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36799\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36751\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36746\ : std_logic;
signal \N__36743\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36739\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36729\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36698\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36569\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36553\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36528\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36501\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36495\ : std_logic;
signal \N__36492\ : std_logic;
signal \N__36489\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36476\ : std_logic;
signal \N__36475\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36458\ : std_logic;
signal \N__36455\ : std_logic;
signal \N__36452\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36443\ : std_logic;
signal \N__36440\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36434\ : std_logic;
signal \N__36429\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36419\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36383\ : std_logic;
signal \N__36380\ : std_logic;
signal \N__36377\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36300\ : std_logic;
signal \N__36297\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36285\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36282\ : std_logic;
signal \N__36275\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36267\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36263\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36248\ : std_logic;
signal \N__36245\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36239\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36212\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36203\ : std_logic;
signal \N__36202\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36193\ : std_logic;
signal \N__36190\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36180\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36157\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35999\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35890\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35879\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35873\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35864\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35791\ : std_logic;
signal \N__35788\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35720\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35709\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35693\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35676\ : std_logic;
signal \N__35673\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35666\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35624\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35609\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35601\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35579\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35501\ : std_logic;
signal \N__35498\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35469\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35466\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35456\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35429\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35373\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35309\ : std_logic;
signal \N__35306\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35253\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35222\ : std_logic;
signal \N__35219\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35201\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35193\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35187\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35138\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35081\ : std_logic;
signal \N__35078\ : std_logic;
signal \N__35075\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35066\ : std_logic;
signal \N__35063\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35052\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35013\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35010\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34972\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34966\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34958\ : std_logic;
signal \N__34957\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34929\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34870\ : std_logic;
signal \N__34867\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34859\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34781\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34775\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34766\ : std_logic;
signal \N__34763\ : std_logic;
signal \N__34760\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34733\ : std_logic;
signal \N__34730\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34706\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34691\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34688\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34684\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34643\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34619\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34603\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34559\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34440\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34429\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34419\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34349\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34338\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34298\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34271\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34253\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34206\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34134\ : std_logic;
signal \N__34131\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34090\ : std_logic;
signal \N__34087\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34070\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33831\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33764\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33732\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33626\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33560\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33554\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33500\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33471\ : std_logic;
signal \N__33468\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33389\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33382\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33380\ : std_logic;
signal \N__33379\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33374\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33311\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33161\ : std_logic;
signal \N__33154\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33020\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32945\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32929\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32816\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32768\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32694\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32679\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32607\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32594\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32571\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32531\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32501\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32495\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32474\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32459\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32454\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32414\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32335\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32282\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32261\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32221\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32116\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32048\ : std_logic;
signal \N__32047\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32024\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__32000\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31937\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31867\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31843\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31802\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31658\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31565\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31485\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31473\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31467\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31420\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31417\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31382\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31313\ : std_logic;
signal \N__31310\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31209\ : std_logic;
signal \N__31206\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31077\ : std_logic;
signal \N__31074\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31070\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31064\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31043\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31022\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30995\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30968\ : std_logic;
signal \N__30965\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30949\ : std_logic;
signal \N__30946\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30897\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30881\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30864\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30827\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30808\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30737\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30563\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30530\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30404\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30361\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30353\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30313\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30286\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30234\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30060\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30008\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29963\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29904\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29891\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29807\ : std_logic;
signal \N__29804\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29780\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29396\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29349\ : std_logic;
signal \N__29346\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29339\ : std_logic;
signal \N__29336\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29121\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29058\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28969\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28869\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28839\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28832\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28823\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28691\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28622\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28475\ : std_logic;
signal \N__28472\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28358\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28250\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28238\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28232\ : std_logic;
signal \N__28229\ : std_logic;
signal \N__28226\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27941\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27813\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27699\ : std_logic;
signal \N__27696\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27576\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27488\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27323\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27168\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27077\ : std_logic;
signal \N__27072\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27042\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26874\ : std_logic;
signal \N__26871\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26701\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26394\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26319\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26274\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26250\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26217\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26085\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26067\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26046\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26034\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25730\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25689\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25634\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25427\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25397\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25339\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25327\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25006\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24759\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24590\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24403\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24296\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24215\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24080\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23727\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23559\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22709\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22454\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22167\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22161\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21626\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20753\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20538\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19868\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18634\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18312\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18267\ : std_logic;
signal \N__18264\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17898\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15663\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.count_rst_6\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_6_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_14\ : std_logic;
signal \PCH_PWRGD.count_i_0_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_0\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_9_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_13\ : std_logic;
signal \PCH_PWRGD.count_i_0\ : std_logic;
signal \PCH_PWRGD.N_1_i_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_7\ : std_logic;
signal \PCH_PWRGD.count_rst_3\ : std_logic;
signal \PCH_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_4\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_14\ : std_logic;
signal \RSMRST_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_5_9\ : std_logic;
signal \RSMRST_PWRGD.count_rst_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_5_10\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_9\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_12\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_5\ : std_logic;
signal \RSMRST_PWRGD.count_5_14\ : std_logic;
signal \RSMRST_PWRGD.count_rst_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.count_rst_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_5_5\ : std_logic;
signal \RSMRST_PWRGD.count_rst_0\ : std_logic;
signal \RSMRST_PWRGD.count_5_11\ : std_logic;
signal \RSMRST_PWRGD.N_240_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.count_rst_1\ : std_logic;
signal \RSMRST_PWRGD.count_5_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_4\ : std_logic;
signal \RSMRST_PWRGD.count_5_15\ : std_logic;
signal \POWERLED.func_state_enZ0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_0\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \POWERLED.func_state_1_m2_0_cascade_\ : std_logic;
signal vccst_en : std_logic;
signal \POWERLED.un1_func_state25_6_0_a3_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \POWERLED.N_189_i_cascade_\ : std_logic;
signal \POWERLED.N_238\ : std_logic;
signal \POWERLED.N_189_i\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.dutycycle_eena_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_0\ : std_logic;
signal \POWERLED.N_120_f0_1\ : std_logic;
signal \POWERLED.dutycycle_eena_0\ : std_logic;
signal \POWERLED.dutycycle_eena_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_1\ : std_logic;
signal \POWERLED.g0_18_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_0\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \POWERLED.g2_1\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m0_0\ : std_logic;
signal \POWERLED.g2_0_0_1_0_cascade_\ : std_logic;
signal \POWERLED.N_237\ : std_logic;
signal \POWERLED.N_3297_0_0_0_cascade_\ : std_logic;
signal \POWERLED.g1_0_1_0_1\ : std_logic;
signal \POWERLED.N_3297_0_0_2\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m3_0_0_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_o2_0_0_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_164_0\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1_0_cascade_\ : std_logic;
signal \POWERLED.g0_0_m2_1\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1_1_0\ : std_logic;
signal \POWERLED.N_134\ : std_logic;
signal \POWERLED.un1_dutycycle_168_0_0_1\ : std_logic;
signal \POWERLED.g1_1_0\ : std_logic;
signal \POWERLED.g2_0_1_cascade_\ : std_logic;
signal \POWERLED.g0_10_0_0_1\ : std_logic;
signal \POWERLED.g2_0_cascade_\ : std_logic;
signal \POWERLED.g0_10_0_0_0\ : std_logic;
signal \POWERLED.g0_8_1\ : std_logic;
signal \POWERLED.g1_1_0_1_0\ : std_logic;
signal \POWERLED.un1_dutycycle_inv_4_0\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_5\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.count_rst_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_5_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.count_rst_11\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_0\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.count_rst_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \RSMRST_PWRGD.count_rst_8\ : std_logic;
signal \RSMRST_PWRGD.count_5_3\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.count_5_13\ : std_logic;
signal \RSMRST_PWRGD.count_rst_2_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_13_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_5_8\ : std_logic;
signal \RSMRST_PWRGD.count_rst_11\ : std_logic;
signal \RSMRST_PWRGD.count_5_6\ : std_logic;
signal \RSMRST_PWRGD.count_5_7\ : std_logic;
signal \RSMRST_PWRGD.count_rst_12\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_4_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_rst_9\ : std_logic;
signal \RSMRST_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_1\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.count_5_2\ : std_logic;
signal \RSMRST_PWRGD.count_rst_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_3\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_4\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \RSMRST_PWRGD.count_5_4\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_1_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_4\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_5\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_11_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_12\ : std_logic;
signal \RSMRST_PWRGD.count_5_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \RSMRST_PWRGD.count_rst_6\ : std_logic;
signal \RSMRST_PWRGD.count_5_1\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\ : std_logic;
signal \RSMRST_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un12_clk_100khz_2\ : std_logic;
signal \POWERLED.func_state_RNIAE974Z0Z_0\ : std_logic;
signal \POWERLED.func_state_1_m2_am_1_1_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_1_cascade_\ : std_logic;
signal \POWERLED.N_79\ : std_logic;
signal \POWERLED.func_state_RNIQTLM2Z0Z_1\ : std_logic;
signal \POWERLED.N_79_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_1\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.func_state_enZ0\ : std_logic;
signal \POWERLED.func_state_1_m2_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_set_0_0\ : std_logic;
signal \POWERLED.dutycycle_set_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.N_346_cascade_\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIQBTF3_0Z0Z_1\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o2_1\ : std_logic;
signal \POWERLED.func_state_RNIQBTF3_1Z0Z_1\ : std_logic;
signal \POWERLED.N_343\ : std_logic;
signal \POWERLED.N_118_f0\ : std_logic;
signal \POWERLED.dutycycle_eena_3_0_0_sx_cascade_\ : std_logic;
signal \POWERLED.N_393\ : std_logic;
signal \POWERLED.func_state_0_sqmuxa_0_oZ0Z2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI0DTG7Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_0_2\ : std_logic;
signal \POWERLED.dutycycle_RNIHGUM6Z0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\ : std_logic;
signal \POWERLED.N_301\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_a2_0_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_2\ : std_logic;
signal \POWERLED.dutycycle_set_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_set_1\ : std_logic;
signal \POWERLED.dutycycle_eena_14_0_0_1\ : std_logic;
signal \POWERLED.dutycycle_0_5\ : std_logic;
signal \POWERLED.dutycycle_er_RNIT8CS1Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_i3_mux\ : std_logic;
signal \POWERLED.N_235_N_cascade_\ : std_logic;
signal \POWERLED.N_434_N\ : std_logic;
signal \POWERLED.N_235_N\ : std_logic;
signal \POWERLED.un1_clk_100khz_42_and_i_a2_3_0\ : std_logic;
signal \POWERLED.N_371\ : std_logic;
signal \POWERLED.N_371_cascade_\ : std_logic;
signal \POWERLED.N_372_cascade_\ : std_logic;
signal \POWERLED.un1_m5_2_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_30_0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_30_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_a0_2_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_11Z0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_34_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_34_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_36_0\ : std_logic;
signal \POWERLED.un1_m2_0_a0_0_cascade_\ : std_logic;
signal \POWERLED.un1_m2_0_a0_1\ : std_logic;
signal \PCH_PWRGD.N_3120_i_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_7_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_1_0\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.curr_state_7_1_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.N_3122_i\ : std_logic;
signal \PCH_PWRGD.N_3120_i\ : std_logic;
signal \PCH_PWRGD.N_413\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_413_cascade_\ : std_logic;
signal \PCH_PWRGD.N_277_0\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0\ : std_logic;
signal \PCH_PWRGD.N_277_0_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0_cascade_\ : std_logic;
signal \PCH_PWRGD.un12_clk_100khz_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.N_278_0\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \RSMRST_PWRGD.N_423_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \curr_state_RNIR5QD1_0_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_state_1_1\ : std_logic;
signal \RSMRST_PWRGD.curr_state_2_0\ : std_logic;
signal \RSMRST_PWRGD.m4_0_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_423\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_state_7_1\ : std_logic;
signal \POWERLED.count_off_1_0_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.count_off_0_3\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \POWERLED.func_state_RNI3IN21_2Z0Z_1\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\ : std_logic;
signal \POWERLED.N_425_cascade_\ : std_logic;
signal \POWERLED.N_175_cascade_\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_bm_1\ : std_logic;
signal \POWERLED.count_clk_en_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_en_2\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_0_o3_out\ : std_logic;
signal \POWERLED.un1_clk_100khz_2_i_o3_0\ : std_logic;
signal \POWERLED.func_state_RNI3IN21_1Z0Z_1_cascade_\ : std_logic;
signal \clk_100Khz_signalkeep_4_rep1\ : std_logic;
signal \POWERLED.func_state_0_sqmuxa_0_o2_xZ0\ : std_logic;
signal \POWERLED.N_233_N\ : std_logic;
signal \curr_state_RNIR5QD1_0_0\ : std_logic;
signal \clk_100Khz_signalkeep_4_fast\ : std_logic;
signal \RSMRST_PWRGD_RSMRSTn_fast\ : std_logic;
signal \rsmrstn_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_42_and_i_o2_1_1_cascade_\ : std_logic;
signal \POWERLED.N_171\ : std_logic;
signal \POWERLED.N_171_cascade_\ : std_logic;
signal \POWERLED.N_387\ : std_logic;
signal \POWERLED.dutycycle_m1_0_a2_0_cascade_\ : std_logic;
signal \POWERLED.N_145_N\ : std_logic;
signal \POWERLED.g1Z0Z_3\ : std_logic;
signal \POWERLED.g2_2\ : std_logic;
signal \POWERLED.func_state_1_m2_am_1_0\ : std_logic;
signal slp_s4n : std_logic;
signal slp_s3n : std_logic;
signal \POWERLED.un1_clk_100khz_42_and_i_o2_1_1\ : std_logic;
signal \POWERLED.func_state_RNI8H551Z0Z_0_cascade_\ : std_logic;
signal rsmrstn : std_logic;
signal \POWERLED.N_143_N_cascade_\ : std_logic;
signal \POWERLED.N_116_f0\ : std_logic;
signal \POWERLED.N_116_f0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_erZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_en_2\ : std_logic;
signal \POWERLED.N_3168_i\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_a0_1_a1_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_a0_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_13_1_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_a0_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_12\ : std_logic;
signal \POWERLED.func_state_RNI8H551Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNIANIR7Z0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIANIR7Z0Z_10\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \POWERLED.dutycycle_eena_3_d_0\ : std_logic;
signal \POWERLED.dutycycle_eena_3_0_0\ : std_logic;
signal \POWERLED.dutycycle_RNIANIR7Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIANIR7Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_10Z0Z_3\ : std_logic;
signal \POWERLED.func_state_RNI8H551_0Z0Z_0\ : std_logic;
signal \POWERLED.N_372\ : std_logic;
signal \POWERLED.func_state_RNIZ0Z_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_a2_6_0_0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_39_c_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_10_cascade_\ : std_logic;
signal v1p8a_ok : std_logic;
signal v5a_ok : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \N_392_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRSTn_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13_cascade_\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_2\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \HDA_STRAP.i4_mux_cascade_\ : std_logic;
signal \HDA_STRAP.curr_state_i_2_cascade_\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \HDA_STRAP.curr_state_3_1\ : std_logic;
signal \HDA_STRAP.N_208\ : std_logic;
signal \HDA_STRAP.curr_state_i_2\ : std_logic;
signal \HDA_STRAP.HDA_SDO_ATP_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.count_offZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_9_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.un34_clk_100khz_8\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_1_5\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.count_off_0_2\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \POWERLED.count_clk_0_10\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal \RSMRST_PWRGD.count_RNI166B31Z0Z_12\ : std_logic;
signal \RSMRST_PWRGD.count_0_sqmuxa\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.count_rst_5\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.N_388_N\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_1\ : std_logic;
signal \POWERLED.un1_func_state25_4_i_a2_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_1_1\ : std_logic;
signal \POWERLED.N_425\ : std_logic;
signal \POWERLED.count_clk_RNI0TA81Z0Z_7\ : std_logic;
signal \POWERLED.count_clk_RNI0TA81Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.N_128\ : std_logic;
signal \POWERLED.N_431_cascade_\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_0\ : std_logic;
signal \POWERLED.N_321\ : std_logic;
signal \POWERLED.un1_clk_100khz_43_and_i_0_d_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_40_and_i_0_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.dutycycle_en_8_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_40_and_i_0_0_0\ : std_logic;
signal \POWERLED.un1_clk_100khz_40_and_i_0_d_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_6\ : std_logic;
signal \POWERLED.dutycycle_en_6_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNIZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_cZ0\ : std_logic;
signal \POWERLED.N_308\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_7_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_44_d_c_1_s_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_2_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_44_d_1_0_tz\ : std_logic;
signal \POWERLED.dutycycle_er_RNIZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.N_297_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_ok_cascade_\ : std_logic;
signal vccst_pwrgd : std_logic;
signal pch_pwrok : std_logic;
signal \VPP_VDDQ.count_2_0_6\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_0\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11_cascade_\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_1\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \POWERLED.count_off_0_9\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_11\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_off_1_10\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.count_off_0_11\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \POWERLED.count_off_1_12\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.count_off_1_13\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_off_1_14\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNIPVUTZ0Z2\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.un34_clk_100khz_10\ : std_logic;
signal \POWERLED.count_off_0_6\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_12\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.un1_N_1_i\ : std_logic;
signal \POWERLED.g3_0_3_0_0\ : std_logic;
signal \POWERLED.N_164\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_1_0\ : std_logic;
signal \POWERLED.N_228\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\ : std_logic;
signal \POWERLED.func_state\ : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_1\ : std_logic;
signal \POWERLED.dutycycle_eena_5_d_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0\ : std_logic;
signal \POWERLED.dutycycle_RNIB8FGCZ0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNIB8FGCZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.N_158_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_11\ : std_logic;
signal \POWERLED.dutycycle_en_11_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HHZ0Z1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_11\ : std_logic;
signal \POWERLED.dutycycle_eena_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.dutycycle_eena_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_i1_mux\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_11_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_12_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.N_156_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_10\ : std_logic;
signal \POWERLED.dutycycle_en_10_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_13\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.N_143_N\ : std_logic;
signal \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\ : std_logic;
signal \POWERLED.N_161_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_en_12\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\ : std_logic;
signal \POWERLED.func_state_RNI3IN21_1Z0Z_1\ : std_logic;
signal \POWERLED.dutycycle_en_12_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.N_229_iZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_49_0_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_49_0_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_9_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_1_0_tz\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_13_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.count_2_0_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_rst_8_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_rst_7_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.count_2_rst_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2_rst_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.count_2_rst_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_10\ : std_logic;
signal \VPP_VDDQ.count_2_rst_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_12\ : std_logic;
signal \VPP_VDDQ.count_2_rst_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_14\ : std_logic;
signal \VPP_VDDQ.count_2_rst_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \PCH_PWRGD.N_424\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \POWERLED.count_0_5\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.count_0_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_15_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.N_193\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.N_178\ : std_logic;
signal \POWERLED.count_clkZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.N_385\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_1\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.count_clk_1_9\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.func_state_RNI43L44_0_0\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal \POWERLED.count_clk_en\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_6\ : std_logic;
signal \POWERLED.N_175\ : std_logic;
signal \POWERLED.N_175_i\ : std_logic;
signal \POWERLED.N_428\ : std_logic;
signal \POWERLED.func_state_RNI_5Z0Z_0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3_cZ0\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_11\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_11\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_15\ : std_logic;
signal \POWERLED.un1_dutycycle_53_44_d_1_a0_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.N_361\ : std_logic;
signal \POWERLED.dutycycle_er_RNIZ0Z_9\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_a2_1_4_cascade_\ : std_logic;
signal \POWERLED.N_369\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.un1_m2_2_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_rst_6\ : std_logic;
signal \VPP_VDDQ.count_2_rst_6_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.count_2_rst_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\ : std_logic;
signal \VPP_VDDQ.count_2_rst_3_cascade_\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_12\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_11\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_5_cascade_\ : std_logic;
signal \VPP_VDDQ.un29_clk_100khz_4\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\ : std_logic;
signal \VPP_VDDQ.N_1_i_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_sqmuxa\ : std_logic;
signal \VPP_VDDQ.count_2_rst_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.count_2_rst_3\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_5\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \HDA_STRAP.N_51\ : std_logic;
signal \HDA_STRAP.N_53\ : std_logic;
signal \HDA_STRAP.count_enZ0\ : std_logic;
signal \HDA_STRAP.N_3252_i\ : std_logic;
signal \N_414_cascade_\ : std_logic;
signal \HDA_STRAP.N_285\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \N_227\ : std_logic;
signal \HDA_STRAP.m6_i_0\ : std_logic;
signal \HDA_STRAP.m6_i_0_cascade_\ : std_logic;
signal \N_414\ : std_logic;
signal \HDA_STRAP.curr_state_4_0\ : std_logic;
signal \POWERLED.un79_clk_100khzlt6_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_3\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8_cascade_\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.count_1_3\ : std_logic;
signal \POWERLED.un1_count_cry_2\ : std_logic;
signal \POWERLED.un1_count_cry_3\ : std_logic;
signal \POWERLED.count_1_5\ : std_logic;
signal \POWERLED.un1_count_cry_4\ : std_logic;
signal \POWERLED.count_1_6\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.count_1_7\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.count_1_8\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \POWERLED.count_1_9\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.count_1_11\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.count_1_12\ : std_logic;
signal \POWERLED.un1_count_cry_11\ : std_logic;
signal \POWERLED.count_1_13\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.count_1_14\ : std_logic;
signal \POWERLED.un1_count_cry_13\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5\ : std_logic;
signal \DSW_PWRGD.curr_state_7_1_cascade_\ : std_logic;
signal \DSW_PWRGD.curr_state_2_1\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \DSW_PWRGD.curr_state_3_0\ : std_logic;
signal \DSW_PWRGD.curr_state_7_0_cascade_\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \bfn_8_9_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2_c\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_c\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_c\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_c\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_c\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.count_off_0_7\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.count_off_1_8\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \POWERLED.dutycycle_RNIBADV5Z0Z_0\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_4_sf\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un47_sum_s_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3_1_0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.un1_i3_mux_cascade_\ : std_logic;
signal \POWERLED.d_i3_mux\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_3140_i_cascade_\ : std_logic;
signal \VPP_VDDQ.m4_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.N_3140_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal vddq_ok : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_1\ : std_logic;
signal \DSW_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_5_cascade_\ : std_logic;
signal \DSW_PWRGD.count_rst_9\ : std_logic;
signal \DSW_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \DSW_PWRGD.count_1_5\ : std_logic;
signal \DSW_PWRGD.count_rst_4_cascade_\ : std_logic;
signal \VPP_VDDQ.N_3160_i\ : std_logic;
signal \DSW_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_6_cascade_\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_5\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \DSW_PWRGD.count_rst_6\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_8_cascade_\ : std_logic;
signal \DSW_PWRGD.count_1_8\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_13\ : std_logic;
signal \DSW_PWRGD.N_1_i_cascade_\ : std_logic;
signal \DSW_PWRGD.count_1_10\ : std_logic;
signal \POWERLED.g0_i_o3_0_cascade_\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \POWERLED.N_8\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal \POWERLED.g0_i_o3_0\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.curr_state_3_0_cascade_\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \POWERLED.count_1_0_cascade_\ : std_logic;
signal \POWERLED.count_1_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_0_1\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal \POWERLED.count_1_10\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal \POWERLED.count_1_2\ : std_logic;
signal \POWERLED.count_0_2\ : std_logic;
signal \DSW_PWRGD.count_1_6\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.count_rst_0\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \POWERLED.count_0_4\ : std_logic;
signal \POWERLED.count_1_4\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.un1_count_cry_0_i\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.N_6478_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.N_6479_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.N_6480_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.N_6481_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.N_6482_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.N_6483_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.un85_clk_100khz_7\ : std_logic;
signal \POWERLED.N_6484_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.un85_clk_100khz_8\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.N_6485_i\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_8\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.N_6486_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.N_6487_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.N_6488_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.N_6489_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.N_6490_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.N_6491_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_6492_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_8\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un47_sum\ : std_logic;
signal \POWERLED.mult1_un47_sum_i\ : std_logic;
signal v33a_ok : std_logic;
signal slp_susn : std_logic;
signal v1p8a_en : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_3119\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_0\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_4\ : std_logic;
signal \DSW_PWRGD.count_rst_12\ : std_logic;
signal \DSW_PWRGD.count_rst_12_cascade_\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_2_cascade_\ : std_logic;
signal \DSW_PWRGD.count_1_2\ : std_logic;
signal \DSW_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_3_cascade_\ : std_logic;
signal \DSW_PWRGD.count_1_3\ : std_logic;
signal \DSW_PWRGD.count_1_7\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_0\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_1_THRU_CO\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \DSW_PWRGD.countZ0Z_3\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_5\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \DSW_PWRGD.count_rst_8\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \DSW_PWRGD.countZ0Z_7\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_8\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \DSW_PWRGD.countZ0Z_10\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_10_cascade_\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_i_cascade_\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_8\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_9\ : std_logic;
signal \VPP_VDDQ.count_4_0\ : std_logic;
signal \VPP_VDDQ.count_rst_5_cascade_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_4_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_rst_6\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.curr_state_0_0\ : std_logic;
signal \VPP_VDDQ.count_2_rst_9\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.count_4_14\ : std_logic;
signal \VPP_VDDQ.count_4_5\ : std_logic;
signal \VPP_VDDQ.count_4_15\ : std_logic;
signal \VPP_VDDQ.count_4_6\ : std_logic;
signal \DSW_PWRGD.DSW_PWROK_0\ : std_logic;
signal dsw_pwrok : std_logic;
signal v5s_ok : std_logic;
signal \dsw_pwrok_cascade_\ : std_logic;
signal vccin_en : std_logic;
signal \VPP_VDDQ_delayed_vddq_pwrgd_en\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal v33dsw_ok : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \DSW_PWRGD.curr_state_RNI3E27Z0Z_0\ : std_logic;
signal v33s_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal v5s_enn : std_logic;
signal \N_392\ : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_3\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_0_1\ : std_logic;
signal \clk_100Khz_signalkeep_4\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_0\ : std_logic;
signal \VPP_VDDQ.count_4_10\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.N_188\ : std_logic;
signal \POWERLED.N_388\ : std_logic;
signal \POWERLED.un85_clk_100khz_6\ : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.m4_0_a2\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un85_clk_100khz_5\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_1\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_2\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \HDA_STRAP.count_3_14\ : std_logic;
signal \HDA_STRAP.count_3_4\ : std_logic;
signal \HDA_STRAP.count_3_7\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_5_cZ0\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_7\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_15\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_16\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \HDA_STRAP.count_0_17\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_15\ : std_logic;
signal \HDA_STRAP.count_1_6\ : std_logic;
signal \HDA_STRAP.count_3_6\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.count_3_15\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0\ : std_logic;
signal \HDA_STRAP.countZ0Z_6_cascade_\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_16\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.count_1_16\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_0\ : std_logic;
signal \DSW_PWRGD.count_rst_14\ : std_logic;
signal \DSW_PWRGD.count_rst_14_cascade_\ : std_logic;
signal \DSW_PWRGD.count_i_0_cascade_\ : std_logic;
signal \DSW_PWRGD.count_1_0\ : std_logic;
signal \DSW_PWRGD.count_rst_3_cascade_\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_11\ : std_logic;
signal \DSW_PWRGD.N_1_i\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_11_cascade_\ : std_logic;
signal \DSW_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \DSW_PWRGD.count_rst_3\ : std_logic;
signal \DSW_PWRGD.count_1_11\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_7\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_9\ : std_logic;
signal \DSW_PWRGD.count_1_12\ : std_logic;
signal \DSW_PWRGD.count_rst_2\ : std_logic;
signal \DSW_PWRGD.countZ0Z_12\ : std_logic;
signal \DSW_PWRGD.count_rst_5\ : std_logic;
signal \DSW_PWRGD.count_1_9\ : std_logic;
signal \DSW_PWRGD.countZ0Z_12_cascade_\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_1\ : std_logic;
signal \DSW_PWRGD.un2_count_1_axb_4\ : std_logic;
signal \DSW_PWRGD.count_rst_10\ : std_logic;
signal \DSW_PWRGD.count_1_4\ : std_logic;
signal \DSW_PWRGD.countZ0Z_6\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_0\ : std_logic;
signal \DSW_PWRGD.count_rst_1\ : std_logic;
signal \DSW_PWRGD.count_1_13\ : std_logic;
signal \DSW_PWRGD.count_rst_0\ : std_logic;
signal \DSW_PWRGD.count_1_14\ : std_logic;
signal \DSW_PWRGD.count_0_sqmuxa\ : std_logic;
signal \DSW_PWRGD.count_rst\ : std_logic;
signal \DSW_PWRGD.count_1_15\ : std_logic;
signal \DSW_PWRGD.countZ0Z_15\ : std_logic;
signal \DSW_PWRGD.count_i_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_14\ : std_logic;
signal \DSW_PWRGD.countZ0Z_15_cascade_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_13\ : std_logic;
signal \DSW_PWRGD.un12_clk_100khz_9\ : std_logic;
signal \DSW_PWRGD.count_1_1\ : std_logic;
signal \DSW_PWRGD.curr_state_RNI57NNZ0Z_0\ : std_logic;
signal \DSW_PWRGD.count_rst_13\ : std_logic;
signal \DSW_PWRGD.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_4_7\ : std_logic;
signal \VPP_VDDQ.count_4_8\ : std_logic;
signal \VPP_VDDQ.count_4_9\ : std_logic;
signal \VPP_VDDQ.count_4_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_2_cZ0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.count_rst_10\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.count_rst_11\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.count_rst_12\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.count_rst_13\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.count_rst_14\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \VPP_VDDQ.count_rst\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_i\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.count_rst_0\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.count_rst_3\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0\ : std_logic;
signal \VPP_VDDQ.count_rst_2\ : std_logic;
signal \VPP_VDDQ.count_4_13\ : std_logic;
signal \VPP_VDDQ.count_rst_1\ : std_logic;
signal \VPP_VDDQ.count_4_12\ : std_logic;
signal \VPP_VDDQ.count_rst_8\ : std_logic;
signal \VPP_VDDQ.count_4_3\ : std_logic;
signal \VPP_VDDQ.count_rst_9\ : std_logic;
signal \VPP_VDDQ.count_4_4\ : std_logic;
signal \POWERLED.func_state_RNI_1Z0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI2MQDZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_5\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_0_0\ : std_logic;
signal \VCCST_EN_i_0_o3_0\ : std_logic;
signal vpp_en : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ.N_194\ : std_logic;
signal \VPP_VDDQ.curr_state_0_0\ : std_logic;
signal \VPP_VDDQ.un4_count_1_axb_2\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_pwrgd_en_g\ : std_logic;
signal \VPP_VDDQ.count_en\ : std_logic;
signal \VPP_VDDQ.count_4_2\ : std_logic;
signal \VPP_VDDQ.count_en_cascade_\ : std_logic;
signal \VPP_VDDQ.count_rst_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2_cascade_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.un13_clk_100khz_11\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un145_sum\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un85_clk_100khz_3\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.N_203_i\ : std_logic;
signal \POWERLED.g0_9_0\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.count_3_3\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_2_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_5\ : std_logic;
signal \HDA_STRAP.count_3_13\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_3\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_9\ : std_logic;
signal \HDA_STRAP.count_3_12\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.count_3_9\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84\ : std_logic;
signal \HDA_STRAP.countZ0Z_12_cascade_\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_4\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_5\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\ : std_logic;
signal \HDA_STRAP.count_3_5\ : std_logic;
signal \HDA_STRAP.count_3_10\ : std_logic;
signal \HDA_STRAP.count_1_10\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_1_cascade_\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_1\ : std_logic;
signal \HDA_STRAP.count_RNIZ0Z_1\ : std_logic;
signal \HDA_STRAP.count_3_1\ : std_logic;
signal \HDA_STRAP.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614\ : std_logic;
signal \HDA_STRAP.count_3_2\ : std_logic;
signal \HDA_STRAP.count_1_11\ : std_logic;
signal \HDA_STRAP.count_3_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_0\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_6\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_14\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_7_cascade_\ : std_logic;
signal \HDA_STRAP.un25_clk_100khz_13\ : std_logic;
signal \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_\ : std_logic;
signal \HDA_STRAP.count_1_0_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_0_cascade_\ : std_logic;
signal \HDA_STRAP.count_RNI6OA47Z0Z_8\ : std_logic;
signal \HDA_STRAP.count_3_0\ : std_logic;
signal fpga_osc : std_logic;
signal \HDA_STRAP.count_1_8\ : std_logic;
signal \HDA_STRAP.count_3_8\ : std_logic;
signal \HDA_STRAP.count_en_g\ : std_logic;
signal \HDA_STRAP.un2_count_1_axb_8\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    \SUSWARN_N_wire\ <= SUSWARN_N;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    \VCCINAUX_VR_PE_wire\ <= VCCINAUX_VR_PE;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    \VCCIN_VR_PE_wire\ <= VCCIN_VR_PE;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39256\,
            DIN => \N__39255\,
            DOUT => \N__39254\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39256\,
            PADOUT => \N__39255\,
            PADIN => \N__39254\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39247\,
            DIN => \N__39246\,
            DOUT => \N__39245\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39247\,
            PADOUT => \N__39246\,
            PADIN => \N__39245\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39238\,
            DIN => \N__39237\,
            DOUT => \N__39236\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39238\,
            PADOUT => \N__39237\,
            PADIN => \N__39236\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30897\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39229\,
            DIN => \N__39228\,
            DOUT => \N__39227\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39229\,
            PADOUT => \N__39228\,
            PADIN => \N__39227\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16206\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39220\,
            DIN => \N__39219\,
            DOUT => \N__39218\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39220\,
            PADOUT => \N__39219\,
            PADIN => \N__39218\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39211\,
            DIN => \N__39210\,
            DOUT => \N__39209\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39211\,
            PADOUT => \N__39210\,
            PADIN => \N__39209\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39202\,
            DIN => \N__39201\,
            DOUT => \N__39200\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39202\,
            PADOUT => \N__39201\,
            PADIN => \N__39200\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39193\,
            DIN => \N__39192\,
            DOUT => \N__39191\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39193\,
            PADOUT => \N__39192\,
            PADIN => \N__39191\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39184\,
            DIN => \N__39183\,
            DOUT => \N__39182\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39184\,
            PADOUT => \N__39183\,
            PADIN => \N__39182\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32296\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39175\,
            DIN => \N__39174\,
            DOUT => \N__39173\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39175\,
            PADOUT => \N__39174\,
            PADIN => \N__39173\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39166\,
            DIN => \N__39165\,
            DOUT => \N__39164\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39166\,
            PADOUT => \N__39165\,
            PADIN => \N__39164\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39157\,
            DIN => \N__39156\,
            DOUT => \N__39155\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39157\,
            PADOUT => \N__39156\,
            PADIN => \N__39155\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29493\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39148\,
            DIN => \N__39147\,
            DOUT => \N__39146\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39148\,
            PADOUT => \N__39147\,
            PADIN => \N__39146\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39139\,
            DIN => \N__39138\,
            DOUT => \N__39137\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39139\,
            PADOUT => \N__39138\,
            PADIN => \N__39137\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39130\,
            DIN => \N__39129\,
            DOUT => \N__39128\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39130\,
            PADOUT => \N__39129\,
            PADIN => \N__39128\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39121\,
            DIN => \N__39120\,
            DOUT => \N__39119\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39121\,
            PADOUT => \N__39120\,
            PADIN => \N__39119\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39112\,
            DIN => \N__39111\,
            DOUT => \N__39110\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39112\,
            PADOUT => \N__39111\,
            PADIN => \N__39110\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16095\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39103\,
            DIN => \N__39102\,
            DOUT => \N__39101\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39103\,
            PADOUT => \N__39102\,
            PADIN => \N__39101\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39094\,
            DIN => \N__39093\,
            DOUT => \N__39092\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39094\,
            PADOUT => \N__39093\,
            PADIN => \N__39092\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39085\,
            DIN => \N__39084\,
            DOUT => \N__39083\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39085\,
            PADOUT => \N__39084\,
            PADIN => \N__39083\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39076\,
            DIN => \N__39075\,
            DOUT => \N__39074\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39076\,
            PADOUT => \N__39075\,
            PADIN => \N__39074\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39067\,
            DIN => \N__39066\,
            DOUT => \N__39065\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39067\,
            PADOUT => \N__39066\,
            PADIN => \N__39065\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39058\,
            DIN => \N__39057\,
            DOUT => \N__39056\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39058\,
            PADOUT => \N__39057\,
            PADIN => \N__39056\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__39049\,
            DIN => \N__39048\,
            DOUT => \N__39047\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39049\,
            PADOUT => \N__39048\,
            PADIN => \N__39047\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39040\,
            DIN => \N__39039\,
            DOUT => \N__39038\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39040\,
            PADOUT => \N__39039\,
            PADIN => \N__39038\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18978\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39031\,
            DIN => \N__39030\,
            DOUT => \N__39029\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39031\,
            PADOUT => \N__39030\,
            PADIN => \N__39029\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39022\,
            DIN => \N__39021\,
            DOUT => \N__39020\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39022\,
            PADOUT => \N__39021\,
            PADIN => \N__39020\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21093\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39013\,
            DIN => \N__39012\,
            DOUT => \N__39011\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39013\,
            PADOUT => \N__39012\,
            PADIN => \N__39011\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21087\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__39004\,
            DIN => \N__39003\,
            DOUT => \N__39002\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__39004\,
            PADOUT => \N__39003\,
            PADIN => \N__39002\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38995\,
            DIN => \N__38994\,
            DOUT => \N__38993\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38995\,
            PADOUT => \N__38994\,
            PADIN => \N__38993\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38986\,
            DIN => \N__38985\,
            DOUT => \N__38984\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38986\,
            PADOUT => \N__38985\,
            PADIN => \N__38984\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38977\,
            DIN => \N__38976\,
            DOUT => \N__38975\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38977\,
            PADOUT => \N__38976\,
            PADIN => \N__38975\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38968\,
            DIN => \N__38967\,
            DOUT => \N__38966\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38968\,
            PADOUT => \N__38967\,
            PADIN => \N__38966\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38959\,
            DIN => \N__38958\,
            DOUT => \N__38957\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38959\,
            PADOUT => \N__38958\,
            PADIN => \N__38957\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19845\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38950\,
            DIN => \N__38949\,
            DOUT => \N__38948\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38950\,
            PADOUT => \N__38949\,
            PADIN => \N__38948\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38941\,
            DIN => \N__38940\,
            DOUT => \N__38939\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38941\,
            PADOUT => \N__38940\,
            PADIN => \N__38939\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__36138\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__38932\,
            DIN => \N__38931\,
            DOUT => \N__38930\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38932\,
            PADOUT => \N__38931\,
            PADIN => \N__38930\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38923\,
            DIN => \N__38922\,
            DOUT => \N__38921\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38923\,
            PADOUT => \N__38922\,
            PADIN => \N__38921\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38914\,
            DIN => \N__38913\,
            DOUT => \N__38912\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38914\,
            PADOUT => \N__38913\,
            PADIN => \N__38912\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38905\,
            DIN => \N__38904\,
            DOUT => \N__38903\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38905\,
            PADOUT => \N__38904\,
            PADIN => \N__38903\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38896\,
            DIN => \N__38895\,
            DOUT => \N__38894\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38896\,
            PADOUT => \N__38895\,
            PADIN => \N__38894\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19551\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38887\,
            DIN => \N__38886\,
            DOUT => \N__38885\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38887\,
            PADOUT => \N__38886\,
            PADIN => \N__38885\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38878\,
            DIN => \N__38877\,
            DOUT => \N__38876\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38878\,
            PADOUT => \N__38877\,
            PADIN => \N__38876\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32331\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38869\,
            DIN => \N__38868\,
            DOUT => \N__38867\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38869\,
            PADOUT => \N__38868\,
            PADIN => \N__38867\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38860\,
            DIN => \N__38859\,
            DOUT => \N__38858\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38860\,
            PADOUT => \N__38859\,
            PADIN => \N__38858\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32697\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38851\,
            DIN => \N__38850\,
            DOUT => \N__38849\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38851\,
            PADOUT => \N__38850\,
            PADIN => \N__38849\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30968\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38842\,
            DIN => \N__38841\,
            DOUT => \N__38840\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38842\,
            PADOUT => \N__38841\,
            PADIN => \N__38840\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38833\,
            DIN => \N__38832\,
            DOUT => \N__38831\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38833\,
            PADOUT => \N__38832\,
            PADIN => \N__38831\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__38824\,
            DIN => \N__38823\,
            DOUT => \N__38822\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38824\,
            PADOUT => \N__38823\,
            PADIN => \N__38822\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38815\,
            DIN => \N__38814\,
            DOUT => \N__38813\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38815\,
            PADOUT => \N__38814\,
            PADIN => \N__38813\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38806\,
            DIN => \N__38805\,
            DOUT => \N__38804\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38806\,
            PADOUT => \N__38805\,
            PADIN => \N__38804\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32664\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38797\,
            DIN => \N__38796\,
            DOUT => \N__38795\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38797\,
            PADOUT => \N__38796\,
            PADIN => \N__38795\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38788\,
            DIN => \N__38787\,
            DOUT => \N__38786\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38788\,
            PADOUT => \N__38787\,
            PADIN => \N__38786\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38779\,
            DIN => \N__38778\,
            DOUT => \N__38777\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38779\,
            PADOUT => \N__38778\,
            PADIN => \N__38777\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38770\,
            DIN => \N__38769\,
            DOUT => \N__38768\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38770\,
            PADOUT => \N__38769\,
            PADIN => \N__38768\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38761\,
            DIN => \N__38760\,
            DOUT => \N__38759\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38761\,
            PADOUT => \N__38760\,
            PADIN => \N__38759\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38752\,
            DIN => \N__38751\,
            DOUT => \N__38750\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38752\,
            PADOUT => \N__38751\,
            PADIN => \N__38750\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38743\,
            DIN => \N__38742\,
            DOUT => \N__38741\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38743\,
            PADOUT => \N__38742\,
            PADIN => \N__38741\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21080\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__38734\,
            DIN => \N__38733\,
            DOUT => \N__38732\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__38734\,
            PADOUT => \N__38733\,
            PADIN => \N__38732\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__8999\ : CascadeMux
    port map (
            O => \N__38715\,
            I => \HDA_STRAP.countZ0Z_0_cascade_\
        );

    \I__8998\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38703\
        );

    \I__8997\ : InMux
    port map (
            O => \N__38711\,
            I => \N__38703\
        );

    \I__8996\ : InMux
    port map (
            O => \N__38710\,
            I => \N__38703\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38698\
        );

    \I__8994\ : InMux
    port map (
            O => \N__38702\,
            I => \N__38693\
        );

    \I__8993\ : InMux
    port map (
            O => \N__38701\,
            I => \N__38693\
        );

    \I__8992\ : Span4Mux_s3_v
    port map (
            O => \N__38698\,
            I => \N__38687\
        );

    \I__8991\ : LocalMux
    port map (
            O => \N__38693\,
            I => \N__38682\
        );

    \I__8990\ : InMux
    port map (
            O => \N__38692\,
            I => \N__38679\
        );

    \I__8989\ : InMux
    port map (
            O => \N__38691\,
            I => \N__38674\
        );

    \I__8988\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38674\
        );

    \I__8987\ : Span4Mux_h
    port map (
            O => \N__38687\,
            I => \N__38671\
        );

    \I__8986\ : InMux
    port map (
            O => \N__38686\,
            I => \N__38668\
        );

    \I__8985\ : InMux
    port map (
            O => \N__38685\,
            I => \N__38665\
        );

    \I__8984\ : Span4Mux_h
    port map (
            O => \N__38682\,
            I => \N__38662\
        );

    \I__8983\ : LocalMux
    port map (
            O => \N__38679\,
            I => \N__38657\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__38674\,
            I => \N__38657\
        );

    \I__8981\ : Sp12to4
    port map (
            O => \N__38671\,
            I => \N__38654\
        );

    \I__8980\ : LocalMux
    port map (
            O => \N__38668\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__38665\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__38662\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__8977\ : Odrv4
    port map (
            O => \N__38657\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__8976\ : Odrv12
    port map (
            O => \N__38654\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8\
        );

    \I__8975\ : InMux
    port map (
            O => \N__38643\,
            I => \N__38640\
        );

    \I__8974\ : LocalMux
    port map (
            O => \N__38640\,
            I => \HDA_STRAP.count_3_0\
        );

    \I__8973\ : ClkMux
    port map (
            O => \N__38637\,
            I => \N__38631\
        );

    \I__8972\ : ClkMux
    port map (
            O => \N__38636\,
            I => \N__38628\
        );

    \I__8971\ : ClkMux
    port map (
            O => \N__38635\,
            I => \N__38625\
        );

    \I__8970\ : ClkMux
    port map (
            O => \N__38634\,
            I => \N__38615\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__38631\,
            I => \N__38607\
        );

    \I__8968\ : LocalMux
    port map (
            O => \N__38628\,
            I => \N__38602\
        );

    \I__8967\ : LocalMux
    port map (
            O => \N__38625\,
            I => \N__38602\
        );

    \I__8966\ : ClkMux
    port map (
            O => \N__38624\,
            I => \N__38599\
        );

    \I__8965\ : ClkMux
    port map (
            O => \N__38623\,
            I => \N__38596\
        );

    \I__8964\ : ClkMux
    port map (
            O => \N__38622\,
            I => \N__38591\
        );

    \I__8963\ : ClkMux
    port map (
            O => \N__38621\,
            I => \N__38585\
        );

    \I__8962\ : ClkMux
    port map (
            O => \N__38620\,
            I => \N__38582\
        );

    \I__8961\ : ClkMux
    port map (
            O => \N__38619\,
            I => \N__38578\
        );

    \I__8960\ : ClkMux
    port map (
            O => \N__38618\,
            I => \N__38571\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__38615\,
            I => \N__38568\
        );

    \I__8958\ : ClkMux
    port map (
            O => \N__38614\,
            I => \N__38565\
        );

    \I__8957\ : ClkMux
    port map (
            O => \N__38613\,
            I => \N__38561\
        );

    \I__8956\ : ClkMux
    port map (
            O => \N__38612\,
            I => \N__38558\
        );

    \I__8955\ : ClkMux
    port map (
            O => \N__38611\,
            I => \N__38554\
        );

    \I__8954\ : ClkMux
    port map (
            O => \N__38610\,
            I => \N__38551\
        );

    \I__8953\ : Span4Mux_s2_v
    port map (
            O => \N__38607\,
            I => \N__38538\
        );

    \I__8952\ : Span4Mux_s2_v
    port map (
            O => \N__38602\,
            I => \N__38538\
        );

    \I__8951\ : LocalMux
    port map (
            O => \N__38599\,
            I => \N__38538\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__38596\,
            I => \N__38538\
        );

    \I__8949\ : ClkMux
    port map (
            O => \N__38595\,
            I => \N__38535\
        );

    \I__8948\ : ClkMux
    port map (
            O => \N__38594\,
            I => \N__38530\
        );

    \I__8947\ : LocalMux
    port map (
            O => \N__38591\,
            I => \N__38526\
        );

    \I__8946\ : ClkMux
    port map (
            O => \N__38590\,
            I => \N__38523\
        );

    \I__8945\ : ClkMux
    port map (
            O => \N__38589\,
            I => \N__38519\
        );

    \I__8944\ : ClkMux
    port map (
            O => \N__38588\,
            I => \N__38516\
        );

    \I__8943\ : LocalMux
    port map (
            O => \N__38585\,
            I => \N__38509\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__38582\,
            I => \N__38509\
        );

    \I__8941\ : ClkMux
    port map (
            O => \N__38581\,
            I => \N__38506\
        );

    \I__8940\ : LocalMux
    port map (
            O => \N__38578\,
            I => \N__38503\
        );

    \I__8939\ : ClkMux
    port map (
            O => \N__38577\,
            I => \N__38500\
        );

    \I__8938\ : ClkMux
    port map (
            O => \N__38576\,
            I => \N__38497\
        );

    \I__8937\ : ClkMux
    port map (
            O => \N__38575\,
            I => \N__38494\
        );

    \I__8936\ : ClkMux
    port map (
            O => \N__38574\,
            I => \N__38490\
        );

    \I__8935\ : LocalMux
    port map (
            O => \N__38571\,
            I => \N__38482\
        );

    \I__8934\ : Span4Mux_s2_h
    port map (
            O => \N__38568\,
            I => \N__38477\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__38565\,
            I => \N__38477\
        );

    \I__8932\ : ClkMux
    port map (
            O => \N__38564\,
            I => \N__38474\
        );

    \I__8931\ : LocalMux
    port map (
            O => \N__38561\,
            I => \N__38470\
        );

    \I__8930\ : LocalMux
    port map (
            O => \N__38558\,
            I => \N__38467\
        );

    \I__8929\ : ClkMux
    port map (
            O => \N__38557\,
            I => \N__38464\
        );

    \I__8928\ : LocalMux
    port map (
            O => \N__38554\,
            I => \N__38458\
        );

    \I__8927\ : LocalMux
    port map (
            O => \N__38551\,
            I => \N__38458\
        );

    \I__8926\ : ClkMux
    port map (
            O => \N__38550\,
            I => \N__38453\
        );

    \I__8925\ : ClkMux
    port map (
            O => \N__38549\,
            I => \N__38450\
        );

    \I__8924\ : ClkMux
    port map (
            O => \N__38548\,
            I => \N__38446\
        );

    \I__8923\ : ClkMux
    port map (
            O => \N__38547\,
            I => \N__38442\
        );

    \I__8922\ : Span4Mux_v
    port map (
            O => \N__38538\,
            I => \N__38436\
        );

    \I__8921\ : LocalMux
    port map (
            O => \N__38535\,
            I => \N__38436\
        );

    \I__8920\ : ClkMux
    port map (
            O => \N__38534\,
            I => \N__38433\
        );

    \I__8919\ : ClkMux
    port map (
            O => \N__38533\,
            I => \N__38429\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__38530\,
            I => \N__38426\
        );

    \I__8917\ : ClkMux
    port map (
            O => \N__38529\,
            I => \N__38423\
        );

    \I__8916\ : Span4Mux_s3_h
    port map (
            O => \N__38526\,
            I => \N__38414\
        );

    \I__8915\ : LocalMux
    port map (
            O => \N__38523\,
            I => \N__38414\
        );

    \I__8914\ : ClkMux
    port map (
            O => \N__38522\,
            I => \N__38409\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__38519\,
            I => \N__38406\
        );

    \I__8912\ : LocalMux
    port map (
            O => \N__38516\,
            I => \N__38403\
        );

    \I__8911\ : ClkMux
    port map (
            O => \N__38515\,
            I => \N__38400\
        );

    \I__8910\ : ClkMux
    port map (
            O => \N__38514\,
            I => \N__38397\
        );

    \I__8909\ : Span4Mux_v
    port map (
            O => \N__38509\,
            I => \N__38391\
        );

    \I__8908\ : LocalMux
    port map (
            O => \N__38506\,
            I => \N__38391\
        );

    \I__8907\ : Span4Mux_s3_v
    port map (
            O => \N__38503\,
            I => \N__38386\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__38500\,
            I => \N__38386\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__38497\,
            I => \N__38383\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__38494\,
            I => \N__38380\
        );

    \I__8903\ : ClkMux
    port map (
            O => \N__38493\,
            I => \N__38377\
        );

    \I__8902\ : LocalMux
    port map (
            O => \N__38490\,
            I => \N__38374\
        );

    \I__8901\ : ClkMux
    port map (
            O => \N__38489\,
            I => \N__38371\
        );

    \I__8900\ : ClkMux
    port map (
            O => \N__38488\,
            I => \N__38368\
        );

    \I__8899\ : ClkMux
    port map (
            O => \N__38487\,
            I => \N__38363\
        );

    \I__8898\ : ClkMux
    port map (
            O => \N__38486\,
            I => \N__38360\
        );

    \I__8897\ : ClkMux
    port map (
            O => \N__38485\,
            I => \N__38356\
        );

    \I__8896\ : Span4Mux_h
    port map (
            O => \N__38482\,
            I => \N__38345\
        );

    \I__8895\ : Span4Mux_h
    port map (
            O => \N__38477\,
            I => \N__38345\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__38474\,
            I => \N__38345\
        );

    \I__8893\ : ClkMux
    port map (
            O => \N__38473\,
            I => \N__38342\
        );

    \I__8892\ : Span4Mux_v
    port map (
            O => \N__38470\,
            I => \N__38335\
        );

    \I__8891\ : Span4Mux_v
    port map (
            O => \N__38467\,
            I => \N__38335\
        );

    \I__8890\ : LocalMux
    port map (
            O => \N__38464\,
            I => \N__38332\
        );

    \I__8889\ : ClkMux
    port map (
            O => \N__38463\,
            I => \N__38329\
        );

    \I__8888\ : Span4Mux_s2_v
    port map (
            O => \N__38458\,
            I => \N__38325\
        );

    \I__8887\ : ClkMux
    port map (
            O => \N__38457\,
            I => \N__38322\
        );

    \I__8886\ : ClkMux
    port map (
            O => \N__38456\,
            I => \N__38316\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__38453\,
            I => \N__38310\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__38450\,
            I => \N__38305\
        );

    \I__8883\ : ClkMux
    port map (
            O => \N__38449\,
            I => \N__38302\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__38446\,
            I => \N__38299\
        );

    \I__8881\ : ClkMux
    port map (
            O => \N__38445\,
            I => \N__38296\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__38442\,
            I => \N__38293\
        );

    \I__8879\ : ClkMux
    port map (
            O => \N__38441\,
            I => \N__38290\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__38436\,
            I => \N__38285\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__38433\,
            I => \N__38285\
        );

    \I__8876\ : ClkMux
    port map (
            O => \N__38432\,
            I => \N__38282\
        );

    \I__8875\ : LocalMux
    port map (
            O => \N__38429\,
            I => \N__38279\
        );

    \I__8874\ : Span4Mux_h
    port map (
            O => \N__38426\,
            I => \N__38276\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__38423\,
            I => \N__38273\
        );

    \I__8872\ : ClkMux
    port map (
            O => \N__38422\,
            I => \N__38270\
        );

    \I__8871\ : ClkMux
    port map (
            O => \N__38421\,
            I => \N__38267\
        );

    \I__8870\ : ClkMux
    port map (
            O => \N__38420\,
            I => \N__38264\
        );

    \I__8869\ : ClkMux
    port map (
            O => \N__38419\,
            I => \N__38257\
        );

    \I__8868\ : Span4Mux_h
    port map (
            O => \N__38414\,
            I => \N__38254\
        );

    \I__8867\ : ClkMux
    port map (
            O => \N__38413\,
            I => \N__38251\
        );

    \I__8866\ : ClkMux
    port map (
            O => \N__38412\,
            I => \N__38248\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__38409\,
            I => \N__38245\
        );

    \I__8864\ : Span4Mux_h
    port map (
            O => \N__38406\,
            I => \N__38238\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__38403\,
            I => \N__38238\
        );

    \I__8862\ : LocalMux
    port map (
            O => \N__38400\,
            I => \N__38238\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__38397\,
            I => \N__38235\
        );

    \I__8860\ : ClkMux
    port map (
            O => \N__38396\,
            I => \N__38232\
        );

    \I__8859\ : Span4Mux_v
    port map (
            O => \N__38391\,
            I => \N__38229\
        );

    \I__8858\ : Span4Mux_v
    port map (
            O => \N__38386\,
            I => \N__38220\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__38383\,
            I => \N__38220\
        );

    \I__8856\ : Span4Mux_h
    port map (
            O => \N__38380\,
            I => \N__38220\
        );

    \I__8855\ : LocalMux
    port map (
            O => \N__38377\,
            I => \N__38220\
        );

    \I__8854\ : Span4Mux_h
    port map (
            O => \N__38374\,
            I => \N__38213\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__38371\,
            I => \N__38213\
        );

    \I__8852\ : LocalMux
    port map (
            O => \N__38368\,
            I => \N__38213\
        );

    \I__8851\ : ClkMux
    port map (
            O => \N__38367\,
            I => \N__38210\
        );

    \I__8850\ : ClkMux
    port map (
            O => \N__38366\,
            I => \N__38207\
        );

    \I__8849\ : LocalMux
    port map (
            O => \N__38363\,
            I => \N__38201\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__38360\,
            I => \N__38201\
        );

    \I__8847\ : ClkMux
    port map (
            O => \N__38359\,
            I => \N__38198\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__38356\,
            I => \N__38195\
        );

    \I__8845\ : ClkMux
    port map (
            O => \N__38355\,
            I => \N__38192\
        );

    \I__8844\ : ClkMux
    port map (
            O => \N__38354\,
            I => \N__38189\
        );

    \I__8843\ : ClkMux
    port map (
            O => \N__38353\,
            I => \N__38186\
        );

    \I__8842\ : ClkMux
    port map (
            O => \N__38352\,
            I => \N__38183\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__38345\,
            I => \N__38179\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__38342\,
            I => \N__38176\
        );

    \I__8839\ : ClkMux
    port map (
            O => \N__38341\,
            I => \N__38173\
        );

    \I__8838\ : ClkMux
    port map (
            O => \N__38340\,
            I => \N__38170\
        );

    \I__8837\ : Span4Mux_v
    port map (
            O => \N__38335\,
            I => \N__38163\
        );

    \I__8836\ : Span4Mux_h
    port map (
            O => \N__38332\,
            I => \N__38163\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__38329\,
            I => \N__38163\
        );

    \I__8834\ : ClkMux
    port map (
            O => \N__38328\,
            I => \N__38160\
        );

    \I__8833\ : Span4Mux_h
    port map (
            O => \N__38325\,
            I => \N__38155\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__38322\,
            I => \N__38155\
        );

    \I__8831\ : ClkMux
    port map (
            O => \N__38321\,
            I => \N__38152\
        );

    \I__8830\ : ClkMux
    port map (
            O => \N__38320\,
            I => \N__38149\
        );

    \I__8829\ : ClkMux
    port map (
            O => \N__38319\,
            I => \N__38146\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__38316\,
            I => \N__38143\
        );

    \I__8827\ : ClkMux
    port map (
            O => \N__38315\,
            I => \N__38140\
        );

    \I__8826\ : ClkMux
    port map (
            O => \N__38314\,
            I => \N__38137\
        );

    \I__8825\ : ClkMux
    port map (
            O => \N__38313\,
            I => \N__38134\
        );

    \I__8824\ : Span4Mux_v
    port map (
            O => \N__38310\,
            I => \N__38130\
        );

    \I__8823\ : ClkMux
    port map (
            O => \N__38309\,
            I => \N__38127\
        );

    \I__8822\ : ClkMux
    port map (
            O => \N__38308\,
            I => \N__38124\
        );

    \I__8821\ : Span4Mux_s1_h
    port map (
            O => \N__38305\,
            I => \N__38117\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__38302\,
            I => \N__38117\
        );

    \I__8819\ : Span4Mux_v
    port map (
            O => \N__38299\,
            I => \N__38112\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__38296\,
            I => \N__38112\
        );

    \I__8817\ : Span4Mux_v
    port map (
            O => \N__38293\,
            I => \N__38107\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__38290\,
            I => \N__38107\
        );

    \I__8815\ : IoSpan4Mux
    port map (
            O => \N__38285\,
            I => \N__38104\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__38282\,
            I => \N__38101\
        );

    \I__8813\ : Span4Mux_v
    port map (
            O => \N__38279\,
            I => \N__38092\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__38276\,
            I => \N__38092\
        );

    \I__8811\ : Span4Mux_s2_h
    port map (
            O => \N__38273\,
            I => \N__38092\
        );

    \I__8810\ : LocalMux
    port map (
            O => \N__38270\,
            I => \N__38092\
        );

    \I__8809\ : LocalMux
    port map (
            O => \N__38267\,
            I => \N__38089\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__38264\,
            I => \N__38086\
        );

    \I__8807\ : ClkMux
    port map (
            O => \N__38263\,
            I => \N__38083\
        );

    \I__8806\ : ClkMux
    port map (
            O => \N__38262\,
            I => \N__38080\
        );

    \I__8805\ : ClkMux
    port map (
            O => \N__38261\,
            I => \N__38077\
        );

    \I__8804\ : ClkMux
    port map (
            O => \N__38260\,
            I => \N__38072\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__38257\,
            I => \N__38067\
        );

    \I__8802\ : Span4Mux_h
    port map (
            O => \N__38254\,
            I => \N__38067\
        );

    \I__8801\ : LocalMux
    port map (
            O => \N__38251\,
            I => \N__38064\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38061\
        );

    \I__8799\ : Span4Mux_v
    port map (
            O => \N__38245\,
            I => \N__38052\
        );

    \I__8798\ : Span4Mux_v
    port map (
            O => \N__38238\,
            I => \N__38052\
        );

    \I__8797\ : Span4Mux_h
    port map (
            O => \N__38235\,
            I => \N__38052\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__38232\,
            I => \N__38052\
        );

    \I__8795\ : Span4Mux_h
    port map (
            O => \N__38229\,
            I => \N__38043\
        );

    \I__8794\ : Span4Mux_v
    port map (
            O => \N__38220\,
            I => \N__38043\
        );

    \I__8793\ : Span4Mux_v
    port map (
            O => \N__38213\,
            I => \N__38043\
        );

    \I__8792\ : LocalMux
    port map (
            O => \N__38210\,
            I => \N__38043\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__38207\,
            I => \N__38040\
        );

    \I__8790\ : ClkMux
    port map (
            O => \N__38206\,
            I => \N__38037\
        );

    \I__8789\ : Span4Mux_v
    port map (
            O => \N__38201\,
            I => \N__38026\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__38198\,
            I => \N__38026\
        );

    \I__8787\ : Span4Mux_s3_h
    port map (
            O => \N__38195\,
            I => \N__38026\
        );

    \I__8786\ : LocalMux
    port map (
            O => \N__38192\,
            I => \N__38026\
        );

    \I__8785\ : LocalMux
    port map (
            O => \N__38189\,
            I => \N__38026\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__38186\,
            I => \N__38023\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__38183\,
            I => \N__38020\
        );

    \I__8782\ : ClkMux
    port map (
            O => \N__38182\,
            I => \N__38017\
        );

    \I__8781\ : Span4Mux_v
    port map (
            O => \N__38179\,
            I => \N__38008\
        );

    \I__8780\ : Span4Mux_h
    port map (
            O => \N__38176\,
            I => \N__38008\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__38173\,
            I => \N__38008\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__38170\,
            I => \N__38008\
        );

    \I__8777\ : Span4Mux_v
    port map (
            O => \N__38163\,
            I => \N__37999\
        );

    \I__8776\ : LocalMux
    port map (
            O => \N__38160\,
            I => \N__37999\
        );

    \I__8775\ : Span4Mux_h
    port map (
            O => \N__38155\,
            I => \N__37999\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__38152\,
            I => \N__37999\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__38149\,
            I => \N__37994\
        );

    \I__8772\ : LocalMux
    port map (
            O => \N__38146\,
            I => \N__37994\
        );

    \I__8771\ : Span4Mux_h
    port map (
            O => \N__38143\,
            I => \N__37985\
        );

    \I__8770\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__37985\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__38137\,
            I => \N__37985\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__38134\,
            I => \N__37985\
        );

    \I__8767\ : ClkMux
    port map (
            O => \N__38133\,
            I => \N__37982\
        );

    \I__8766\ : Span4Mux_h
    port map (
            O => \N__38130\,
            I => \N__37975\
        );

    \I__8765\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__37975\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__38124\,
            I => \N__37975\
        );

    \I__8763\ : ClkMux
    port map (
            O => \N__38123\,
            I => \N__37972\
        );

    \I__8762\ : ClkMux
    port map (
            O => \N__38122\,
            I => \N__37969\
        );

    \I__8761\ : Span4Mux_v
    port map (
            O => \N__38117\,
            I => \N__37965\
        );

    \I__8760\ : Span4Mux_v
    port map (
            O => \N__38112\,
            I => \N__37960\
        );

    \I__8759\ : Span4Mux_v
    port map (
            O => \N__38107\,
            I => \N__37960\
        );

    \I__8758\ : IoSpan4Mux
    port map (
            O => \N__38104\,
            I => \N__37955\
        );

    \I__8757\ : IoSpan4Mux
    port map (
            O => \N__38101\,
            I => \N__37955\
        );

    \I__8756\ : Span4Mux_v
    port map (
            O => \N__38092\,
            I => \N__37952\
        );

    \I__8755\ : Span4Mux_v
    port map (
            O => \N__38089\,
            I => \N__37941\
        );

    \I__8754\ : Span4Mux_v
    port map (
            O => \N__38086\,
            I => \N__37941\
        );

    \I__8753\ : LocalMux
    port map (
            O => \N__38083\,
            I => \N__37941\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__37941\
        );

    \I__8751\ : LocalMux
    port map (
            O => \N__38077\,
            I => \N__37941\
        );

    \I__8750\ : ClkMux
    port map (
            O => \N__38076\,
            I => \N__37938\
        );

    \I__8749\ : ClkMux
    port map (
            O => \N__38075\,
            I => \N__37935\
        );

    \I__8748\ : LocalMux
    port map (
            O => \N__38072\,
            I => \N__37932\
        );

    \I__8747\ : IoSpan4Mux
    port map (
            O => \N__38067\,
            I => \N__37929\
        );

    \I__8746\ : Span4Mux_v
    port map (
            O => \N__38064\,
            I => \N__37920\
        );

    \I__8745\ : Span4Mux_h
    port map (
            O => \N__38061\,
            I => \N__37920\
        );

    \I__8744\ : IoSpan4Mux
    port map (
            O => \N__38052\,
            I => \N__37920\
        );

    \I__8743\ : Span4Mux_v
    port map (
            O => \N__38043\,
            I => \N__37920\
        );

    \I__8742\ : Span4Mux_s3_h
    port map (
            O => \N__38040\,
            I => \N__37913\
        );

    \I__8741\ : LocalMux
    port map (
            O => \N__38037\,
            I => \N__37913\
        );

    \I__8740\ : Span4Mux_v
    port map (
            O => \N__38026\,
            I => \N__37913\
        );

    \I__8739\ : IoSpan4Mux
    port map (
            O => \N__38023\,
            I => \N__37910\
        );

    \I__8738\ : Span4Mux_v
    port map (
            O => \N__38020\,
            I => \N__37905\
        );

    \I__8737\ : LocalMux
    port map (
            O => \N__38017\,
            I => \N__37905\
        );

    \I__8736\ : Span4Mux_v
    port map (
            O => \N__38008\,
            I => \N__37894\
        );

    \I__8735\ : IoSpan4Mux
    port map (
            O => \N__37999\,
            I => \N__37894\
        );

    \I__8734\ : Span4Mux_h
    port map (
            O => \N__37994\,
            I => \N__37894\
        );

    \I__8733\ : Span4Mux_v
    port map (
            O => \N__37985\,
            I => \N__37894\
        );

    \I__8732\ : LocalMux
    port map (
            O => \N__37982\,
            I => \N__37894\
        );

    \I__8731\ : Span4Mux_v
    port map (
            O => \N__37975\,
            I => \N__37887\
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__37972\,
            I => \N__37887\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__37969\,
            I => \N__37887\
        );

    \I__8728\ : ClkMux
    port map (
            O => \N__37968\,
            I => \N__37884\
        );

    \I__8727\ : IoSpan4Mux
    port map (
            O => \N__37965\,
            I => \N__37874\
        );

    \I__8726\ : IoSpan4Mux
    port map (
            O => \N__37960\,
            I => \N__37874\
        );

    \I__8725\ : IoSpan4Mux
    port map (
            O => \N__37955\,
            I => \N__37874\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__37952\,
            I => \N__37869\
        );

    \I__8723\ : Span4Mux_v
    port map (
            O => \N__37941\,
            I => \N__37869\
        );

    \I__8722\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37862\
        );

    \I__8721\ : LocalMux
    port map (
            O => \N__37935\,
            I => \N__37862\
        );

    \I__8720\ : Sp12to4
    port map (
            O => \N__37932\,
            I => \N__37862\
        );

    \I__8719\ : IoSpan4Mux
    port map (
            O => \N__37929\,
            I => \N__37855\
        );

    \I__8718\ : IoSpan4Mux
    port map (
            O => \N__37920\,
            I => \N__37855\
        );

    \I__8717\ : IoSpan4Mux
    port map (
            O => \N__37913\,
            I => \N__37855\
        );

    \I__8716\ : IoSpan4Mux
    port map (
            O => \N__37910\,
            I => \N__37848\
        );

    \I__8715\ : IoSpan4Mux
    port map (
            O => \N__37905\,
            I => \N__37848\
        );

    \I__8714\ : IoSpan4Mux
    port map (
            O => \N__37894\,
            I => \N__37848\
        );

    \I__8713\ : Span4Mux_v
    port map (
            O => \N__37887\,
            I => \N__37843\
        );

    \I__8712\ : LocalMux
    port map (
            O => \N__37884\,
            I => \N__37843\
        );

    \I__8711\ : ClkMux
    port map (
            O => \N__37883\,
            I => \N__37840\
        );

    \I__8710\ : ClkMux
    port map (
            O => \N__37882\,
            I => \N__37837\
        );

    \I__8709\ : ClkMux
    port map (
            O => \N__37881\,
            I => \N__37834\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__37874\,
            I => fpga_osc
        );

    \I__8707\ : Odrv4
    port map (
            O => \N__37869\,
            I => fpga_osc
        );

    \I__8706\ : Odrv12
    port map (
            O => \N__37862\,
            I => fpga_osc
        );

    \I__8705\ : Odrv4
    port map (
            O => \N__37855\,
            I => fpga_osc
        );

    \I__8704\ : Odrv4
    port map (
            O => \N__37848\,
            I => fpga_osc
        );

    \I__8703\ : Odrv4
    port map (
            O => \N__37843\,
            I => fpga_osc
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__37840\,
            I => fpga_osc
        );

    \I__8701\ : LocalMux
    port map (
            O => \N__37837\,
            I => fpga_osc
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__37834\,
            I => fpga_osc
        );

    \I__8699\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37806\
        );

    \I__8698\ : InMux
    port map (
            O => \N__37814\,
            I => \N__37806\
        );

    \I__8697\ : InMux
    port map (
            O => \N__37813\,
            I => \N__37806\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__37806\,
            I => \N__37803\
        );

    \I__8695\ : Odrv4
    port map (
            O => \N__37803\,
            I => \HDA_STRAP.count_1_8\
        );

    \I__8694\ : CascadeMux
    port map (
            O => \N__37800\,
            I => \N__37797\
        );

    \I__8693\ : InMux
    port map (
            O => \N__37797\,
            I => \N__37793\
        );

    \I__8692\ : InMux
    port map (
            O => \N__37796\,
            I => \N__37790\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__37793\,
            I => \HDA_STRAP.count_3_8\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__37790\,
            I => \HDA_STRAP.count_3_8\
        );

    \I__8689\ : CascadeMux
    port map (
            O => \N__37785\,
            I => \N__37777\
        );

    \I__8688\ : InMux
    port map (
            O => \N__37784\,
            I => \N__37748\
        );

    \I__8687\ : InMux
    port map (
            O => \N__37783\,
            I => \N__37748\
        );

    \I__8686\ : InMux
    port map (
            O => \N__37782\,
            I => \N__37748\
        );

    \I__8685\ : InMux
    port map (
            O => \N__37781\,
            I => \N__37748\
        );

    \I__8684\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37745\
        );

    \I__8683\ : InMux
    port map (
            O => \N__37777\,
            I => \N__37734\
        );

    \I__8682\ : InMux
    port map (
            O => \N__37776\,
            I => \N__37734\
        );

    \I__8681\ : InMux
    port map (
            O => \N__37775\,
            I => \N__37734\
        );

    \I__8680\ : InMux
    port map (
            O => \N__37774\,
            I => \N__37734\
        );

    \I__8679\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37734\
        );

    \I__8678\ : InMux
    port map (
            O => \N__37772\,
            I => \N__37727\
        );

    \I__8677\ : InMux
    port map (
            O => \N__37771\,
            I => \N__37727\
        );

    \I__8676\ : InMux
    port map (
            O => \N__37770\,
            I => \N__37727\
        );

    \I__8675\ : InMux
    port map (
            O => \N__37769\,
            I => \N__37716\
        );

    \I__8674\ : InMux
    port map (
            O => \N__37768\,
            I => \N__37716\
        );

    \I__8673\ : InMux
    port map (
            O => \N__37767\,
            I => \N__37716\
        );

    \I__8672\ : InMux
    port map (
            O => \N__37766\,
            I => \N__37716\
        );

    \I__8671\ : InMux
    port map (
            O => \N__37765\,
            I => \N__37716\
        );

    \I__8670\ : InMux
    port map (
            O => \N__37764\,
            I => \N__37705\
        );

    \I__8669\ : InMux
    port map (
            O => \N__37763\,
            I => \N__37705\
        );

    \I__8668\ : InMux
    port map (
            O => \N__37762\,
            I => \N__37705\
        );

    \I__8667\ : InMux
    port map (
            O => \N__37761\,
            I => \N__37705\
        );

    \I__8666\ : InMux
    port map (
            O => \N__37760\,
            I => \N__37705\
        );

    \I__8665\ : InMux
    port map (
            O => \N__37759\,
            I => \N__37698\
        );

    \I__8664\ : InMux
    port map (
            O => \N__37758\,
            I => \N__37698\
        );

    \I__8663\ : InMux
    port map (
            O => \N__37757\,
            I => \N__37698\
        );

    \I__8662\ : LocalMux
    port map (
            O => \N__37748\,
            I => \N__37689\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__37745\,
            I => \N__37686\
        );

    \I__8660\ : LocalMux
    port map (
            O => \N__37734\,
            I => \N__37683\
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__37727\,
            I => \N__37680\
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__37716\,
            I => \N__37677\
        );

    \I__8657\ : LocalMux
    port map (
            O => \N__37705\,
            I => \N__37674\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__37698\,
            I => \N__37671\
        );

    \I__8655\ : CEMux
    port map (
            O => \N__37697\,
            I => \N__37644\
        );

    \I__8654\ : CEMux
    port map (
            O => \N__37696\,
            I => \N__37644\
        );

    \I__8653\ : CEMux
    port map (
            O => \N__37695\,
            I => \N__37644\
        );

    \I__8652\ : CEMux
    port map (
            O => \N__37694\,
            I => \N__37644\
        );

    \I__8651\ : CEMux
    port map (
            O => \N__37693\,
            I => \N__37644\
        );

    \I__8650\ : CEMux
    port map (
            O => \N__37692\,
            I => \N__37644\
        );

    \I__8649\ : Glb2LocalMux
    port map (
            O => \N__37689\,
            I => \N__37644\
        );

    \I__8648\ : Glb2LocalMux
    port map (
            O => \N__37686\,
            I => \N__37644\
        );

    \I__8647\ : Glb2LocalMux
    port map (
            O => \N__37683\,
            I => \N__37644\
        );

    \I__8646\ : Glb2LocalMux
    port map (
            O => \N__37680\,
            I => \N__37644\
        );

    \I__8645\ : Glb2LocalMux
    port map (
            O => \N__37677\,
            I => \N__37644\
        );

    \I__8644\ : Glb2LocalMux
    port map (
            O => \N__37674\,
            I => \N__37644\
        );

    \I__8643\ : Glb2LocalMux
    port map (
            O => \N__37671\,
            I => \N__37644\
        );

    \I__8642\ : GlobalMux
    port map (
            O => \N__37644\,
            I => \N__37641\
        );

    \I__8641\ : gio2CtrlBuf
    port map (
            O => \N__37641\,
            I => \HDA_STRAP.count_en_g\
        );

    \I__8640\ : InMux
    port map (
            O => \N__37638\,
            I => \N__37635\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__37635\,
            I => \N__37632\
        );

    \I__8638\ : Span4Mux_h
    port map (
            O => \N__37632\,
            I => \N__37629\
        );

    \I__8637\ : Odrv4
    port map (
            O => \N__37629\,
            I => \HDA_STRAP.un2_count_1_axb_8\
        );

    \I__8636\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37620\
        );

    \I__8635\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37620\
        );

    \I__8634\ : LocalMux
    port map (
            O => \N__37620\,
            I => \HDA_STRAP.count_3_1\
        );

    \I__8633\ : CascadeMux
    port map (
            O => \N__37617\,
            I => \HDA_STRAP.count_RNIZ0Z_1_cascade_\
        );

    \I__8632\ : InMux
    port map (
            O => \N__37614\,
            I => \N__37610\
        );

    \I__8631\ : InMux
    port map (
            O => \N__37613\,
            I => \N__37607\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__37610\,
            I => \N__37604\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__37607\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__8628\ : Odrv4
    port map (
            O => \N__37604\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__8627\ : InMux
    port map (
            O => \N__37599\,
            I => \N__37593\
        );

    \I__8626\ : InMux
    port map (
            O => \N__37598\,
            I => \N__37593\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__37593\,
            I => \N__37590\
        );

    \I__8624\ : Odrv4
    port map (
            O => \N__37590\,
            I => \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614\
        );

    \I__8623\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37584\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__37584\,
            I => \HDA_STRAP.count_3_2\
        );

    \I__8621\ : InMux
    port map (
            O => \N__37581\,
            I => \N__37577\
        );

    \I__8620\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37574\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__37577\,
            I => \HDA_STRAP.count_1_11\
        );

    \I__8618\ : LocalMux
    port map (
            O => \N__37574\,
            I => \HDA_STRAP.count_1_11\
        );

    \I__8617\ : InMux
    port map (
            O => \N__37569\,
            I => \N__37566\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__37566\,
            I => \HDA_STRAP.count_3_11\
        );

    \I__8615\ : InMux
    port map (
            O => \N__37563\,
            I => \N__37559\
        );

    \I__8614\ : InMux
    port map (
            O => \N__37562\,
            I => \N__37556\
        );

    \I__8613\ : LocalMux
    port map (
            O => \N__37559\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__8612\ : LocalMux
    port map (
            O => \N__37556\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__8611\ : InMux
    port map (
            O => \N__37551\,
            I => \N__37548\
        );

    \I__8610\ : LocalMux
    port map (
            O => \N__37548\,
            I => \HDA_STRAP.un25_clk_100khz_0\
        );

    \I__8609\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37542\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__37542\,
            I => \HDA_STRAP.un25_clk_100khz_1\
        );

    \I__8607\ : InMux
    port map (
            O => \N__37539\,
            I => \N__37536\
        );

    \I__8606\ : LocalMux
    port map (
            O => \N__37536\,
            I => \N__37533\
        );

    \I__8605\ : Span4Mux_s0_h
    port map (
            O => \N__37533\,
            I => \N__37529\
        );

    \I__8604\ : InMux
    port map (
            O => \N__37532\,
            I => \N__37526\
        );

    \I__8603\ : Odrv4
    port map (
            O => \N__37529\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__8602\ : LocalMux
    port map (
            O => \N__37526\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__8601\ : InMux
    port map (
            O => \N__37521\,
            I => \N__37518\
        );

    \I__8600\ : LocalMux
    port map (
            O => \N__37518\,
            I => \N__37515\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__37515\,
            I => \HDA_STRAP.un25_clk_100khz_6\
        );

    \I__8598\ : InMux
    port map (
            O => \N__37512\,
            I => \N__37509\
        );

    \I__8597\ : LocalMux
    port map (
            O => \N__37509\,
            I => \N__37506\
        );

    \I__8596\ : Odrv4
    port map (
            O => \N__37506\,
            I => \HDA_STRAP.un25_clk_100khz_14\
        );

    \I__8595\ : CascadeMux
    port map (
            O => \N__37503\,
            I => \HDA_STRAP.un25_clk_100khz_7_cascade_\
        );

    \I__8594\ : InMux
    port map (
            O => \N__37500\,
            I => \N__37497\
        );

    \I__8593\ : LocalMux
    port map (
            O => \N__37497\,
            I => \HDA_STRAP.un25_clk_100khz_13\
        );

    \I__8592\ : CascadeMux
    port map (
            O => \N__37494\,
            I => \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_\
        );

    \I__8591\ : CascadeMux
    port map (
            O => \N__37491\,
            I => \HDA_STRAP.count_1_0_cascade_\
        );

    \I__8590\ : CascadeMux
    port map (
            O => \N__37488\,
            I => \N__37484\
        );

    \I__8589\ : CascadeMux
    port map (
            O => \N__37487\,
            I => \N__37480\
        );

    \I__8588\ : InMux
    port map (
            O => \N__37484\,
            I => \N__37477\
        );

    \I__8587\ : InMux
    port map (
            O => \N__37483\,
            I => \N__37470\
        );

    \I__8586\ : InMux
    port map (
            O => \N__37480\,
            I => \N__37470\
        );

    \I__8585\ : LocalMux
    port map (
            O => \N__37477\,
            I => \N__37467\
        );

    \I__8584\ : InMux
    port map (
            O => \N__37476\,
            I => \N__37462\
        );

    \I__8583\ : InMux
    port map (
            O => \N__37475\,
            I => \N__37462\
        );

    \I__8582\ : LocalMux
    port map (
            O => \N__37470\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__8581\ : Odrv4
    port map (
            O => \N__37467\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__37462\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__8579\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37452\
        );

    \I__8578\ : LocalMux
    port map (
            O => \N__37452\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__8577\ : InMux
    port map (
            O => \N__37449\,
            I => \N__37443\
        );

    \I__8576\ : InMux
    port map (
            O => \N__37448\,
            I => \N__37443\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__37443\,
            I => \HDA_STRAP.count_3_9\
        );

    \I__8574\ : InMux
    port map (
            O => \N__37440\,
            I => \N__37431\
        );

    \I__8573\ : InMux
    port map (
            O => \N__37439\,
            I => \N__37431\
        );

    \I__8572\ : InMux
    port map (
            O => \N__37438\,
            I => \N__37431\
        );

    \I__8571\ : LocalMux
    port map (
            O => \N__37431\,
            I => \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84\
        );

    \I__8570\ : CascadeMux
    port map (
            O => \N__37428\,
            I => \HDA_STRAP.countZ0Z_12_cascade_\
        );

    \I__8569\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37422\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__37422\,
            I => \N__37419\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__37419\,
            I => \HDA_STRAP.un25_clk_100khz_4\
        );

    \I__8566\ : InMux
    port map (
            O => \N__37416\,
            I => \N__37413\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__37413\,
            I => \HDA_STRAP.un2_count_1_axb_5\
        );

    \I__8564\ : InMux
    port map (
            O => \N__37410\,
            I => \N__37405\
        );

    \I__8563\ : InMux
    port map (
            O => \N__37409\,
            I => \N__37400\
        );

    \I__8562\ : InMux
    port map (
            O => \N__37408\,
            I => \N__37400\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__37405\,
            I => \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__37400\,
            I => \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__8558\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37388\
        );

    \I__8557\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37385\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__37388\,
            I => \HDA_STRAP.count_3_5\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__37385\,
            I => \HDA_STRAP.count_3_5\
        );

    \I__8554\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37377\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__8552\ : Span4Mux_s3_v
    port map (
            O => \N__37374\,
            I => \N__37371\
        );

    \I__8551\ : Odrv4
    port map (
            O => \N__37371\,
            I => \HDA_STRAP.count_3_10\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__37368\,
            I => \N__37364\
        );

    \I__8549\ : InMux
    port map (
            O => \N__37367\,
            I => \N__37361\
        );

    \I__8548\ : InMux
    port map (
            O => \N__37364\,
            I => \N__37358\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__37361\,
            I => \N__37355\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__37358\,
            I => \HDA_STRAP.count_1_10\
        );

    \I__8545\ : Odrv4
    port map (
            O => \N__37355\,
            I => \HDA_STRAP.count_1_10\
        );

    \I__8544\ : CascadeMux
    port map (
            O => \N__37350\,
            I => \HDA_STRAP.un2_count_1_axb_1_cascade_\
        );

    \I__8543\ : InMux
    port map (
            O => \N__37347\,
            I => \N__37343\
        );

    \I__8542\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37340\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__37343\,
            I => \N__37337\
        );

    \I__8540\ : LocalMux
    port map (
            O => \N__37340\,
            I => \HDA_STRAP.un2_count_1_axb_1\
        );

    \I__8539\ : Odrv4
    port map (
            O => \N__37337\,
            I => \HDA_STRAP.un2_count_1_axb_1\
        );

    \I__8538\ : InMux
    port map (
            O => \N__37332\,
            I => \N__37329\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__37329\,
            I => \HDA_STRAP.count_RNIZ0Z_1\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__37326\,
            I => \HDA_STRAP.un25_clk_100khz_2_cascade_\
        );

    \I__8535\ : InMux
    port map (
            O => \N__37323\,
            I => \N__37319\
        );

    \I__8534\ : InMux
    port map (
            O => \N__37322\,
            I => \N__37316\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__37319\,
            I => \N__37313\
        );

    \I__8532\ : LocalMux
    port map (
            O => \N__37316\,
            I => \N__37310\
        );

    \I__8531\ : Span4Mux_v
    port map (
            O => \N__37313\,
            I => \N__37307\
        );

    \I__8530\ : Span4Mux_s2_h
    port map (
            O => \N__37310\,
            I => \N__37304\
        );

    \I__8529\ : Span4Mux_v
    port map (
            O => \N__37307\,
            I => \N__37301\
        );

    \I__8528\ : Span4Mux_v
    port map (
            O => \N__37304\,
            I => \N__37298\
        );

    \I__8527\ : Odrv4
    port map (
            O => \N__37301\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__37298\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__8525\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37290\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__37290\,
            I => \HDA_STRAP.un25_clk_100khz_5\
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__37287\,
            I => \N__37284\
        );

    \I__8522\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37278\
        );

    \I__8521\ : InMux
    port map (
            O => \N__37283\,
            I => \N__37278\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__37278\,
            I => \N__37275\
        );

    \I__8519\ : Odrv4
    port map (
            O => \N__37275\,
            I => \HDA_STRAP.count_3_13\
        );

    \I__8518\ : InMux
    port map (
            O => \N__37272\,
            I => \N__37265\
        );

    \I__8517\ : InMux
    port map (
            O => \N__37271\,
            I => \N__37265\
        );

    \I__8516\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37262\
        );

    \I__8515\ : LocalMux
    port map (
            O => \N__37265\,
            I => \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__37262\,
            I => \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\
        );

    \I__8513\ : InMux
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__37254\,
            I => \HDA_STRAP.un2_count_1_axb_13\
        );

    \I__8511\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37247\
        );

    \I__8510\ : InMux
    port map (
            O => \N__37250\,
            I => \N__37244\
        );

    \I__8509\ : LocalMux
    port map (
            O => \N__37247\,
            I => \N__37239\
        );

    \I__8508\ : LocalMux
    port map (
            O => \N__37244\,
            I => \N__37239\
        );

    \I__8507\ : Span4Mux_s2_h
    port map (
            O => \N__37239\,
            I => \N__37236\
        );

    \I__8506\ : Span4Mux_v
    port map (
            O => \N__37236\,
            I => \N__37233\
        );

    \I__8505\ : Odrv4
    port map (
            O => \N__37233\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__8504\ : InMux
    port map (
            O => \N__37230\,
            I => \N__37227\
        );

    \I__8503\ : LocalMux
    port map (
            O => \N__37227\,
            I => \HDA_STRAP.un25_clk_100khz_3\
        );

    \I__8502\ : InMux
    port map (
            O => \N__37224\,
            I => \N__37221\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__37221\,
            I => \HDA_STRAP.un2_count_1_axb_9\
        );

    \I__8500\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37215\
        );

    \I__8499\ : LocalMux
    port map (
            O => \N__37215\,
            I => \HDA_STRAP.count_3_12\
        );

    \I__8498\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37206\
        );

    \I__8497\ : InMux
    port map (
            O => \N__37211\,
            I => \N__37206\
        );

    \I__8496\ : LocalMux
    port map (
            O => \N__37206\,
            I => \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3\
        );

    \I__8495\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37200\
        );

    \I__8494\ : LocalMux
    port map (
            O => \N__37200\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__37197\,
            I => \N__37194\
        );

    \I__8492\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37191\
        );

    \I__8491\ : LocalMux
    port map (
            O => \N__37191\,
            I => \N__37188\
        );

    \I__8490\ : Span4Mux_h
    port map (
            O => \N__37188\,
            I => \N__37185\
        );

    \I__8489\ : Span4Mux_v
    port map (
            O => \N__37185\,
            I => \N__37182\
        );

    \I__8488\ : Odrv4
    port map (
            O => \N__37182\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__8487\ : InMux
    port map (
            O => \N__37179\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__8486\ : CascadeMux
    port map (
            O => \N__37176\,
            I => \N__37173\
        );

    \I__8485\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37170\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__37170\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__8483\ : InMux
    port map (
            O => \N__37167\,
            I => \N__37164\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__37164\,
            I => \N__37161\
        );

    \I__8481\ : Span4Mux_h
    port map (
            O => \N__37161\,
            I => \N__37158\
        );

    \I__8480\ : Span4Mux_v
    port map (
            O => \N__37158\,
            I => \N__37155\
        );

    \I__8479\ : Odrv4
    port map (
            O => \N__37155\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__8478\ : InMux
    port map (
            O => \N__37152\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__8477\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37146\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__37146\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__8475\ : CascadeMux
    port map (
            O => \N__37143\,
            I => \N__37140\
        );

    \I__8474\ : InMux
    port map (
            O => \N__37140\,
            I => \N__37137\
        );

    \I__8473\ : LocalMux
    port map (
            O => \N__37137\,
            I => \N__37134\
        );

    \I__8472\ : Span4Mux_v
    port map (
            O => \N__37134\,
            I => \N__37131\
        );

    \I__8471\ : Odrv4
    port map (
            O => \N__37131\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__8470\ : InMux
    port map (
            O => \N__37128\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__8469\ : CascadeMux
    port map (
            O => \N__37125\,
            I => \N__37122\
        );

    \I__8468\ : InMux
    port map (
            O => \N__37122\,
            I => \N__37119\
        );

    \I__8467\ : LocalMux
    port map (
            O => \N__37119\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__8466\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37113\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__37113\,
            I => \N__37110\
        );

    \I__8464\ : Span4Mux_v
    port map (
            O => \N__37110\,
            I => \N__37107\
        );

    \I__8463\ : Odrv4
    port map (
            O => \N__37107\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__8462\ : InMux
    port map (
            O => \N__37104\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__8461\ : InMux
    port map (
            O => \N__37101\,
            I => \N__37098\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__37098\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__8459\ : InMux
    port map (
            O => \N__37095\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__8458\ : CascadeMux
    port map (
            O => \N__37092\,
            I => \N__37089\
        );

    \I__8457\ : InMux
    port map (
            O => \N__37089\,
            I => \N__37080\
        );

    \I__8456\ : InMux
    port map (
            O => \N__37088\,
            I => \N__37080\
        );

    \I__8455\ : InMux
    port map (
            O => \N__37087\,
            I => \N__37080\
        );

    \I__8454\ : LocalMux
    port map (
            O => \N__37080\,
            I => \N__37077\
        );

    \I__8453\ : Span4Mux_v
    port map (
            O => \N__37077\,
            I => \N__37072\
        );

    \I__8452\ : InMux
    port map (
            O => \N__37076\,
            I => \N__37069\
        );

    \I__8451\ : InMux
    port map (
            O => \N__37075\,
            I => \N__37066\
        );

    \I__8450\ : Odrv4
    port map (
            O => \N__37072\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__37069\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__37066\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__8447\ : CascadeMux
    port map (
            O => \N__37059\,
            I => \N__37056\
        );

    \I__8446\ : InMux
    port map (
            O => \N__37056\,
            I => \N__37045\
        );

    \I__8445\ : InMux
    port map (
            O => \N__37055\,
            I => \N__37045\
        );

    \I__8444\ : InMux
    port map (
            O => \N__37054\,
            I => \N__37045\
        );

    \I__8443\ : InMux
    port map (
            O => \N__37053\,
            I => \N__37042\
        );

    \I__8442\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37039\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__37045\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__8440\ : LocalMux
    port map (
            O => \N__37042\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__37039\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__8438\ : CascadeMux
    port map (
            O => \N__37032\,
            I => \N__37028\
        );

    \I__8437\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37020\
        );

    \I__8436\ : InMux
    port map (
            O => \N__37028\,
            I => \N__37020\
        );

    \I__8435\ : InMux
    port map (
            O => \N__37027\,
            I => \N__37020\
        );

    \I__8434\ : LocalMux
    port map (
            O => \N__37020\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__8433\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37014\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__37014\,
            I => \HDA_STRAP.un2_count_1_axb_3\
        );

    \I__8431\ : InMux
    port map (
            O => \N__37011\,
            I => \N__37007\
        );

    \I__8430\ : InMux
    port map (
            O => \N__37010\,
            I => \N__37004\
        );

    \I__8429\ : LocalMux
    port map (
            O => \N__37007\,
            I => \N__36999\
        );

    \I__8428\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__36999\
        );

    \I__8427\ : Span4Mux_v
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__8426\ : Span4Mux_v
    port map (
            O => \N__36996\,
            I => \N__36993\
        );

    \I__8425\ : Odrv4
    port map (
            O => \N__36993\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__36990\,
            I => \N__36987\
        );

    \I__8423\ : InMux
    port map (
            O => \N__36987\,
            I => \N__36981\
        );

    \I__8422\ : InMux
    port map (
            O => \N__36986\,
            I => \N__36981\
        );

    \I__8421\ : LocalMux
    port map (
            O => \N__36981\,
            I => \HDA_STRAP.count_3_3\
        );

    \I__8420\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36969\
        );

    \I__8419\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36969\
        );

    \I__8418\ : InMux
    port map (
            O => \N__36976\,
            I => \N__36969\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__36969\,
            I => \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824\
        );

    \I__8416\ : InMux
    port map (
            O => \N__36966\,
            I => \N__36963\
        );

    \I__8415\ : LocalMux
    port map (
            O => \N__36963\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__8414\ : InMux
    port map (
            O => \N__36960\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__8413\ : CascadeMux
    port map (
            O => \N__36957\,
            I => \N__36954\
        );

    \I__8412\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36951\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__36951\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__8410\ : InMux
    port map (
            O => \N__36948\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__8409\ : InMux
    port map (
            O => \N__36945\,
            I => \N__36942\
        );

    \I__8408\ : LocalMux
    port map (
            O => \N__36942\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__8407\ : InMux
    port map (
            O => \N__36939\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__8406\ : CascadeMux
    port map (
            O => \N__36936\,
            I => \N__36933\
        );

    \I__8405\ : InMux
    port map (
            O => \N__36933\,
            I => \N__36930\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__36930\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__8403\ : InMux
    port map (
            O => \N__36927\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__8402\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36921\
        );

    \I__8401\ : LocalMux
    port map (
            O => \N__36921\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__8400\ : InMux
    port map (
            O => \N__36918\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__8399\ : CascadeMux
    port map (
            O => \N__36915\,
            I => \N__36912\
        );

    \I__8398\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36902\
        );

    \I__8397\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36902\
        );

    \I__8396\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36902\
        );

    \I__8395\ : InMux
    port map (
            O => \N__36909\,
            I => \N__36899\
        );

    \I__8394\ : LocalMux
    port map (
            O => \N__36902\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__36899\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__36894\,
            I => \N__36890\
        );

    \I__8391\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36882\
        );

    \I__8390\ : InMux
    port map (
            O => \N__36890\,
            I => \N__36882\
        );

    \I__8389\ : InMux
    port map (
            O => \N__36889\,
            I => \N__36882\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__36882\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__8387\ : InMux
    port map (
            O => \N__36879\,
            I => \N__36873\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__36878\,
            I => \N__36870\
        );

    \I__8385\ : InMux
    port map (
            O => \N__36877\,
            I => \N__36860\
        );

    \I__8384\ : CascadeMux
    port map (
            O => \N__36876\,
            I => \N__36856\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__36873\,
            I => \N__36851\
        );

    \I__8382\ : InMux
    port map (
            O => \N__36870\,
            I => \N__36842\
        );

    \I__8381\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36842\
        );

    \I__8380\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36842\
        );

    \I__8379\ : InMux
    port map (
            O => \N__36867\,
            I => \N__36842\
        );

    \I__8378\ : InMux
    port map (
            O => \N__36866\,
            I => \N__36833\
        );

    \I__8377\ : InMux
    port map (
            O => \N__36865\,
            I => \N__36833\
        );

    \I__8376\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36833\
        );

    \I__8375\ : InMux
    port map (
            O => \N__36863\,
            I => \N__36833\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__36860\,
            I => \N__36830\
        );

    \I__8373\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36827\
        );

    \I__8372\ : InMux
    port map (
            O => \N__36856\,
            I => \N__36824\
        );

    \I__8371\ : CascadeMux
    port map (
            O => \N__36855\,
            I => \N__36821\
        );

    \I__8370\ : CascadeMux
    port map (
            O => \N__36854\,
            I => \N__36818\
        );

    \I__8369\ : Span4Mux_h
    port map (
            O => \N__36851\,
            I => \N__36812\
        );

    \I__8368\ : LocalMux
    port map (
            O => \N__36842\,
            I => \N__36807\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__36833\,
            I => \N__36807\
        );

    \I__8366\ : Sp12to4
    port map (
            O => \N__36830\,
            I => \N__36802\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__36827\,
            I => \N__36802\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__36824\,
            I => \N__36799\
        );

    \I__8363\ : InMux
    port map (
            O => \N__36821\,
            I => \N__36796\
        );

    \I__8362\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36789\
        );

    \I__8361\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36789\
        );

    \I__8360\ : InMux
    port map (
            O => \N__36816\,
            I => \N__36789\
        );

    \I__8359\ : InMux
    port map (
            O => \N__36815\,
            I => \N__36786\
        );

    \I__8358\ : Span4Mux_h
    port map (
            O => \N__36812\,
            I => \N__36783\
        );

    \I__8357\ : Span12Mux_s11_h
    port map (
            O => \N__36807\,
            I => \N__36780\
        );

    \I__8356\ : Span12Mux_s7_h
    port map (
            O => \N__36802\,
            I => \N__36775\
        );

    \I__8355\ : Span12Mux_s4_v
    port map (
            O => \N__36799\,
            I => \N__36775\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__36796\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__36789\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__36786\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__8351\ : Odrv4
    port map (
            O => \N__36783\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__8350\ : Odrv12
    port map (
            O => \N__36780\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__8349\ : Odrv12
    port map (
            O => \N__36775\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__8348\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36755\
        );

    \I__8347\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36752\
        );

    \I__8346\ : CascadeMux
    port map (
            O => \N__36760\,
            I => \N__36746\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__36759\,
            I => \N__36743\
        );

    \I__8344\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36739\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__36755\,
            I => \N__36733\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__36752\,
            I => \N__36733\
        );

    \I__8341\ : InMux
    port map (
            O => \N__36751\,
            I => \N__36729\
        );

    \I__8340\ : InMux
    port map (
            O => \N__36750\,
            I => \N__36722\
        );

    \I__8339\ : InMux
    port map (
            O => \N__36749\,
            I => \N__36722\
        );

    \I__8338\ : InMux
    port map (
            O => \N__36746\,
            I => \N__36717\
        );

    \I__8337\ : InMux
    port map (
            O => \N__36743\,
            I => \N__36717\
        );

    \I__8336\ : InMux
    port map (
            O => \N__36742\,
            I => \N__36713\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__36739\,
            I => \N__36710\
        );

    \I__8334\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36707\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__36733\,
            I => \N__36704\
        );

    \I__8332\ : InMux
    port map (
            O => \N__36732\,
            I => \N__36701\
        );

    \I__8331\ : LocalMux
    port map (
            O => \N__36729\,
            I => \N__36698\
        );

    \I__8330\ : InMux
    port map (
            O => \N__36728\,
            I => \N__36693\
        );

    \I__8329\ : InMux
    port map (
            O => \N__36727\,
            I => \N__36693\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__36722\,
            I => \N__36688\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__36717\,
            I => \N__36688\
        );

    \I__8326\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36685\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__36713\,
            I => \N__36682\
        );

    \I__8324\ : Span4Mux_h
    port map (
            O => \N__36710\,
            I => \N__36679\
        );

    \I__8323\ : LocalMux
    port map (
            O => \N__36707\,
            I => \N__36675\
        );

    \I__8322\ : Span4Mux_s1_h
    port map (
            O => \N__36704\,
            I => \N__36664\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__36701\,
            I => \N__36664\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__36698\,
            I => \N__36664\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36664\
        );

    \I__8318\ : Span4Mux_v
    port map (
            O => \N__36688\,
            I => \N__36664\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__36685\,
            I => \N__36661\
        );

    \I__8316\ : Span4Mux_v
    port map (
            O => \N__36682\,
            I => \N__36658\
        );

    \I__8315\ : Sp12to4
    port map (
            O => \N__36679\,
            I => \N__36655\
        );

    \I__8314\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36652\
        );

    \I__8313\ : Span4Mux_h
    port map (
            O => \N__36675\,
            I => \N__36649\
        );

    \I__8312\ : Span4Mux_h
    port map (
            O => \N__36664\,
            I => \N__36646\
        );

    \I__8311\ : Span4Mux_s1_h
    port map (
            O => \N__36661\,
            I => \N__36643\
        );

    \I__8310\ : Odrv4
    port map (
            O => \N__36658\,
            I => \POWERLED.N_203_i\
        );

    \I__8309\ : Odrv12
    port map (
            O => \N__36655\,
            I => \POWERLED.N_203_i\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__36652\,
            I => \POWERLED.N_203_i\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__36649\,
            I => \POWERLED.N_203_i\
        );

    \I__8306\ : Odrv4
    port map (
            O => \N__36646\,
            I => \POWERLED.N_203_i\
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__36643\,
            I => \POWERLED.N_203_i\
        );

    \I__8304\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36627\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__36627\,
            I => \N__36624\
        );

    \I__8302\ : Span4Mux_h
    port map (
            O => \N__36624\,
            I => \N__36621\
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__36621\,
            I => \POWERLED.g0_9_0\
        );

    \I__8300\ : CascadeMux
    port map (
            O => \N__36618\,
            I => \N__36615\
        );

    \I__8299\ : InMux
    port map (
            O => \N__36615\,
            I => \N__36612\
        );

    \I__8298\ : LocalMux
    port map (
            O => \N__36612\,
            I => \N__36609\
        );

    \I__8297\ : Span12Mux_s4_h
    port map (
            O => \N__36609\,
            I => \N__36606\
        );

    \I__8296\ : Odrv12
    port map (
            O => \N__36606\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__8295\ : InMux
    port map (
            O => \N__36603\,
            I => \N__36600\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__36600\,
            I => \N__36597\
        );

    \I__8293\ : Span4Mux_v
    port map (
            O => \N__36597\,
            I => \N__36594\
        );

    \I__8292\ : Odrv4
    port map (
            O => \N__36594\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__8291\ : InMux
    port map (
            O => \N__36591\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__8290\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36585\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__36585\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__8288\ : InMux
    port map (
            O => \N__36582\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__8287\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36576\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__36576\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__8285\ : InMux
    port map (
            O => \N__36573\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__8284\ : CascadeMux
    port map (
            O => \N__36570\,
            I => \N__36564\
        );

    \I__8283\ : InMux
    port map (
            O => \N__36569\,
            I => \N__36558\
        );

    \I__8282\ : InMux
    port map (
            O => \N__36568\,
            I => \N__36558\
        );

    \I__8281\ : InMux
    port map (
            O => \N__36567\,
            I => \N__36553\
        );

    \I__8280\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36553\
        );

    \I__8279\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36550\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__36558\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__36553\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__36550\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__36543\,
            I => \N__36540\
        );

    \I__8274\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36537\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__36537\,
            I => \N__36534\
        );

    \I__8272\ : Odrv4
    port map (
            O => \N__36534\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__8271\ : InMux
    port map (
            O => \N__36531\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__8270\ : CascadeMux
    port map (
            O => \N__36528\,
            I => \N__36524\
        );

    \I__8269\ : InMux
    port map (
            O => \N__36527\,
            I => \N__36516\
        );

    \I__8268\ : InMux
    port map (
            O => \N__36524\,
            I => \N__36516\
        );

    \I__8267\ : InMux
    port map (
            O => \N__36523\,
            I => \N__36516\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__36516\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__36513\,
            I => \N__36510\
        );

    \I__8264\ : InMux
    port map (
            O => \N__36510\,
            I => \N__36507\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__36507\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__8262\ : InMux
    port map (
            O => \N__36504\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__8261\ : InMux
    port map (
            O => \N__36501\,
            I => \N__36498\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__36498\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__8259\ : InMux
    port map (
            O => \N__36495\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__8258\ : CascadeMux
    port map (
            O => \N__36492\,
            I => \POWERLED.mult1_un145_sum_s_8_cascade_\
        );

    \I__8257\ : InMux
    port map (
            O => \N__36489\,
            I => \N__36486\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__36486\,
            I => \N__36483\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__36483\,
            I => \N__36480\
        );

    \I__8254\ : Odrv4
    port map (
            O => \N__36480\,
            I => \POWERLED.un85_clk_100khz_3\
        );

    \I__8253\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36472\
        );

    \I__8252\ : CascadeMux
    port map (
            O => \N__36476\,
            I => \N__36469\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__36475\,
            I => \N__36465\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__36472\,
            I => \N__36460\
        );

    \I__8249\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36455\
        );

    \I__8248\ : InMux
    port map (
            O => \N__36468\,
            I => \N__36452\
        );

    \I__8247\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36447\
        );

    \I__8246\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36447\
        );

    \I__8245\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36444\
        );

    \I__8244\ : Span4Mux_s3_h
    port map (
            O => \N__36460\,
            I => \N__36440\
        );

    \I__8243\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36434\
        );

    \I__8242\ : InMux
    port map (
            O => \N__36458\,
            I => \N__36434\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__36455\,
            I => \N__36429\
        );

    \I__8240\ : LocalMux
    port map (
            O => \N__36452\,
            I => \N__36429\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__36447\,
            I => \N__36426\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__36444\,
            I => \N__36423\
        );

    \I__8237\ : InMux
    port map (
            O => \N__36443\,
            I => \N__36420\
        );

    \I__8236\ : Sp12to4
    port map (
            O => \N__36440\,
            I => \N__36415\
        );

    \I__8235\ : InMux
    port map (
            O => \N__36439\,
            I => \N__36412\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__36434\,
            I => \N__36409\
        );

    \I__8233\ : Span4Mux_h
    port map (
            O => \N__36429\,
            I => \N__36406\
        );

    \I__8232\ : Span4Mux_v
    port map (
            O => \N__36426\,
            I => \N__36399\
        );

    \I__8231\ : Span4Mux_s3_v
    port map (
            O => \N__36423\,
            I => \N__36399\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__36420\,
            I => \N__36399\
        );

    \I__8229\ : InMux
    port map (
            O => \N__36419\,
            I => \N__36394\
        );

    \I__8228\ : InMux
    port map (
            O => \N__36418\,
            I => \N__36394\
        );

    \I__8227\ : Span12Mux_s4_v
    port map (
            O => \N__36415\,
            I => \N__36391\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__36412\,
            I => \N__36388\
        );

    \I__8225\ : Span4Mux_v
    port map (
            O => \N__36409\,
            I => \N__36383\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__36406\,
            I => \N__36383\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__36399\,
            I => \N__36380\
        );

    \I__8222\ : LocalMux
    port map (
            O => \N__36394\,
            I => \N__36377\
        );

    \I__8221\ : Odrv12
    port map (
            O => \N__36391\,
            I => \POWERLED.dutycycle\
        );

    \I__8220\ : Odrv4
    port map (
            O => \N__36388\,
            I => \POWERLED.dutycycle\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__36383\,
            I => \POWERLED.dutycycle\
        );

    \I__8218\ : Odrv4
    port map (
            O => \N__36380\,
            I => \POWERLED.dutycycle\
        );

    \I__8217\ : Odrv4
    port map (
            O => \N__36377\,
            I => \POWERLED.dutycycle\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__36366\,
            I => \N__36363\
        );

    \I__8215\ : InMux
    port map (
            O => \N__36363\,
            I => \N__36360\
        );

    \I__8214\ : LocalMux
    port map (
            O => \N__36360\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__8213\ : InMux
    port map (
            O => \N__36357\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__36354\,
            I => \N__36351\
        );

    \I__8211\ : InMux
    port map (
            O => \N__36351\,
            I => \N__36348\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__36348\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__8209\ : InMux
    port map (
            O => \N__36345\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__8208\ : InMux
    port map (
            O => \N__36342\,
            I => \N__36339\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__36339\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__8206\ : InMux
    port map (
            O => \N__36336\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__8205\ : CascadeMux
    port map (
            O => \N__36333\,
            I => \N__36330\
        );

    \I__8204\ : InMux
    port map (
            O => \N__36330\,
            I => \N__36327\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__36327\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__8202\ : InMux
    port map (
            O => \N__36324\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__8201\ : InMux
    port map (
            O => \N__36321\,
            I => \N__36318\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__36318\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__8199\ : InMux
    port map (
            O => \N__36315\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__36312\,
            I => \N__36309\
        );

    \I__8197\ : InMux
    port map (
            O => \N__36309\,
            I => \N__36306\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__36306\,
            I => \N__36303\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__36303\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__8194\ : InMux
    port map (
            O => \N__36300\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__8193\ : InMux
    port map (
            O => \N__36297\,
            I => \N__36294\
        );

    \I__8192\ : LocalMux
    port map (
            O => \N__36294\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__8191\ : InMux
    port map (
            O => \N__36291\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__36288\,
            I => \N__36285\
        );

    \I__8189\ : InMux
    port map (
            O => \N__36285\,
            I => \N__36275\
        );

    \I__8188\ : InMux
    port map (
            O => \N__36284\,
            I => \N__36275\
        );

    \I__8187\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36275\
        );

    \I__8186\ : InMux
    port map (
            O => \N__36282\,
            I => \N__36272\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__36275\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__36272\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__8183\ : CascadeMux
    port map (
            O => \N__36267\,
            I => \N__36263\
        );

    \I__8182\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36255\
        );

    \I__8181\ : InMux
    port map (
            O => \N__36263\,
            I => \N__36255\
        );

    \I__8180\ : InMux
    port map (
            O => \N__36262\,
            I => \N__36255\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__36255\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__8178\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36249\
        );

    \I__8177\ : LocalMux
    port map (
            O => \N__36249\,
            I => \N__36245\
        );

    \I__8176\ : InMux
    port map (
            O => \N__36248\,
            I => \N__36242\
        );

    \I__8175\ : Span4Mux_v
    port map (
            O => \N__36245\,
            I => \N__36239\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__36242\,
            I => \N__36236\
        );

    \I__8173\ : Sp12to4
    port map (
            O => \N__36239\,
            I => \N__36233\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__36236\,
            I => \N__36230\
        );

    \I__8171\ : Odrv12
    port map (
            O => \N__36233\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__8170\ : Odrv4
    port map (
            O => \N__36230\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__8169\ : CascadeMux
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__8168\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36219\
        );

    \I__8167\ : LocalMux
    port map (
            O => \N__36219\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__8166\ : InMux
    port map (
            O => \N__36216\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__8165\ : CascadeMux
    port map (
            O => \N__36213\,
            I => \N__36209\
        );

    \I__8164\ : CascadeMux
    port map (
            O => \N__36212\,
            I => \N__36206\
        );

    \I__8163\ : InMux
    port map (
            O => \N__36209\,
            I => \N__36203\
        );

    \I__8162\ : InMux
    port map (
            O => \N__36206\,
            I => \N__36199\
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__36203\,
            I => \N__36196\
        );

    \I__8160\ : InMux
    port map (
            O => \N__36202\,
            I => \N__36193\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__36199\,
            I => \N__36190\
        );

    \I__8158\ : Span4Mux_s2_h
    port map (
            O => \N__36196\,
            I => \N__36181\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__36193\,
            I => \N__36181\
        );

    \I__8156\ : Span4Mux_s2_h
    port map (
            O => \N__36190\,
            I => \N__36181\
        );

    \I__8155\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36177\
        );

    \I__8154\ : CascadeMux
    port map (
            O => \N__36188\,
            I => \N__36174\
        );

    \I__8153\ : Span4Mux_h
    port map (
            O => \N__36181\,
            I => \N__36168\
        );

    \I__8152\ : InMux
    port map (
            O => \N__36180\,
            I => \N__36165\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__36177\,
            I => \N__36162\
        );

    \I__8150\ : InMux
    port map (
            O => \N__36174\,
            I => \N__36157\
        );

    \I__8149\ : InMux
    port map (
            O => \N__36173\,
            I => \N__36157\
        );

    \I__8148\ : InMux
    port map (
            O => \N__36172\,
            I => \N__36152\
        );

    \I__8147\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36152\
        );

    \I__8146\ : Span4Mux_h
    port map (
            O => \N__36168\,
            I => \N__36147\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__36165\,
            I => \N__36147\
        );

    \I__8144\ : Odrv12
    port map (
            O => \N__36162\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__36157\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__8142\ : LocalMux
    port map (
            O => \N__36152\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__8141\ : Odrv4
    port map (
            O => \N__36147\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__8140\ : IoInMux
    port map (
            O => \N__36138\,
            I => \N__36135\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__36135\,
            I => \N__36132\
        );

    \I__8138\ : Span4Mux_s0_h
    port map (
            O => \N__36132\,
            I => \N__36129\
        );

    \I__8137\ : Span4Mux_v
    port map (
            O => \N__36129\,
            I => \N__36126\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__36126\,
            I => vpp_en
        );

    \I__8135\ : InMux
    port map (
            O => \N__36123\,
            I => \N__36120\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__36120\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__8133\ : InMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__8132\ : LocalMux
    port map (
            O => \N__36114\,
            I => \N__36109\
        );

    \I__8131\ : InMux
    port map (
            O => \N__36113\,
            I => \N__36104\
        );

    \I__8130\ : InMux
    port map (
            O => \N__36112\,
            I => \N__36104\
        );

    \I__8129\ : Span4Mux_v
    port map (
            O => \N__36109\,
            I => \N__36101\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__36104\,
            I => \N__36098\
        );

    \I__8127\ : Span4Mux_h
    port map (
            O => \N__36101\,
            I => \N__36095\
        );

    \I__8126\ : Odrv12
    port map (
            O => \N__36098\,
            I => \VPP_VDDQ.N_194\
        );

    \I__8125\ : Odrv4
    port map (
            O => \N__36095\,
            I => \VPP_VDDQ.N_194\
        );

    \I__8124\ : InMux
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__36087\,
            I => \VPP_VDDQ.curr_state_0_0\
        );

    \I__8122\ : InMux
    port map (
            O => \N__36084\,
            I => \N__36081\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__36081\,
            I => \N__36078\
        );

    \I__8120\ : Odrv12
    port map (
            O => \N__36078\,
            I => \VPP_VDDQ.un4_count_1_axb_2\
        );

    \I__8119\ : InMux
    port map (
            O => \N__36075\,
            I => \N__36068\
        );

    \I__8118\ : InMux
    port map (
            O => \N__36074\,
            I => \N__36059\
        );

    \I__8117\ : InMux
    port map (
            O => \N__36073\,
            I => \N__36059\
        );

    \I__8116\ : InMux
    port map (
            O => \N__36072\,
            I => \N__36059\
        );

    \I__8115\ : InMux
    port map (
            O => \N__36071\,
            I => \N__36059\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__36068\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__36059\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__8112\ : InMux
    port map (
            O => \N__36054\,
            I => \N__36038\
        );

    \I__8111\ : InMux
    port map (
            O => \N__36053\,
            I => \N__36035\
        );

    \I__8110\ : InMux
    port map (
            O => \N__36052\,
            I => \N__36032\
        );

    \I__8109\ : InMux
    port map (
            O => \N__36051\,
            I => \N__36027\
        );

    \I__8108\ : InMux
    port map (
            O => \N__36050\,
            I => \N__36027\
        );

    \I__8107\ : InMux
    port map (
            O => \N__36049\,
            I => \N__36020\
        );

    \I__8106\ : InMux
    port map (
            O => \N__36048\,
            I => \N__36020\
        );

    \I__8105\ : InMux
    port map (
            O => \N__36047\,
            I => \N__36020\
        );

    \I__8104\ : InMux
    port map (
            O => \N__36046\,
            I => \N__36017\
        );

    \I__8103\ : InMux
    port map (
            O => \N__36045\,
            I => \N__36014\
        );

    \I__8102\ : InMux
    port map (
            O => \N__36044\,
            I => \N__36011\
        );

    \I__8101\ : InMux
    port map (
            O => \N__36043\,
            I => \N__36006\
        );

    \I__8100\ : InMux
    port map (
            O => \N__36042\,
            I => \N__36006\
        );

    \I__8099\ : InMux
    port map (
            O => \N__36041\,
            I => \N__36003\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__36038\,
            I => \N__35985\
        );

    \I__8097\ : LocalMux
    port map (
            O => \N__36035\,
            I => \N__35982\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__36032\,
            I => \N__35979\
        );

    \I__8095\ : LocalMux
    port map (
            O => \N__36027\,
            I => \N__35976\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__36020\,
            I => \N__35973\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__36017\,
            I => \N__35970\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__36014\,
            I => \N__35967\
        );

    \I__8091\ : LocalMux
    port map (
            O => \N__36011\,
            I => \N__35964\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__36006\,
            I => \N__35961\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__36003\,
            I => \N__35958\
        );

    \I__8088\ : CEMux
    port map (
            O => \N__36002\,
            I => \N__35907\
        );

    \I__8087\ : CEMux
    port map (
            O => \N__36001\,
            I => \N__35907\
        );

    \I__8086\ : CEMux
    port map (
            O => \N__36000\,
            I => \N__35907\
        );

    \I__8085\ : CEMux
    port map (
            O => \N__35999\,
            I => \N__35907\
        );

    \I__8084\ : CEMux
    port map (
            O => \N__35998\,
            I => \N__35907\
        );

    \I__8083\ : CEMux
    port map (
            O => \N__35997\,
            I => \N__35907\
        );

    \I__8082\ : CEMux
    port map (
            O => \N__35996\,
            I => \N__35907\
        );

    \I__8081\ : CEMux
    port map (
            O => \N__35995\,
            I => \N__35907\
        );

    \I__8080\ : CEMux
    port map (
            O => \N__35994\,
            I => \N__35907\
        );

    \I__8079\ : CEMux
    port map (
            O => \N__35993\,
            I => \N__35907\
        );

    \I__8078\ : CEMux
    port map (
            O => \N__35992\,
            I => \N__35907\
        );

    \I__8077\ : CEMux
    port map (
            O => \N__35991\,
            I => \N__35907\
        );

    \I__8076\ : CEMux
    port map (
            O => \N__35990\,
            I => \N__35907\
        );

    \I__8075\ : CEMux
    port map (
            O => \N__35989\,
            I => \N__35907\
        );

    \I__8074\ : CEMux
    port map (
            O => \N__35988\,
            I => \N__35907\
        );

    \I__8073\ : Glb2LocalMux
    port map (
            O => \N__35985\,
            I => \N__35907\
        );

    \I__8072\ : Glb2LocalMux
    port map (
            O => \N__35982\,
            I => \N__35907\
        );

    \I__8071\ : Glb2LocalMux
    port map (
            O => \N__35979\,
            I => \N__35907\
        );

    \I__8070\ : Glb2LocalMux
    port map (
            O => \N__35976\,
            I => \N__35907\
        );

    \I__8069\ : Glb2LocalMux
    port map (
            O => \N__35973\,
            I => \N__35907\
        );

    \I__8068\ : Glb2LocalMux
    port map (
            O => \N__35970\,
            I => \N__35907\
        );

    \I__8067\ : Glb2LocalMux
    port map (
            O => \N__35967\,
            I => \N__35907\
        );

    \I__8066\ : Glb2LocalMux
    port map (
            O => \N__35964\,
            I => \N__35907\
        );

    \I__8065\ : Glb2LocalMux
    port map (
            O => \N__35961\,
            I => \N__35907\
        );

    \I__8064\ : Glb2LocalMux
    port map (
            O => \N__35958\,
            I => \N__35907\
        );

    \I__8063\ : GlobalMux
    port map (
            O => \N__35907\,
            I => \N__35904\
        );

    \I__8062\ : gio2CtrlBuf
    port map (
            O => \N__35904\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en_g\
        );

    \I__8061\ : CEMux
    port map (
            O => \N__35901\,
            I => \N__35898\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__35898\,
            I => \N__35894\
        );

    \I__8059\ : CEMux
    port map (
            O => \N__35897\,
            I => \N__35873\
        );

    \I__8058\ : Span4Mux_s3_h
    port map (
            O => \N__35894\,
            I => \N__35870\
        );

    \I__8057\ : CEMux
    port map (
            O => \N__35893\,
            I => \N__35867\
        );

    \I__8056\ : CEMux
    port map (
            O => \N__35892\,
            I => \N__35864\
        );

    \I__8055\ : CEMux
    port map (
            O => \N__35891\,
            I => \N__35861\
        );

    \I__8054\ : InMux
    port map (
            O => \N__35890\,
            I => \N__35852\
        );

    \I__8053\ : InMux
    port map (
            O => \N__35889\,
            I => \N__35852\
        );

    \I__8052\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35852\
        );

    \I__8051\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35852\
        );

    \I__8050\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35843\
        );

    \I__8049\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35843\
        );

    \I__8048\ : InMux
    port map (
            O => \N__35884\,
            I => \N__35843\
        );

    \I__8047\ : InMux
    port map (
            O => \N__35883\,
            I => \N__35843\
        );

    \I__8046\ : InMux
    port map (
            O => \N__35882\,
            I => \N__35832\
        );

    \I__8045\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35832\
        );

    \I__8044\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35832\
        );

    \I__8043\ : InMux
    port map (
            O => \N__35879\,
            I => \N__35832\
        );

    \I__8042\ : InMux
    port map (
            O => \N__35878\,
            I => \N__35832\
        );

    \I__8041\ : InMux
    port map (
            O => \N__35877\,
            I => \N__35829\
        );

    \I__8040\ : CEMux
    port map (
            O => \N__35876\,
            I => \N__35826\
        );

    \I__8039\ : LocalMux
    port map (
            O => \N__35873\,
            I => \N__35823\
        );

    \I__8038\ : Span4Mux_h
    port map (
            O => \N__35870\,
            I => \N__35820\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__35867\,
            I => \N__35815\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__35864\,
            I => \N__35802\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__35861\,
            I => \N__35802\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__35852\,
            I => \N__35802\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__35843\,
            I => \N__35802\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__35832\,
            I => \N__35802\
        );

    \I__8031\ : LocalMux
    port map (
            O => \N__35829\,
            I => \N__35802\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__35826\,
            I => \N__35797\
        );

    \I__8029\ : Span4Mux_v
    port map (
            O => \N__35823\,
            I => \N__35797\
        );

    \I__8028\ : Span4Mux_v
    port map (
            O => \N__35820\,
            I => \N__35794\
        );

    \I__8027\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35791\
        );

    \I__8026\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35788\
        );

    \I__8025\ : Span4Mux_v
    port map (
            O => \N__35815\,
            I => \N__35783\
        );

    \I__8024\ : Span4Mux_v
    port map (
            O => \N__35802\,
            I => \N__35783\
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__35797\,
            I => \VPP_VDDQ.count_en\
        );

    \I__8022\ : Odrv4
    port map (
            O => \N__35794\,
            I => \VPP_VDDQ.count_en\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__35791\,
            I => \VPP_VDDQ.count_en\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__35788\,
            I => \VPP_VDDQ.count_en\
        );

    \I__8019\ : Odrv4
    port map (
            O => \N__35783\,
            I => \VPP_VDDQ.count_en\
        );

    \I__8018\ : InMux
    port map (
            O => \N__35772\,
            I => \N__35766\
        );

    \I__8017\ : InMux
    port map (
            O => \N__35771\,
            I => \N__35766\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__35766\,
            I => \VPP_VDDQ.count_4_2\
        );

    \I__8015\ : CascadeMux
    port map (
            O => \N__35763\,
            I => \VPP_VDDQ.count_en_cascade_\
        );

    \I__8014\ : InMux
    port map (
            O => \N__35760\,
            I => \N__35755\
        );

    \I__8013\ : InMux
    port map (
            O => \N__35759\,
            I => \N__35750\
        );

    \I__8012\ : InMux
    port map (
            O => \N__35758\,
            I => \N__35750\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35745\
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__35750\,
            I => \N__35745\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__35745\,
            I => \N__35742\
        );

    \I__8008\ : Odrv4
    port map (
            O => \N__35742\,
            I => \VPP_VDDQ.count_rst_7\
        );

    \I__8007\ : InMux
    port map (
            O => \N__35739\,
            I => \N__35735\
        );

    \I__8006\ : InMux
    port map (
            O => \N__35738\,
            I => \N__35732\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__35735\,
            I => \N__35729\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__35732\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__8003\ : Odrv4
    port map (
            O => \N__35729\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__8002\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35721\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__35721\,
            I => \N__35717\
        );

    \I__8000\ : InMux
    port map (
            O => \N__35720\,
            I => \N__35714\
        );

    \I__7999\ : Odrv4
    port map (
            O => \N__35717\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__35714\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__7997\ : CascadeMux
    port map (
            O => \N__35709\,
            I => \VPP_VDDQ.countZ0Z_2_cascade_\
        );

    \I__7996\ : CascadeMux
    port map (
            O => \N__35706\,
            I => \N__35702\
        );

    \I__7995\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35699\
        );

    \I__7994\ : InMux
    port map (
            O => \N__35702\,
            I => \N__35696\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__35699\,
            I => \N__35693\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__35696\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__7991\ : Odrv4
    port map (
            O => \N__35693\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__7990\ : InMux
    port map (
            O => \N__35688\,
            I => \N__35685\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__35685\,
            I => \N__35682\
        );

    \I__7988\ : Span4Mux_v
    port map (
            O => \N__35682\,
            I => \N__35679\
        );

    \I__7987\ : Odrv4
    port map (
            O => \N__35679\,
            I => \VPP_VDDQ.un13_clk_100khz_11\
        );

    \I__7986\ : InMux
    port map (
            O => \N__35676\,
            I => \N__35673\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__35673\,
            I => \N__35669\
        );

    \I__7984\ : InMux
    port map (
            O => \N__35672\,
            I => \N__35666\
        );

    \I__7983\ : Span4Mux_s1_h
    port map (
            O => \N__35669\,
            I => \N__35661\
        );

    \I__7982\ : LocalMux
    port map (
            O => \N__35666\,
            I => \N__35661\
        );

    \I__7981\ : Span4Mux_v
    port map (
            O => \N__35661\,
            I => \N__35658\
        );

    \I__7980\ : Odrv4
    port map (
            O => \N__35658\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__7979\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35652\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__35652\,
            I => \N__35648\
        );

    \I__7977\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35645\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__35648\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__7975\ : LocalMux
    port map (
            O => \N__35645\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__7974\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35634\
        );

    \I__7973\ : InMux
    port map (
            O => \N__35639\,
            I => \N__35634\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__35634\,
            I => \VPP_VDDQ.count_rst_3\
        );

    \I__7971\ : InMux
    port map (
            O => \N__35631\,
            I => \VPP_VDDQ.un4_count_1_cry_13\
        );

    \I__7970\ : InMux
    port map (
            O => \N__35628\,
            I => \N__35624\
        );

    \I__7969\ : InMux
    port map (
            O => \N__35627\,
            I => \N__35621\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__35624\,
            I => \N__35618\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__35621\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__7966\ : Odrv4
    port map (
            O => \N__35618\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__7965\ : InMux
    port map (
            O => \N__35613\,
            I => \VPP_VDDQ.un4_count_1_cry_14\
        );

    \I__7964\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35604\
        );

    \I__7963\ : InMux
    port map (
            O => \N__35609\,
            I => \N__35604\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__35604\,
            I => \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0\
        );

    \I__7961\ : InMux
    port map (
            O => \N__35601\,
            I => \N__35597\
        );

    \I__7960\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35594\
        );

    \I__7959\ : LocalMux
    port map (
            O => \N__35597\,
            I => \VPP_VDDQ.count_rst_2\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__35594\,
            I => \VPP_VDDQ.count_rst_2\
        );

    \I__7957\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35586\
        );

    \I__7956\ : LocalMux
    port map (
            O => \N__35586\,
            I => \VPP_VDDQ.count_4_13\
        );

    \I__7955\ : InMux
    port map (
            O => \N__35583\,
            I => \N__35579\
        );

    \I__7954\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35576\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__35579\,
            I => \VPP_VDDQ.count_rst_1\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__35576\,
            I => \VPP_VDDQ.count_rst_1\
        );

    \I__7951\ : InMux
    port map (
            O => \N__35571\,
            I => \N__35568\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__35568\,
            I => \N__35565\
        );

    \I__7949\ : Odrv4
    port map (
            O => \N__35565\,
            I => \VPP_VDDQ.count_4_12\
        );

    \I__7948\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35559\
        );

    \I__7947\ : LocalMux
    port map (
            O => \N__35559\,
            I => \N__35555\
        );

    \I__7946\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35552\
        );

    \I__7945\ : Odrv4
    port map (
            O => \N__35555\,
            I => \VPP_VDDQ.count_rst_8\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__35552\,
            I => \VPP_VDDQ.count_rst_8\
        );

    \I__7943\ : InMux
    port map (
            O => \N__35547\,
            I => \N__35544\
        );

    \I__7942\ : LocalMux
    port map (
            O => \N__35544\,
            I => \N__35541\
        );

    \I__7941\ : Odrv4
    port map (
            O => \N__35541\,
            I => \VPP_VDDQ.count_4_3\
        );

    \I__7940\ : InMux
    port map (
            O => \N__35538\,
            I => \N__35534\
        );

    \I__7939\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35531\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__35534\,
            I => \N__35528\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__35531\,
            I => \VPP_VDDQ.count_rst_9\
        );

    \I__7936\ : Odrv12
    port map (
            O => \N__35528\,
            I => \VPP_VDDQ.count_rst_9\
        );

    \I__7935\ : InMux
    port map (
            O => \N__35523\,
            I => \N__35520\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35517\
        );

    \I__7933\ : Odrv4
    port map (
            O => \N__35517\,
            I => \VPP_VDDQ.count_4_4\
        );

    \I__7932\ : InMux
    port map (
            O => \N__35514\,
            I => \N__35510\
        );

    \I__7931\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35507\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__35510\,
            I => \N__35504\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__35507\,
            I => \N__35501\
        );

    \I__7928\ : Span4Mux_v
    port map (
            O => \N__35504\,
            I => \N__35498\
        );

    \I__7927\ : Span4Mux_v
    port map (
            O => \N__35501\,
            I => \N__35494\
        );

    \I__7926\ : Span4Mux_v
    port map (
            O => \N__35498\,
            I => \N__35491\
        );

    \I__7925\ : InMux
    port map (
            O => \N__35497\,
            I => \N__35488\
        );

    \I__7924\ : Sp12to4
    port map (
            O => \N__35494\,
            I => \N__35483\
        );

    \I__7923\ : Sp12to4
    port map (
            O => \N__35491\,
            I => \N__35483\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__35488\,
            I => \N__35480\
        );

    \I__7921\ : Odrv12
    port map (
            O => \N__35483\,
            I => \POWERLED.func_state_RNI_1Z0Z_1\
        );

    \I__7920\ : Odrv12
    port map (
            O => \N__35480\,
            I => \POWERLED.func_state_RNI_1Z0Z_1\
        );

    \I__7919\ : InMux
    port map (
            O => \N__35475\,
            I => \N__35472\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__35472\,
            I => \N__35469\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__35469\,
            I => \N__35462\
        );

    \I__7916\ : InMux
    port map (
            O => \N__35468\,
            I => \N__35459\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__35467\,
            I => \N__35456\
        );

    \I__7914\ : InMux
    port map (
            O => \N__35466\,
            I => \N__35451\
        );

    \I__7913\ : InMux
    port map (
            O => \N__35465\,
            I => \N__35451\
        );

    \I__7912\ : Sp12to4
    port map (
            O => \N__35462\,
            I => \N__35448\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__35459\,
            I => \N__35445\
        );

    \I__7910\ : InMux
    port map (
            O => \N__35456\,
            I => \N__35442\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__35451\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_0\
        );

    \I__7908\ : Odrv12
    port map (
            O => \N__35448\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_0\
        );

    \I__7907\ : Odrv4
    port map (
            O => \N__35445\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_0\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__35442\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_0\
        );

    \I__7905\ : CascadeMux
    port map (
            O => \N__35433\,
            I => \N__35429\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__35432\,
            I => \N__35425\
        );

    \I__7903\ : InMux
    port map (
            O => \N__35429\,
            I => \N__35422\
        );

    \I__7902\ : InMux
    port map (
            O => \N__35428\,
            I => \N__35419\
        );

    \I__7901\ : InMux
    port map (
            O => \N__35425\,
            I => \N__35416\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__35422\,
            I => \N__35413\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__35419\,
            I => \N__35410\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35407\
        );

    \I__7897\ : Span4Mux_h
    port map (
            O => \N__35413\,
            I => \N__35404\
        );

    \I__7896\ : Span12Mux_v
    port map (
            O => \N__35410\,
            I => \N__35401\
        );

    \I__7895\ : Span4Mux_v
    port map (
            O => \N__35407\,
            I => \N__35398\
        );

    \I__7894\ : Odrv4
    port map (
            O => \N__35404\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_5\
        );

    \I__7893\ : Odrv12
    port map (
            O => \N__35401\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_5\
        );

    \I__7892\ : Odrv4
    port map (
            O => \N__35398\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_5\
        );

    \I__7891\ : InMux
    port map (
            O => \N__35391\,
            I => \N__35388\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__35388\,
            I => \N__35385\
        );

    \I__7889\ : Span4Mux_v
    port map (
            O => \N__35385\,
            I => \N__35382\
        );

    \I__7888\ : Span4Mux_h
    port map (
            O => \N__35382\,
            I => \N__35379\
        );

    \I__7887\ : Span4Mux_h
    port map (
            O => \N__35379\,
            I => \N__35376\
        );

    \I__7886\ : Odrv4
    port map (
            O => \N__35376\,
            I => \POWERLED.un1_clk_100khz_51_and_i_0_0\
        );

    \I__7885\ : InMux
    port map (
            O => \N__35373\,
            I => \N__35367\
        );

    \I__7884\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35367\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__35367\,
            I => \VPP_VDDQ.count_rst_11\
        );

    \I__7882\ : InMux
    port map (
            O => \N__35364\,
            I => \VPP_VDDQ.un4_count_1_cry_5\
        );

    \I__7881\ : CascadeMux
    port map (
            O => \N__35361\,
            I => \N__35358\
        );

    \I__7880\ : InMux
    port map (
            O => \N__35358\,
            I => \N__35354\
        );

    \I__7879\ : InMux
    port map (
            O => \N__35357\,
            I => \N__35351\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__35354\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__35351\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__7876\ : InMux
    port map (
            O => \N__35346\,
            I => \N__35340\
        );

    \I__7875\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35340\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__35340\,
            I => \VPP_VDDQ.count_rst_12\
        );

    \I__7873\ : InMux
    port map (
            O => \N__35337\,
            I => \VPP_VDDQ.un4_count_1_cry_6\
        );

    \I__7872\ : InMux
    port map (
            O => \N__35334\,
            I => \N__35330\
        );

    \I__7871\ : InMux
    port map (
            O => \N__35333\,
            I => \N__35327\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__35330\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__35327\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__7868\ : InMux
    port map (
            O => \N__35322\,
            I => \N__35316\
        );

    \I__7867\ : InMux
    port map (
            O => \N__35321\,
            I => \N__35316\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__35316\,
            I => \VPP_VDDQ.count_rst_13\
        );

    \I__7865\ : InMux
    port map (
            O => \N__35313\,
            I => \VPP_VDDQ.un4_count_1_cry_7\
        );

    \I__7864\ : InMux
    port map (
            O => \N__35310\,
            I => \N__35306\
        );

    \I__7863\ : CascadeMux
    port map (
            O => \N__35309\,
            I => \N__35303\
        );

    \I__7862\ : LocalMux
    port map (
            O => \N__35306\,
            I => \N__35300\
        );

    \I__7861\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35297\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__35300\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__7859\ : LocalMux
    port map (
            O => \N__35297\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__7858\ : InMux
    port map (
            O => \N__35292\,
            I => \N__35286\
        );

    \I__7857\ : InMux
    port map (
            O => \N__35291\,
            I => \N__35286\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__35286\,
            I => \N__35283\
        );

    \I__7855\ : Odrv12
    port map (
            O => \N__35283\,
            I => \VPP_VDDQ.count_rst_14\
        );

    \I__7854\ : InMux
    port map (
            O => \N__35280\,
            I => \bfn_12_6_0_\
        );

    \I__7853\ : InMux
    port map (
            O => \N__35277\,
            I => \N__35271\
        );

    \I__7852\ : InMux
    port map (
            O => \N__35276\,
            I => \N__35271\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__35271\,
            I => \N__35268\
        );

    \I__7850\ : Span4Mux_v
    port map (
            O => \N__35268\,
            I => \N__35265\
        );

    \I__7849\ : Odrv4
    port map (
            O => \N__35265\,
            I => \VPP_VDDQ.count_rst\
        );

    \I__7848\ : InMux
    port map (
            O => \N__35262\,
            I => \VPP_VDDQ.un4_count_1_cry_9\
        );

    \I__7847\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35245\
        );

    \I__7846\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35245\
        );

    \I__7845\ : InMux
    port map (
            O => \N__35257\,
            I => \N__35240\
        );

    \I__7844\ : InMux
    port map (
            O => \N__35256\,
            I => \N__35240\
        );

    \I__7843\ : InMux
    port map (
            O => \N__35255\,
            I => \N__35237\
        );

    \I__7842\ : InMux
    port map (
            O => \N__35254\,
            I => \N__35232\
        );

    \I__7841\ : InMux
    port map (
            O => \N__35253\,
            I => \N__35232\
        );

    \I__7840\ : InMux
    port map (
            O => \N__35252\,
            I => \N__35225\
        );

    \I__7839\ : InMux
    port map (
            O => \N__35251\,
            I => \N__35225\
        );

    \I__7838\ : InMux
    port map (
            O => \N__35250\,
            I => \N__35225\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__35245\,
            I => \N__35222\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__35240\,
            I => \N__35219\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__35237\,
            I => \VPP_VDDQ.un13_clk_100khz_i\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__35232\,
            I => \VPP_VDDQ.un13_clk_100khz_i\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__35225\,
            I => \VPP_VDDQ.un13_clk_100khz_i\
        );

    \I__7832\ : Odrv4
    port map (
            O => \N__35222\,
            I => \VPP_VDDQ.un13_clk_100khz_i\
        );

    \I__7831\ : Odrv12
    port map (
            O => \N__35219\,
            I => \VPP_VDDQ.un13_clk_100khz_i\
        );

    \I__7830\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35205\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__35205\,
            I => \N__35201\
        );

    \I__7828\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35198\
        );

    \I__7827\ : Odrv4
    port map (
            O => \N__35201\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__7826\ : LocalMux
    port map (
            O => \N__35198\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__7825\ : InMux
    port map (
            O => \N__35193\,
            I => \N__35187\
        );

    \I__7824\ : InMux
    port map (
            O => \N__35192\,
            I => \N__35187\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__35187\,
            I => \N__35184\
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__35184\,
            I => \VPP_VDDQ.count_rst_0\
        );

    \I__7821\ : InMux
    port map (
            O => \N__35181\,
            I => \VPP_VDDQ.un4_count_1_cry_10\
        );

    \I__7820\ : InMux
    port map (
            O => \N__35178\,
            I => \VPP_VDDQ.un4_count_1_cry_11\
        );

    \I__7819\ : CascadeMux
    port map (
            O => \N__35175\,
            I => \N__35172\
        );

    \I__7818\ : InMux
    port map (
            O => \N__35172\,
            I => \N__35168\
        );

    \I__7817\ : InMux
    port map (
            O => \N__35171\,
            I => \N__35165\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__35168\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__35165\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__7814\ : InMux
    port map (
            O => \N__35160\,
            I => \VPP_VDDQ.un4_count_1_cry_12\
        );

    \I__7813\ : InMux
    port map (
            O => \N__35157\,
            I => \N__35154\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__35154\,
            I => \VPP_VDDQ.count_4_9\
        );

    \I__7811\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35148\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__35148\,
            I => \VPP_VDDQ.count_4_11\
        );

    \I__7809\ : InMux
    port map (
            O => \N__35145\,
            I => \N__35138\
        );

    \I__7808\ : InMux
    port map (
            O => \N__35144\,
            I => \N__35138\
        );

    \I__7807\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35135\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__35138\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__35135\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__7804\ : CascadeMux
    port map (
            O => \N__35130\,
            I => \N__35124\
        );

    \I__7803\ : InMux
    port map (
            O => \N__35129\,
            I => \N__35116\
        );

    \I__7802\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35116\
        );

    \I__7801\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35116\
        );

    \I__7800\ : InMux
    port map (
            O => \N__35124\,
            I => \N__35113\
        );

    \I__7799\ : InMux
    port map (
            O => \N__35123\,
            I => \N__35110\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__35116\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__35113\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__35110\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__7795\ : InMux
    port map (
            O => \N__35103\,
            I => \VPP_VDDQ.un4_count_1_cry_1\
        );

    \I__7794\ : InMux
    port map (
            O => \N__35100\,
            I => \N__35096\
        );

    \I__7793\ : InMux
    port map (
            O => \N__35099\,
            I => \N__35093\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__35096\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__35093\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__7790\ : InMux
    port map (
            O => \N__35088\,
            I => \VPP_VDDQ.un4_count_1_cry_2_cZ0\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__35085\,
            I => \N__35082\
        );

    \I__7788\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35078\
        );

    \I__7787\ : InMux
    port map (
            O => \N__35081\,
            I => \N__35075\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__35078\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__7785\ : LocalMux
    port map (
            O => \N__35075\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__7784\ : InMux
    port map (
            O => \N__35070\,
            I => \VPP_VDDQ.un4_count_1_cry_3\
        );

    \I__7783\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35063\
        );

    \I__7782\ : InMux
    port map (
            O => \N__35066\,
            I => \N__35060\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__35063\,
            I => \N__35057\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__35060\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__7779\ : Odrv4
    port map (
            O => \N__35057\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__7778\ : InMux
    port map (
            O => \N__35052\,
            I => \N__35046\
        );

    \I__7777\ : InMux
    port map (
            O => \N__35051\,
            I => \N__35046\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__35046\,
            I => \VPP_VDDQ.count_rst_10\
        );

    \I__7775\ : InMux
    port map (
            O => \N__35043\,
            I => \VPP_VDDQ.un4_count_1_cry_4\
        );

    \I__7774\ : InMux
    port map (
            O => \N__35040\,
            I => \N__35034\
        );

    \I__7773\ : InMux
    port map (
            O => \N__35039\,
            I => \N__35034\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__35034\,
            I => \DSW_PWRGD.count_rst_0\
        );

    \I__7771\ : InMux
    port map (
            O => \N__35031\,
            I => \N__35028\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__35028\,
            I => \DSW_PWRGD.count_1_14\
        );

    \I__7769\ : InMux
    port map (
            O => \N__35025\,
            I => \N__35005\
        );

    \I__7768\ : SRMux
    port map (
            O => \N__35024\,
            I => \N__35005\
        );

    \I__7767\ : SRMux
    port map (
            O => \N__35023\,
            I => \N__35002\
        );

    \I__7766\ : InMux
    port map (
            O => \N__35022\,
            I => \N__34995\
        );

    \I__7765\ : InMux
    port map (
            O => \N__35021\,
            I => \N__34995\
        );

    \I__7764\ : InMux
    port map (
            O => \N__35020\,
            I => \N__34995\
        );

    \I__7763\ : InMux
    port map (
            O => \N__35019\,
            I => \N__34990\
        );

    \I__7762\ : InMux
    port map (
            O => \N__35018\,
            I => \N__34990\
        );

    \I__7761\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34985\
        );

    \I__7760\ : InMux
    port map (
            O => \N__35016\,
            I => \N__34985\
        );

    \I__7759\ : InMux
    port map (
            O => \N__35015\,
            I => \N__34982\
        );

    \I__7758\ : InMux
    port map (
            O => \N__35014\,
            I => \N__34975\
        );

    \I__7757\ : SRMux
    port map (
            O => \N__35013\,
            I => \N__34975\
        );

    \I__7756\ : SRMux
    port map (
            O => \N__35012\,
            I => \N__34972\
        );

    \I__7755\ : SRMux
    port map (
            O => \N__35011\,
            I => \N__34969\
        );

    \I__7754\ : CascadeMux
    port map (
            O => \N__35010\,
            I => \N__34960\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__35005\,
            I => \N__34952\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__35002\,
            I => \N__34949\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__34995\,
            I => \N__34940\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__34990\,
            I => \N__34940\
        );

    \I__7749\ : LocalMux
    port map (
            O => \N__34985\,
            I => \N__34940\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__34982\,
            I => \N__34940\
        );

    \I__7747\ : SRMux
    port map (
            O => \N__34981\,
            I => \N__34932\
        );

    \I__7746\ : InMux
    port map (
            O => \N__34980\,
            I => \N__34932\
        );

    \I__7745\ : LocalMux
    port map (
            O => \N__34975\,
            I => \N__34929\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__34972\,
            I => \N__34926\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__34969\,
            I => \N__34923\
        );

    \I__7742\ : SRMux
    port map (
            O => \N__34968\,
            I => \N__34920\
        );

    \I__7741\ : InMux
    port map (
            O => \N__34967\,
            I => \N__34915\
        );

    \I__7740\ : InMux
    port map (
            O => \N__34966\,
            I => \N__34915\
        );

    \I__7739\ : InMux
    port map (
            O => \N__34965\,
            I => \N__34908\
        );

    \I__7738\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34908\
        );

    \I__7737\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34908\
        );

    \I__7736\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34905\
        );

    \I__7735\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34900\
        );

    \I__7734\ : InMux
    port map (
            O => \N__34958\,
            I => \N__34900\
        );

    \I__7733\ : InMux
    port map (
            O => \N__34957\,
            I => \N__34893\
        );

    \I__7732\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34893\
        );

    \I__7731\ : InMux
    port map (
            O => \N__34955\,
            I => \N__34893\
        );

    \I__7730\ : Span4Mux_s1_h
    port map (
            O => \N__34952\,
            I => \N__34886\
        );

    \I__7729\ : Span4Mux_s1_h
    port map (
            O => \N__34949\,
            I => \N__34886\
        );

    \I__7728\ : Span4Mux_v
    port map (
            O => \N__34940\,
            I => \N__34886\
        );

    \I__7727\ : InMux
    port map (
            O => \N__34939\,
            I => \N__34881\
        );

    \I__7726\ : InMux
    port map (
            O => \N__34938\,
            I => \N__34881\
        );

    \I__7725\ : SRMux
    port map (
            O => \N__34937\,
            I => \N__34878\
        );

    \I__7724\ : LocalMux
    port map (
            O => \N__34932\,
            I => \N__34875\
        );

    \I__7723\ : Span4Mux_s1_v
    port map (
            O => \N__34929\,
            I => \N__34870\
        );

    \I__7722\ : Span4Mux_s3_h
    port map (
            O => \N__34926\,
            I => \N__34870\
        );

    \I__7721\ : Span4Mux_s3_h
    port map (
            O => \N__34923\,
            I => \N__34867\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__34920\,
            I => \N__34864\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__34915\,
            I => \N__34859\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__34908\,
            I => \N__34859\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__34905\,
            I => \N__34848\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__34900\,
            I => \N__34848\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__34893\,
            I => \N__34848\
        );

    \I__7714\ : Sp12to4
    port map (
            O => \N__34886\,
            I => \N__34848\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__34881\,
            I => \N__34848\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__34878\,
            I => \N__34841\
        );

    \I__7711\ : Span4Mux_v
    port map (
            O => \N__34875\,
            I => \N__34841\
        );

    \I__7710\ : Span4Mux_v
    port map (
            O => \N__34870\,
            I => \N__34841\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__34867\,
            I => \N__34838\
        );

    \I__7708\ : Span4Mux_s3_v
    port map (
            O => \N__34864\,
            I => \N__34833\
        );

    \I__7707\ : Span4Mux_s3_v
    port map (
            O => \N__34859\,
            I => \N__34833\
        );

    \I__7706\ : Span12Mux_s4_h
    port map (
            O => \N__34848\,
            I => \N__34830\
        );

    \I__7705\ : Odrv4
    port map (
            O => \N__34841\,
            I => \DSW_PWRGD.count_0_sqmuxa\
        );

    \I__7704\ : Odrv4
    port map (
            O => \N__34838\,
            I => \DSW_PWRGD.count_0_sqmuxa\
        );

    \I__7703\ : Odrv4
    port map (
            O => \N__34833\,
            I => \DSW_PWRGD.count_0_sqmuxa\
        );

    \I__7702\ : Odrv12
    port map (
            O => \N__34830\,
            I => \DSW_PWRGD.count_0_sqmuxa\
        );

    \I__7701\ : InMux
    port map (
            O => \N__34821\,
            I => \N__34815\
        );

    \I__7700\ : InMux
    port map (
            O => \N__34820\,
            I => \N__34815\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__34815\,
            I => \DSW_PWRGD.count_rst\
        );

    \I__7698\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34809\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__34809\,
            I => \DSW_PWRGD.count_1_15\
        );

    \I__7696\ : InMux
    port map (
            O => \N__34806\,
            I => \N__34803\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__34803\,
            I => \N__34800\
        );

    \I__7694\ : Odrv12
    port map (
            O => \N__34800\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__7693\ : InMux
    port map (
            O => \N__34797\,
            I => \N__34794\
        );

    \I__7692\ : LocalMux
    port map (
            O => \N__34794\,
            I => \N__34790\
        );

    \I__7691\ : InMux
    port map (
            O => \N__34793\,
            I => \N__34787\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__34790\,
            I => \DSW_PWRGD.count_i_0\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__34787\,
            I => \DSW_PWRGD.count_i_0\
        );

    \I__7688\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34778\
        );

    \I__7687\ : InMux
    port map (
            O => \N__34781\,
            I => \N__34775\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__34778\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__34775\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__7684\ : CascadeMux
    port map (
            O => \N__34770\,
            I => \DSW_PWRGD.countZ0Z_15_cascade_\
        );

    \I__7683\ : InMux
    port map (
            O => \N__34767\,
            I => \N__34763\
        );

    \I__7682\ : InMux
    port map (
            O => \N__34766\,
            I => \N__34760\
        );

    \I__7681\ : LocalMux
    port map (
            O => \N__34763\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__34760\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__7679\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34752\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34749\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__34749\,
            I => \N__34746\
        );

    \I__7676\ : Odrv4
    port map (
            O => \N__34746\,
            I => \DSW_PWRGD.un12_clk_100khz_9\
        );

    \I__7675\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34740\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__34740\,
            I => \N__34737\
        );

    \I__7673\ : Odrv4
    port map (
            O => \N__34737\,
            I => \DSW_PWRGD.count_1_1\
        );

    \I__7672\ : CEMux
    port map (
            O => \N__34734\,
            I => \N__34730\
        );

    \I__7671\ : CEMux
    port map (
            O => \N__34733\,
            I => \N__34719\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__34730\,
            I => \N__34715\
        );

    \I__7669\ : CEMux
    port map (
            O => \N__34729\,
            I => \N__34712\
        );

    \I__7668\ : CEMux
    port map (
            O => \N__34728\,
            I => \N__34709\
        );

    \I__7667\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34697\
        );

    \I__7666\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34697\
        );

    \I__7665\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34697\
        );

    \I__7664\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34697\
        );

    \I__7663\ : CEMux
    port map (
            O => \N__34723\,
            I => \N__34694\
        );

    \I__7662\ : CEMux
    port map (
            O => \N__34722\,
            I => \N__34691\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__34719\,
            I => \N__34671\
        );

    \I__7660\ : CEMux
    port map (
            O => \N__34718\,
            I => \N__34668\
        );

    \I__7659\ : Span4Mux_h
    port map (
            O => \N__34715\,
            I => \N__34665\
        );

    \I__7658\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34662\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34659\
        );

    \I__7656\ : InMux
    port map (
            O => \N__34708\,
            I => \N__34654\
        );

    \I__7655\ : InMux
    port map (
            O => \N__34707\,
            I => \N__34654\
        );

    \I__7654\ : InMux
    port map (
            O => \N__34706\,
            I => \N__34651\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34648\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__34694\,
            I => \N__34643\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__34691\,
            I => \N__34643\
        );

    \I__7650\ : InMux
    port map (
            O => \N__34690\,
            I => \N__34638\
        );

    \I__7649\ : CEMux
    port map (
            O => \N__34689\,
            I => \N__34638\
        );

    \I__7648\ : InMux
    port map (
            O => \N__34688\,
            I => \N__34633\
        );

    \I__7647\ : InMux
    port map (
            O => \N__34687\,
            I => \N__34633\
        );

    \I__7646\ : InMux
    port map (
            O => \N__34686\,
            I => \N__34626\
        );

    \I__7645\ : InMux
    port map (
            O => \N__34685\,
            I => \N__34626\
        );

    \I__7644\ : InMux
    port map (
            O => \N__34684\,
            I => \N__34626\
        );

    \I__7643\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34619\
        );

    \I__7642\ : InMux
    port map (
            O => \N__34682\,
            I => \N__34619\
        );

    \I__7641\ : InMux
    port map (
            O => \N__34681\,
            I => \N__34619\
        );

    \I__7640\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34612\
        );

    \I__7639\ : InMux
    port map (
            O => \N__34679\,
            I => \N__34612\
        );

    \I__7638\ : InMux
    port map (
            O => \N__34678\,
            I => \N__34612\
        );

    \I__7637\ : InMux
    port map (
            O => \N__34677\,
            I => \N__34603\
        );

    \I__7636\ : InMux
    port map (
            O => \N__34676\,
            I => \N__34603\
        );

    \I__7635\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34603\
        );

    \I__7634\ : InMux
    port map (
            O => \N__34674\,
            I => \N__34603\
        );

    \I__7633\ : Span4Mux_h
    port map (
            O => \N__34671\,
            I => \N__34600\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__34668\,
            I => \N__34597\
        );

    \I__7631\ : Span4Mux_s0_h
    port map (
            O => \N__34665\,
            I => \N__34594\
        );

    \I__7630\ : Span4Mux_s2_v
    port map (
            O => \N__34662\,
            I => \N__34583\
        );

    \I__7629\ : Span4Mux_h
    port map (
            O => \N__34659\,
            I => \N__34583\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__34654\,
            I => \N__34583\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__34651\,
            I => \N__34583\
        );

    \I__7626\ : Span4Mux_s2_v
    port map (
            O => \N__34648\,
            I => \N__34583\
        );

    \I__7625\ : Span4Mux_s2_v
    port map (
            O => \N__34643\,
            I => \N__34578\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__34638\,
            I => \N__34578\
        );

    \I__7623\ : LocalMux
    port map (
            O => \N__34633\,
            I => \N__34567\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__34626\,
            I => \N__34567\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__34619\,
            I => \N__34567\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__34612\,
            I => \N__34567\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__34603\,
            I => \N__34567\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__34600\,
            I => \N__34564\
        );

    \I__7617\ : Span4Mux_s3_v
    port map (
            O => \N__34597\,
            I => \N__34559\
        );

    \I__7616\ : Span4Mux_h
    port map (
            O => \N__34594\,
            I => \N__34559\
        );

    \I__7615\ : Span4Mux_v
    port map (
            O => \N__34583\,
            I => \N__34556\
        );

    \I__7614\ : Span4Mux_s0_h
    port map (
            O => \N__34578\,
            I => \N__34551\
        );

    \I__7613\ : Span4Mux_s2_v
    port map (
            O => \N__34567\,
            I => \N__34551\
        );

    \I__7612\ : Odrv4
    port map (
            O => \N__34564\,
            I => \DSW_PWRGD.curr_state_RNI57NNZ0Z_0\
        );

    \I__7611\ : Odrv4
    port map (
            O => \N__34559\,
            I => \DSW_PWRGD.curr_state_RNI57NNZ0Z_0\
        );

    \I__7610\ : Odrv4
    port map (
            O => \N__34556\,
            I => \DSW_PWRGD.curr_state_RNI57NNZ0Z_0\
        );

    \I__7609\ : Odrv4
    port map (
            O => \N__34551\,
            I => \DSW_PWRGD.curr_state_RNI57NNZ0Z_0\
        );

    \I__7608\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34539\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__7606\ : Span4Mux_h
    port map (
            O => \N__34536\,
            I => \N__34532\
        );

    \I__7605\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34529\
        );

    \I__7604\ : Odrv4
    port map (
            O => \N__34532\,
            I => \DSW_PWRGD.count_rst_13\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__34529\,
            I => \DSW_PWRGD.count_rst_13\
        );

    \I__7602\ : CascadeMux
    port map (
            O => \N__34524\,
            I => \N__34521\
        );

    \I__7601\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34518\
        );

    \I__7600\ : LocalMux
    port map (
            O => \N__34518\,
            I => \N__34514\
        );

    \I__7599\ : InMux
    port map (
            O => \N__34517\,
            I => \N__34511\
        );

    \I__7598\ : Odrv4
    port map (
            O => \N__34514\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__34511\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__7596\ : InMux
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__34503\,
            I => \VPP_VDDQ.count_4_7\
        );

    \I__7594\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34497\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__34497\,
            I => \VPP_VDDQ.count_4_8\
        );

    \I__7592\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34491\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__34491\,
            I => \DSW_PWRGD.count_1_12\
        );

    \I__7590\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34482\
        );

    \I__7589\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34482\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__34482\,
            I => \DSW_PWRGD.count_rst_2\
        );

    \I__7587\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34476\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__34476\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__7585\ : InMux
    port map (
            O => \N__34473\,
            I => \N__34464\
        );

    \I__7584\ : InMux
    port map (
            O => \N__34472\,
            I => \N__34464\
        );

    \I__7583\ : InMux
    port map (
            O => \N__34471\,
            I => \N__34464\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__34464\,
            I => \DSW_PWRGD.count_rst_5\
        );

    \I__7581\ : InMux
    port map (
            O => \N__34461\,
            I => \N__34455\
        );

    \I__7580\ : InMux
    port map (
            O => \N__34460\,
            I => \N__34455\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__34455\,
            I => \DSW_PWRGD.count_1_9\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__34452\,
            I => \DSW_PWRGD.countZ0Z_12_cascade_\
        );

    \I__7577\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34446\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__34446\,
            I => \N__34443\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__34443\,
            I => \N__34440\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__34440\,
            I => \DSW_PWRGD.un12_clk_100khz_1\
        );

    \I__7573\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34434\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__34434\,
            I => \DSW_PWRGD.un2_count_1_axb_4\
        );

    \I__7571\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34422\
        );

    \I__7570\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34422\
        );

    \I__7569\ : InMux
    port map (
            O => \N__34429\,
            I => \N__34422\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__34422\,
            I => \DSW_PWRGD.count_rst_10\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__34419\,
            I => \N__34416\
        );

    \I__7566\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34410\
        );

    \I__7565\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34410\
        );

    \I__7564\ : LocalMux
    port map (
            O => \N__34410\,
            I => \DSW_PWRGD.count_1_4\
        );

    \I__7563\ : InMux
    port map (
            O => \N__34407\,
            I => \N__34403\
        );

    \I__7562\ : InMux
    port map (
            O => \N__34406\,
            I => \N__34400\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34395\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__34400\,
            I => \N__34395\
        );

    \I__7559\ : Span4Mux_s2_v
    port map (
            O => \N__34395\,
            I => \N__34392\
        );

    \I__7558\ : Span4Mux_v
    port map (
            O => \N__34392\,
            I => \N__34389\
        );

    \I__7557\ : Odrv4
    port map (
            O => \N__34389\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__7556\ : CascadeMux
    port map (
            O => \N__34386\,
            I => \N__34383\
        );

    \I__7555\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34380\
        );

    \I__7554\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34377\
        );

    \I__7553\ : Span4Mux_h
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__34374\,
            I => \DSW_PWRGD.un12_clk_100khz_0\
        );

    \I__7551\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34365\
        );

    \I__7550\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34365\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__34365\,
            I => \DSW_PWRGD.count_rst_1\
        );

    \I__7548\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34359\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__34359\,
            I => \DSW_PWRGD.count_1_13\
        );

    \I__7546\ : CascadeMux
    port map (
            O => \N__34356\,
            I => \DSW_PWRGD.count_rst_14_cascade_\
        );

    \I__7545\ : CascadeMux
    port map (
            O => \N__34353\,
            I => \DSW_PWRGD.count_i_0_cascade_\
        );

    \I__7544\ : InMux
    port map (
            O => \N__34350\,
            I => \N__34346\
        );

    \I__7543\ : InMux
    port map (
            O => \N__34349\,
            I => \N__34343\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__34346\,
            I => \DSW_PWRGD.count_1_0\
        );

    \I__7541\ : LocalMux
    port map (
            O => \N__34343\,
            I => \DSW_PWRGD.count_1_0\
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__34338\,
            I => \DSW_PWRGD.count_rst_3_cascade_\
        );

    \I__7539\ : CascadeMux
    port map (
            O => \N__34335\,
            I => \N__34332\
        );

    \I__7538\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34328\
        );

    \I__7537\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34325\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__34328\,
            I => \N__34322\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__34325\,
            I => \DSW_PWRGD.un2_count_1_axb_11\
        );

    \I__7534\ : Odrv4
    port map (
            O => \N__34322\,
            I => \DSW_PWRGD.un2_count_1_axb_11\
        );

    \I__7533\ : CascadeMux
    port map (
            O => \N__34317\,
            I => \N__34309\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__34316\,
            I => \N__34306\
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__34315\,
            I => \N__34299\
        );

    \I__7530\ : InMux
    port map (
            O => \N__34314\,
            I => \N__34289\
        );

    \I__7529\ : InMux
    port map (
            O => \N__34313\,
            I => \N__34289\
        );

    \I__7528\ : InMux
    port map (
            O => \N__34312\,
            I => \N__34289\
        );

    \I__7527\ : InMux
    port map (
            O => \N__34309\,
            I => \N__34284\
        );

    \I__7526\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34284\
        );

    \I__7525\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34275\
        );

    \I__7524\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34275\
        );

    \I__7523\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34275\
        );

    \I__7522\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34275\
        );

    \I__7521\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34260\
        );

    \I__7520\ : InMux
    port map (
            O => \N__34298\,
            I => \N__34260\
        );

    \I__7519\ : InMux
    port map (
            O => \N__34297\,
            I => \N__34260\
        );

    \I__7518\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34260\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__34289\,
            I => \N__34253\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__34284\,
            I => \N__34253\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__34275\,
            I => \N__34253\
        );

    \I__7514\ : InMux
    port map (
            O => \N__34274\,
            I => \N__34244\
        );

    \I__7513\ : InMux
    port map (
            O => \N__34273\,
            I => \N__34244\
        );

    \I__7512\ : InMux
    port map (
            O => \N__34272\,
            I => \N__34244\
        );

    \I__7511\ : InMux
    port map (
            O => \N__34271\,
            I => \N__34244\
        );

    \I__7510\ : InMux
    port map (
            O => \N__34270\,
            I => \N__34239\
        );

    \I__7509\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34239\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__34260\,
            I => \N__34234\
        );

    \I__7507\ : Span4Mux_s2_h
    port map (
            O => \N__34253\,
            I => \N__34234\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__34244\,
            I => \N__34231\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__34239\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__7504\ : Odrv4
    port map (
            O => \N__34234\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__7503\ : Odrv4
    port map (
            O => \N__34231\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__7502\ : CascadeMux
    port map (
            O => \N__34224\,
            I => \DSW_PWRGD.un2_count_1_axb_11_cascade_\
        );

    \I__7501\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34215\
        );

    \I__7500\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34215\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__34215\,
            I => \N__34212\
        );

    \I__7498\ : Odrv4
    port map (
            O => \N__34212\,
            I => \DSW_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__7497\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34206\
        );

    \I__7496\ : LocalMux
    port map (
            O => \N__34206\,
            I => \DSW_PWRGD.count_rst_3\
        );

    \I__7495\ : InMux
    port map (
            O => \N__34203\,
            I => \N__34197\
        );

    \I__7494\ : InMux
    port map (
            O => \N__34202\,
            I => \N__34197\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__34197\,
            I => \DSW_PWRGD.count_1_11\
        );

    \I__7492\ : InMux
    port map (
            O => \N__34194\,
            I => \N__34191\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__34191\,
            I => \N__34188\
        );

    \I__7490\ : Span4Mux_v
    port map (
            O => \N__34188\,
            I => \N__34185\
        );

    \I__7489\ : Odrv4
    port map (
            O => \N__34185\,
            I => \DSW_PWRGD.un12_clk_100khz_7\
        );

    \I__7488\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34179\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__34179\,
            I => \DSW_PWRGD.un2_count_1_axb_9\
        );

    \I__7486\ : InMux
    port map (
            O => \N__34176\,
            I => \N__34173\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__34173\,
            I => \N__34170\
        );

    \I__7484\ : Odrv4
    port map (
            O => \N__34170\,
            I => \HDA_STRAP.un2_count_1_axb_15\
        );

    \I__7483\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34161\
        );

    \I__7482\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34161\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__34161\,
            I => \N__34158\
        );

    \I__7480\ : Odrv12
    port map (
            O => \N__34158\,
            I => \HDA_STRAP.count_1_6\
        );

    \I__7479\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34152\
        );

    \I__7478\ : LocalMux
    port map (
            O => \N__34152\,
            I => \HDA_STRAP.count_3_6\
        );

    \I__7477\ : InMux
    port map (
            O => \N__34149\,
            I => \N__34146\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__34146\,
            I => \N__34143\
        );

    \I__7475\ : Odrv4
    port map (
            O => \N__34143\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__7474\ : InMux
    port map (
            O => \N__34140\,
            I => \N__34134\
        );

    \I__7473\ : InMux
    port map (
            O => \N__34139\,
            I => \N__34134\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__34134\,
            I => \HDA_STRAP.count_3_15\
        );

    \I__7471\ : InMux
    port map (
            O => \N__34131\,
            I => \N__34122\
        );

    \I__7470\ : InMux
    port map (
            O => \N__34130\,
            I => \N__34122\
        );

    \I__7469\ : InMux
    port map (
            O => \N__34129\,
            I => \N__34122\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__34122\,
            I => \N__34119\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__34119\,
            I => \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0\
        );

    \I__7466\ : CascadeMux
    port map (
            O => \N__34116\,
            I => \HDA_STRAP.countZ0Z_6_cascade_\
        );

    \I__7465\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34110\
        );

    \I__7464\ : LocalMux
    port map (
            O => \N__34110\,
            I => \N__34107\
        );

    \I__7463\ : Odrv4
    port map (
            O => \N__34107\,
            I => \HDA_STRAP.un2_count_1_axb_16\
        );

    \I__7462\ : InMux
    port map (
            O => \N__34104\,
            I => \N__34098\
        );

    \I__7461\ : InMux
    port map (
            O => \N__34103\,
            I => \N__34098\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__34098\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__7459\ : CascadeMux
    port map (
            O => \N__34095\,
            I => \N__34091\
        );

    \I__7458\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34087\
        );

    \I__7457\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34082\
        );

    \I__7456\ : InMux
    port map (
            O => \N__34090\,
            I => \N__34082\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__34087\,
            I => \N__34077\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__34082\,
            I => \N__34077\
        );

    \I__7453\ : Odrv4
    port map (
            O => \N__34077\,
            I => \HDA_STRAP.count_1_16\
        );

    \I__7452\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34070\
        );

    \I__7451\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34067\
        );

    \I__7450\ : LocalMux
    port map (
            O => \N__34070\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__34067\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__7448\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34059\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__34059\,
            I => \DSW_PWRGD.un2_count_1_axb_0\
        );

    \I__7446\ : InMux
    port map (
            O => \N__34056\,
            I => \N__34053\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__34053\,
            I => \DSW_PWRGD.count_rst_14\
        );

    \I__7444\ : InMux
    port map (
            O => \N__34050\,
            I => \HDA_STRAP.un2_count_1_cry_10\
        );

    \I__7443\ : InMux
    port map (
            O => \N__34047\,
            I => \HDA_STRAP.un2_count_1_cry_11\
        );

    \I__7442\ : InMux
    port map (
            O => \N__34044\,
            I => \HDA_STRAP.un2_count_1_cry_12\
        );

    \I__7441\ : InMux
    port map (
            O => \N__34041\,
            I => \N__34037\
        );

    \I__7440\ : InMux
    port map (
            O => \N__34040\,
            I => \N__34034\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__34037\,
            I => \N__34031\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__34034\,
            I => \N__34026\
        );

    \I__7437\ : Span12Mux_s10_h
    port map (
            O => \N__34031\,
            I => \N__34026\
        );

    \I__7436\ : Odrv12
    port map (
            O => \N__34026\,
            I => \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3\
        );

    \I__7435\ : InMux
    port map (
            O => \N__34023\,
            I => \HDA_STRAP.un2_count_1_cry_13\
        );

    \I__7434\ : InMux
    port map (
            O => \N__34020\,
            I => \HDA_STRAP.un2_count_1_cry_14\
        );

    \I__7433\ : InMux
    port map (
            O => \N__34017\,
            I => \HDA_STRAP.un2_count_1_cry_15\
        );

    \I__7432\ : InMux
    port map (
            O => \N__34014\,
            I => \bfn_11_15_0_\
        );

    \I__7431\ : InMux
    port map (
            O => \N__34011\,
            I => \N__34008\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__7429\ : Odrv12
    port map (
            O => \N__34005\,
            I => \HDA_STRAP.count_0_17\
        );

    \I__7428\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33999\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__33999\,
            I => \N__33995\
        );

    \I__7426\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33992\
        );

    \I__7425\ : Odrv4
    port map (
            O => \N__33995\,
            I => \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__33992\,
            I => \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\
        );

    \I__7423\ : InMux
    port map (
            O => \N__33987\,
            I => \HDA_STRAP.un2_count_1_cry_1\
        );

    \I__7422\ : InMux
    port map (
            O => \N__33984\,
            I => \HDA_STRAP.un2_count_1_cry_2\
        );

    \I__7421\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33978\
        );

    \I__7420\ : LocalMux
    port map (
            O => \N__33978\,
            I => \N__33975\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__33975\,
            I => \N__33971\
        );

    \I__7418\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33968\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__33971\,
            I => \N__33965\
        );

    \I__7416\ : LocalMux
    port map (
            O => \N__33968\,
            I => \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__33965\,
            I => \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\
        );

    \I__7414\ : InMux
    port map (
            O => \N__33960\,
            I => \HDA_STRAP.un2_count_1_cry_3\
        );

    \I__7413\ : InMux
    port map (
            O => \N__33957\,
            I => \HDA_STRAP.un2_count_1_cry_4\
        );

    \I__7412\ : InMux
    port map (
            O => \N__33954\,
            I => \HDA_STRAP.un2_count_1_cry_5_cZ0\
        );

    \I__7411\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33948\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__33948\,
            I => \N__33944\
        );

    \I__7409\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33941\
        );

    \I__7408\ : Span12Mux_s10_h
    port map (
            O => \N__33944\,
            I => \N__33938\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__33941\,
            I => \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\
        );

    \I__7406\ : Odrv12
    port map (
            O => \N__33938\,
            I => \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\
        );

    \I__7405\ : InMux
    port map (
            O => \N__33933\,
            I => \HDA_STRAP.un2_count_1_cry_6\
        );

    \I__7404\ : InMux
    port map (
            O => \N__33930\,
            I => \HDA_STRAP.un2_count_1_cry_7\
        );

    \I__7403\ : InMux
    port map (
            O => \N__33927\,
            I => \bfn_11_14_0_\
        );

    \I__7402\ : InMux
    port map (
            O => \N__33924\,
            I => \HDA_STRAP.un2_count_1_cry_9\
        );

    \I__7401\ : CascadeMux
    port map (
            O => \N__33921\,
            I => \N__33918\
        );

    \I__7400\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33915\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__7398\ : Span4Mux_v
    port map (
            O => \N__33912\,
            I => \N__33909\
        );

    \I__7397\ : Odrv4
    port map (
            O => \N__33909\,
            I => \POWERLED.un85_clk_100khz_2\
        );

    \I__7396\ : InMux
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__7395\ : LocalMux
    port map (
            O => \N__33903\,
            I => \N__33899\
        );

    \I__7394\ : InMux
    port map (
            O => \N__33902\,
            I => \N__33896\
        );

    \I__7393\ : Span4Mux_v
    port map (
            O => \N__33899\,
            I => \N__33893\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__33896\,
            I => \N__33890\
        );

    \I__7391\ : Odrv4
    port map (
            O => \N__33893\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__33890\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__7389\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33882\
        );

    \I__7388\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33879\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__33879\,
            I => \N__33876\
        );

    \I__7386\ : Odrv12
    port map (
            O => \N__33876\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__7385\ : InMux
    port map (
            O => \N__33873\,
            I => \N__33870\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__33870\,
            I => \N__33867\
        );

    \I__7383\ : Span4Mux_v
    port map (
            O => \N__33867\,
            I => \N__33864\
        );

    \I__7382\ : Span4Mux_v
    port map (
            O => \N__33864\,
            I => \N__33861\
        );

    \I__7381\ : Odrv4
    port map (
            O => \N__33861\,
            I => \HDA_STRAP.count_3_14\
        );

    \I__7380\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33855\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__33855\,
            I => \N__33852\
        );

    \I__7378\ : Span4Mux_v
    port map (
            O => \N__33852\,
            I => \N__33849\
        );

    \I__7377\ : Span4Mux_v
    port map (
            O => \N__33849\,
            I => \N__33846\
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__33846\,
            I => \HDA_STRAP.count_3_4\
        );

    \I__7375\ : InMux
    port map (
            O => \N__33843\,
            I => \N__33840\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__7373\ : Span4Mux_h
    port map (
            O => \N__33837\,
            I => \N__33834\
        );

    \I__7372\ : Span4Mux_v
    port map (
            O => \N__33834\,
            I => \N__33831\
        );

    \I__7371\ : Odrv4
    port map (
            O => \N__33831\,
            I => \HDA_STRAP.count_3_7\
        );

    \I__7370\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33824\
        );

    \I__7369\ : InMux
    port map (
            O => \N__33827\,
            I => \N__33821\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__33824\,
            I => \N__33818\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__33821\,
            I => \N__33815\
        );

    \I__7366\ : Span4Mux_v
    port map (
            O => \N__33818\,
            I => \N__33812\
        );

    \I__7365\ : Span4Mux_v
    port map (
            O => \N__33815\,
            I => \N__33809\
        );

    \I__7364\ : Odrv4
    port map (
            O => \N__33812\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__7363\ : Odrv4
    port map (
            O => \N__33809\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__7362\ : CascadeMux
    port map (
            O => \N__33804\,
            I => \N__33801\
        );

    \I__7361\ : InMux
    port map (
            O => \N__33801\,
            I => \N__33798\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__33798\,
            I => \N__33795\
        );

    \I__7359\ : Span4Mux_v
    port map (
            O => \N__33795\,
            I => \N__33792\
        );

    \I__7358\ : Odrv4
    port map (
            O => \N__33792\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__7357\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33786\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__33786\,
            I => \N__33782\
        );

    \I__7355\ : InMux
    port map (
            O => \N__33785\,
            I => \N__33779\
        );

    \I__7354\ : Span4Mux_s1_h
    port map (
            O => \N__33782\,
            I => \N__33774\
        );

    \I__7353\ : LocalMux
    port map (
            O => \N__33779\,
            I => \N__33774\
        );

    \I__7352\ : Span4Mux_v
    port map (
            O => \N__33774\,
            I => \N__33771\
        );

    \I__7351\ : Odrv4
    port map (
            O => \N__33771\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__7350\ : InMux
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33761\
        );

    \I__7348\ : InMux
    port map (
            O => \N__33764\,
            I => \N__33758\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__33761\,
            I => \N__33753\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__33758\,
            I => \N__33753\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__7344\ : Span4Mux_v
    port map (
            O => \N__33750\,
            I => \N__33747\
        );

    \I__7343\ : Odrv4
    port map (
            O => \N__33747\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__7342\ : InMux
    port map (
            O => \N__33744\,
            I => \N__33741\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__33741\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__7340\ : CascadeMux
    port map (
            O => \N__33738\,
            I => \N__33735\
        );

    \I__7339\ : InMux
    port map (
            O => \N__33735\,
            I => \N__33732\
        );

    \I__7338\ : LocalMux
    port map (
            O => \N__33732\,
            I => \N__33729\
        );

    \I__7337\ : Span4Mux_h
    port map (
            O => \N__33729\,
            I => \N__33726\
        );

    \I__7336\ : Span4Mux_s1_h
    port map (
            O => \N__33726\,
            I => \N__33723\
        );

    \I__7335\ : Odrv4
    port map (
            O => \N__33723\,
            I => \POWERLED.un85_clk_100khz_4\
        );

    \I__7334\ : InMux
    port map (
            O => \N__33720\,
            I => \N__33717\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__33717\,
            I => \N__33713\
        );

    \I__7332\ : CascadeMux
    port map (
            O => \N__33716\,
            I => \N__33709\
        );

    \I__7331\ : Span4Mux_h
    port map (
            O => \N__33713\,
            I => \N__33704\
        );

    \I__7330\ : InMux
    port map (
            O => \N__33712\,
            I => \N__33697\
        );

    \I__7329\ : InMux
    port map (
            O => \N__33709\,
            I => \N__33697\
        );

    \I__7328\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33697\
        );

    \I__7327\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33694\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__33704\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__33697\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__33694\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__7323\ : CascadeMux
    port map (
            O => \N__33687\,
            I => \N__33684\
        );

    \I__7322\ : InMux
    port map (
            O => \N__33684\,
            I => \N__33681\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__33681\,
            I => \N__33678\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__33678\,
            I => \POWERLED.mult1_un96_sum_i_8\
        );

    \I__7319\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33672\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33669\
        );

    \I__7317\ : Span4Mux_v
    port map (
            O => \N__33669\,
            I => \N__33666\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__33666\,
            I => \POWERLED.un85_clk_100khz_1\
        );

    \I__7315\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33660\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__33660\,
            I => \N__33656\
        );

    \I__7313\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33653\
        );

    \I__7312\ : Span4Mux_v
    port map (
            O => \N__33656\,
            I => \N__33648\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__33653\,
            I => \N__33648\
        );

    \I__7310\ : Span4Mux_h
    port map (
            O => \N__33648\,
            I => \N__33645\
        );

    \I__7309\ : Odrv4
    port map (
            O => \N__33645\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__7308\ : InMux
    port map (
            O => \N__33642\,
            I => \N__33639\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__33639\,
            I => \N__33636\
        );

    \I__7306\ : Odrv4
    port map (
            O => \N__33636\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__7305\ : InMux
    port map (
            O => \N__33633\,
            I => \N__33630\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__33630\,
            I => \N__33627\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__33627\,
            I => \N__33623\
        );

    \I__7302\ : InMux
    port map (
            O => \N__33626\,
            I => \N__33619\
        );

    \I__7301\ : Span4Mux_v
    port map (
            O => \N__33623\,
            I => \N__33616\
        );

    \I__7300\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33613\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__33619\,
            I => \N__33610\
        );

    \I__7298\ : Odrv4
    port map (
            O => \N__33616\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__33613\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7296\ : Odrv4
    port map (
            O => \N__33610\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7295\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33597\
        );

    \I__7294\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33597\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__33597\,
            I => \N__33594\
        );

    \I__7292\ : Span4Mux_h
    port map (
            O => \N__33594\,
            I => \N__33591\
        );

    \I__7291\ : Span4Mux_v
    port map (
            O => \N__33591\,
            I => \N__33588\
        );

    \I__7290\ : Odrv4
    port map (
            O => \N__33588\,
            I => \VPP_VDDQ.m4_0_a2\
        );

    \I__7289\ : CascadeMux
    port map (
            O => \N__33585\,
            I => \N__33582\
        );

    \I__7288\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33579\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__33579\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__7286\ : InMux
    port map (
            O => \N__33576\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__7285\ : InMux
    port map (
            O => \N__33573\,
            I => \N__33570\
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__33570\,
            I => \POWERLED.mult1_un131_sum_axb_4_l_fx\
        );

    \I__7283\ : CascadeMux
    port map (
            O => \N__33567\,
            I => \N__33564\
        );

    \I__7282\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33561\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__33561\,
            I => \N__33557\
        );

    \I__7280\ : InMux
    port map (
            O => \N__33560\,
            I => \N__33554\
        );

    \I__7279\ : Span4Mux_v
    port map (
            O => \N__33557\,
            I => \N__33551\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__33554\,
            I => \N__33548\
        );

    \I__7277\ : Odrv4
    port map (
            O => \N__33551\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__7276\ : Odrv4
    port map (
            O => \N__33548\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__7275\ : InMux
    port map (
            O => \N__33543\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__7274\ : CascadeMux
    port map (
            O => \N__33540\,
            I => \N__33537\
        );

    \I__7273\ : InMux
    port map (
            O => \N__33537\,
            I => \N__33534\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__7271\ : Span4Mux_v
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__7270\ : Odrv4
    port map (
            O => \N__33528\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__7269\ : InMux
    port map (
            O => \N__33525\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__7268\ : InMux
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__33519\,
            I => \N__33516\
        );

    \I__7266\ : Span4Mux_v
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__33513\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__7264\ : CascadeMux
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__7263\ : InMux
    port map (
            O => \N__33507\,
            I => \N__33501\
        );

    \I__7262\ : InMux
    port map (
            O => \N__33506\,
            I => \N__33501\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__33501\,
            I => \N__33494\
        );

    \I__7260\ : InMux
    port map (
            O => \N__33500\,
            I => \N__33485\
        );

    \I__7259\ : InMux
    port map (
            O => \N__33499\,
            I => \N__33485\
        );

    \I__7258\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33485\
        );

    \I__7257\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33485\
        );

    \I__7256\ : Span4Mux_v
    port map (
            O => \N__33494\,
            I => \N__33479\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__33485\,
            I => \N__33479\
        );

    \I__7254\ : InMux
    port map (
            O => \N__33484\,
            I => \N__33476\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__33479\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__33476\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__7251\ : InMux
    port map (
            O => \N__33471\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__7250\ : InMux
    port map (
            O => \N__33468\,
            I => \N__33465\
        );

    \I__7249\ : LocalMux
    port map (
            O => \N__33465\,
            I => \POWERLED.mult1_un131_sum_axb_7_l_fx\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__33462\,
            I => \N__33459\
        );

    \I__7247\ : InMux
    port map (
            O => \N__33459\,
            I => \N__33456\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__33456\,
            I => \N__33452\
        );

    \I__7245\ : InMux
    port map (
            O => \N__33455\,
            I => \N__33449\
        );

    \I__7244\ : Span4Mux_v
    port map (
            O => \N__33452\,
            I => \N__33446\
        );

    \I__7243\ : LocalMux
    port map (
            O => \N__33449\,
            I => \N__33443\
        );

    \I__7242\ : Odrv4
    port map (
            O => \N__33446\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__7241\ : Odrv12
    port map (
            O => \N__33443\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__7240\ : InMux
    port map (
            O => \N__33438\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__7239\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33432\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__33432\,
            I => \N__33429\
        );

    \I__7237\ : Span4Mux_v
    port map (
            O => \N__33429\,
            I => \N__33426\
        );

    \I__7236\ : Odrv4
    port map (
            O => \N__33426\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__7235\ : InMux
    port map (
            O => \N__33423\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__7234\ : CascadeMux
    port map (
            O => \N__33420\,
            I => \POWERLED.mult1_un131_sum_s_8_cascade_\
        );

    \I__7233\ : CascadeMux
    port map (
            O => \N__33417\,
            I => \N__33414\
        );

    \I__7232\ : InMux
    port map (
            O => \N__33414\,
            I => \N__33411\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__33411\,
            I => \N__33408\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__7229\ : Odrv4
    port map (
            O => \N__33405\,
            I => \POWERLED.un85_clk_100khz_5\
        );

    \I__7228\ : CascadeMux
    port map (
            O => \N__33402\,
            I => \VPP_VDDQ.curr_stateZ0Z_1_cascade_\
        );

    \I__7227\ : CascadeMux
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__7226\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__33393\,
            I => \VPP_VDDQ.curr_state_0_1\
        );

    \I__7224\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33383\
        );

    \I__7223\ : CascadeMux
    port map (
            O => \N__33389\,
            I => \N__33371\
        );

    \I__7222\ : CascadeMux
    port map (
            O => \N__33388\,
            I => \N__33364\
        );

    \I__7221\ : InMux
    port map (
            O => \N__33387\,
            I => \N__33355\
        );

    \I__7220\ : InMux
    port map (
            O => \N__33386\,
            I => \N__33352\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__33383\,
            I => \N__33349\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__33382\,
            I => \N__33345\
        );

    \I__7217\ : CascadeMux
    port map (
            O => \N__33381\,
            I => \N__33342\
        );

    \I__7216\ : InMux
    port map (
            O => \N__33380\,
            I => \N__33339\
        );

    \I__7215\ : InMux
    port map (
            O => \N__33379\,
            I => \N__33332\
        );

    \I__7214\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33332\
        );

    \I__7213\ : InMux
    port map (
            O => \N__33377\,
            I => \N__33332\
        );

    \I__7212\ : CascadeMux
    port map (
            O => \N__33376\,
            I => \N__33326\
        );

    \I__7211\ : InMux
    port map (
            O => \N__33375\,
            I => \N__33317\
        );

    \I__7210\ : InMux
    port map (
            O => \N__33374\,
            I => \N__33317\
        );

    \I__7209\ : InMux
    port map (
            O => \N__33371\,
            I => \N__33303\
        );

    \I__7208\ : InMux
    port map (
            O => \N__33370\,
            I => \N__33303\
        );

    \I__7207\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33303\
        );

    \I__7206\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33297\
        );

    \I__7205\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33294\
        );

    \I__7204\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33281\
        );

    \I__7203\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33276\
        );

    \I__7202\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33276\
        );

    \I__7201\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33271\
        );

    \I__7200\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33271\
        );

    \I__7199\ : CascadeMux
    port map (
            O => \N__33359\,
            I => \N__33268\
        );

    \I__7198\ : CascadeMux
    port map (
            O => \N__33358\,
            I => \N__33265\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__33355\,
            I => \N__33260\
        );

    \I__7196\ : LocalMux
    port map (
            O => \N__33352\,
            I => \N__33257\
        );

    \I__7195\ : Span4Mux_v
    port map (
            O => \N__33349\,
            I => \N__33254\
        );

    \I__7194\ : InMux
    port map (
            O => \N__33348\,
            I => \N__33251\
        );

    \I__7193\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33246\
        );

    \I__7192\ : InMux
    port map (
            O => \N__33342\,
            I => \N__33246\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__33339\,
            I => \N__33241\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33241\
        );

    \I__7189\ : InMux
    port map (
            O => \N__33331\,
            I => \N__33234\
        );

    \I__7188\ : InMux
    port map (
            O => \N__33330\,
            I => \N__33234\
        );

    \I__7187\ : InMux
    port map (
            O => \N__33329\,
            I => \N__33234\
        );

    \I__7186\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33225\
        );

    \I__7185\ : InMux
    port map (
            O => \N__33325\,
            I => \N__33225\
        );

    \I__7184\ : InMux
    port map (
            O => \N__33324\,
            I => \N__33225\
        );

    \I__7183\ : InMux
    port map (
            O => \N__33323\,
            I => \N__33225\
        );

    \I__7182\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33222\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__33317\,
            I => \N__33219\
        );

    \I__7180\ : InMux
    port map (
            O => \N__33316\,
            I => \N__33214\
        );

    \I__7179\ : InMux
    port map (
            O => \N__33315\,
            I => \N__33214\
        );

    \I__7178\ : InMux
    port map (
            O => \N__33314\,
            I => \N__33211\
        );

    \I__7177\ : InMux
    port map (
            O => \N__33313\,
            I => \N__33202\
        );

    \I__7176\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33202\
        );

    \I__7175\ : InMux
    port map (
            O => \N__33311\,
            I => \N__33202\
        );

    \I__7174\ : InMux
    port map (
            O => \N__33310\,
            I => \N__33202\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33199\
        );

    \I__7172\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33192\
        );

    \I__7171\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33192\
        );

    \I__7170\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33192\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__33297\,
            I => \N__33189\
        );

    \I__7168\ : LocalMux
    port map (
            O => \N__33294\,
            I => \N__33186\
        );

    \I__7167\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33177\
        );

    \I__7166\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33177\
        );

    \I__7165\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33177\
        );

    \I__7164\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33166\
        );

    \I__7163\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33166\
        );

    \I__7162\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33166\
        );

    \I__7161\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33166\
        );

    \I__7160\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33166\
        );

    \I__7159\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33161\
        );

    \I__7158\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33161\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__33281\,
            I => \N__33154\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__33276\,
            I => \N__33154\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__33271\,
            I => \N__33154\
        );

    \I__7154\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33149\
        );

    \I__7153\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33149\
        );

    \I__7152\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33142\
        );

    \I__7151\ : InMux
    port map (
            O => \N__33263\,
            I => \N__33142\
        );

    \I__7150\ : Span4Mux_v
    port map (
            O => \N__33260\,
            I => \N__33136\
        );

    \I__7149\ : Span4Mux_v
    port map (
            O => \N__33257\,
            I => \N__33136\
        );

    \I__7148\ : Span4Mux_h
    port map (
            O => \N__33254\,
            I => \N__33129\
        );

    \I__7147\ : LocalMux
    port map (
            O => \N__33251\,
            I => \N__33129\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__33246\,
            I => \N__33129\
        );

    \I__7145\ : Span4Mux_v
    port map (
            O => \N__33241\,
            I => \N__33124\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__33234\,
            I => \N__33124\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__33225\,
            I => \N__33121\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__33222\,
            I => \N__33112\
        );

    \I__7141\ : Span4Mux_s2_v
    port map (
            O => \N__33219\,
            I => \N__33112\
        );

    \I__7140\ : LocalMux
    port map (
            O => \N__33214\,
            I => \N__33112\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__33211\,
            I => \N__33112\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__33202\,
            I => \N__33105\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__33199\,
            I => \N__33105\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__33192\,
            I => \N__33105\
        );

    \I__7135\ : Span4Mux_v
    port map (
            O => \N__33189\,
            I => \N__33100\
        );

    \I__7134\ : Span4Mux_s2_h
    port map (
            O => \N__33186\,
            I => \N__33100\
        );

    \I__7133\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33095\
        );

    \I__7132\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33095\
        );

    \I__7131\ : LocalMux
    port map (
            O => \N__33177\,
            I => \N__33084\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__33166\,
            I => \N__33084\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__33161\,
            I => \N__33084\
        );

    \I__7128\ : Span4Mux_v
    port map (
            O => \N__33154\,
            I => \N__33084\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__33149\,
            I => \N__33084\
        );

    \I__7126\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33079\
        );

    \I__7125\ : InMux
    port map (
            O => \N__33147\,
            I => \N__33079\
        );

    \I__7124\ : LocalMux
    port map (
            O => \N__33142\,
            I => \N__33076\
        );

    \I__7123\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33073\
        );

    \I__7122\ : Span4Mux_h
    port map (
            O => \N__33136\,
            I => \N__33070\
        );

    \I__7121\ : Span4Mux_v
    port map (
            O => \N__33129\,
            I => \N__33061\
        );

    \I__7120\ : Span4Mux_h
    port map (
            O => \N__33124\,
            I => \N__33061\
        );

    \I__7119\ : Span4Mux_v
    port map (
            O => \N__33121\,
            I => \N__33061\
        );

    \I__7118\ : Span4Mux_h
    port map (
            O => \N__33112\,
            I => \N__33061\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__33105\,
            I => \N__33052\
        );

    \I__7116\ : Span4Mux_v
    port map (
            O => \N__33100\,
            I => \N__33052\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__33095\,
            I => \N__33052\
        );

    \I__7114\ : Span4Mux_v
    port map (
            O => \N__33084\,
            I => \N__33052\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__33079\,
            I => \N__33045\
        );

    \I__7112\ : Span12Mux_s1_v
    port map (
            O => \N__33076\,
            I => \N__33045\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__33073\,
            I => \N__33045\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__33070\,
            I => \clk_100Khz_signalkeep_4\
        );

    \I__7109\ : Odrv4
    port map (
            O => \N__33061\,
            I => \clk_100Khz_signalkeep_4\
        );

    \I__7108\ : Odrv4
    port map (
            O => \N__33052\,
            I => \clk_100Khz_signalkeep_4\
        );

    \I__7107\ : Odrv12
    port map (
            O => \N__33045\,
            I => \clk_100Khz_signalkeep_4\
        );

    \I__7106\ : InMux
    port map (
            O => \N__33036\,
            I => \N__33033\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__33033\,
            I => \VPP_VDDQ.curr_stateZ0Z_0\
        );

    \I__7104\ : InMux
    port map (
            O => \N__33030\,
            I => \N__33027\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__33027\,
            I => \VPP_VDDQ.count_4_10\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__33024\,
            I => \N__33020\
        );

    \I__7101\ : InMux
    port map (
            O => \N__33023\,
            I => \N__33015\
        );

    \I__7100\ : InMux
    port map (
            O => \N__33020\,
            I => \N__33015\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__33015\,
            I => \N__33008\
        );

    \I__7098\ : CascadeMux
    port map (
            O => \N__33014\,
            I => \N__33005\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__33013\,
            I => \N__33002\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__33012\,
            I => \N__32999\
        );

    \I__7095\ : InMux
    port map (
            O => \N__33011\,
            I => \N__32994\
        );

    \I__7094\ : Span4Mux_v
    port map (
            O => \N__33008\,
            I => \N__32991\
        );

    \I__7093\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32988\
        );

    \I__7092\ : InMux
    port map (
            O => \N__33002\,
            I => \N__32985\
        );

    \I__7091\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32980\
        );

    \I__7090\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32980\
        );

    \I__7089\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32977\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__32994\,
            I => \N__32967\
        );

    \I__7087\ : IoSpan4Mux
    port map (
            O => \N__32991\,
            I => \N__32967\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__32988\,
            I => \N__32958\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__32985\,
            I => \N__32958\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__32980\,
            I => \N__32958\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__32977\,
            I => \N__32958\
        );

    \I__7082\ : InMux
    port map (
            O => \N__32976\,
            I => \N__32955\
        );

    \I__7081\ : InMux
    port map (
            O => \N__32975\,
            I => \N__32952\
        );

    \I__7080\ : InMux
    port map (
            O => \N__32974\,
            I => \N__32945\
        );

    \I__7079\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32945\
        );

    \I__7078\ : InMux
    port map (
            O => \N__32972\,
            I => \N__32945\
        );

    \I__7077\ : Span4Mux_s3_h
    port map (
            O => \N__32967\,
            I => \N__32938\
        );

    \I__7076\ : Span4Mux_v
    port map (
            O => \N__32958\,
            I => \N__32938\
        );

    \I__7075\ : LocalMux
    port map (
            O => \N__32955\,
            I => \N__32938\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__32952\,
            I => \N__32932\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__32945\,
            I => \N__32932\
        );

    \I__7072\ : Span4Mux_h
    port map (
            O => \N__32938\,
            I => \N__32929\
        );

    \I__7071\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32925\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__32932\,
            I => \N__32922\
        );

    \I__7069\ : Span4Mux_h
    port map (
            O => \N__32929\,
            I => \N__32919\
        );

    \I__7068\ : InMux
    port map (
            O => \N__32928\,
            I => \N__32916\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32913\
        );

    \I__7066\ : Span4Mux_v
    port map (
            O => \N__32922\,
            I => \N__32910\
        );

    \I__7065\ : Span4Mux_v
    port map (
            O => \N__32919\,
            I => \N__32905\
        );

    \I__7064\ : LocalMux
    port map (
            O => \N__32916\,
            I => \N__32905\
        );

    \I__7063\ : Span12Mux_v
    port map (
            O => \N__32913\,
            I => \N__32900\
        );

    \I__7062\ : Sp12to4
    port map (
            O => \N__32910\,
            I => \N__32900\
        );

    \I__7061\ : Span4Mux_v
    port map (
            O => \N__32905\,
            I => \N__32897\
        );

    \I__7060\ : Odrv12
    port map (
            O => \N__32900\,
            I => gpio_fpga_soc_4
        );

    \I__7059\ : Odrv4
    port map (
            O => \N__32897\,
            I => gpio_fpga_soc_4
        );

    \I__7058\ : InMux
    port map (
            O => \N__32892\,
            I => \N__32887\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__32891\,
            I => \N__32884\
        );

    \I__7056\ : InMux
    port map (
            O => \N__32890\,
            I => \N__32881\
        );

    \I__7055\ : LocalMux
    port map (
            O => \N__32887\,
            I => \N__32878\
        );

    \I__7054\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32875\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32872\
        );

    \I__7052\ : Span4Mux_v
    port map (
            O => \N__32878\,
            I => \N__32869\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__32875\,
            I => \N__32864\
        );

    \I__7050\ : Span4Mux_v
    port map (
            O => \N__32872\,
            I => \N__32859\
        );

    \I__7049\ : Span4Mux_h
    port map (
            O => \N__32869\,
            I => \N__32859\
        );

    \I__7048\ : InMux
    port map (
            O => \N__32868\,
            I => \N__32856\
        );

    \I__7047\ : CascadeMux
    port map (
            O => \N__32867\,
            I => \N__32852\
        );

    \I__7046\ : Span4Mux_h
    port map (
            O => \N__32864\,
            I => \N__32849\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__32859\,
            I => \N__32844\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__32856\,
            I => \N__32844\
        );

    \I__7043\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32839\
        );

    \I__7042\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32839\
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__32849\,
            I => \POWERLED.N_188\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__32844\,
            I => \POWERLED.N_188\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__32839\,
            I => \POWERLED.N_188\
        );

    \I__7038\ : CascadeMux
    port map (
            O => \N__32832\,
            I => \N__32829\
        );

    \I__7037\ : InMux
    port map (
            O => \N__32829\,
            I => \N__32825\
        );

    \I__7036\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32822\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__32825\,
            I => \N__32817\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__32822\,
            I => \N__32817\
        );

    \I__7033\ : Span4Mux_v
    port map (
            O => \N__32817\,
            I => \N__32813\
        );

    \I__7032\ : InMux
    port map (
            O => \N__32816\,
            I => \N__32810\
        );

    \I__7031\ : Span4Mux_h
    port map (
            O => \N__32813\,
            I => \N__32807\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__32810\,
            I => \N__32804\
        );

    \I__7029\ : Sp12to4
    port map (
            O => \N__32807\,
            I => \N__32799\
        );

    \I__7028\ : Span12Mux_s8_v
    port map (
            O => \N__32804\,
            I => \N__32799\
        );

    \I__7027\ : Odrv12
    port map (
            O => \N__32799\,
            I => \POWERLED.N_388\
        );

    \I__7026\ : CascadeMux
    port map (
            O => \N__32796\,
            I => \N__32793\
        );

    \I__7025\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32790\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32787\
        );

    \I__7023\ : Span4Mux_v
    port map (
            O => \N__32787\,
            I => \N__32784\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__32784\,
            I => \N__32781\
        );

    \I__7021\ : Odrv4
    port map (
            O => \N__32781\,
            I => \POWERLED.un85_clk_100khz_6\
        );

    \I__7020\ : InMux
    port map (
            O => \N__32778\,
            I => \N__32773\
        );

    \I__7019\ : CascadeMux
    port map (
            O => \N__32777\,
            I => \N__32770\
        );

    \I__7018\ : CascadeMux
    port map (
            O => \N__32776\,
            I => \N__32761\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__32773\,
            I => \N__32755\
        );

    \I__7016\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32750\
        );

    \I__7015\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32750\
        );

    \I__7014\ : InMux
    port map (
            O => \N__32768\,
            I => \N__32747\
        );

    \I__7013\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32742\
        );

    \I__7012\ : InMux
    port map (
            O => \N__32766\,
            I => \N__32742\
        );

    \I__7011\ : InMux
    port map (
            O => \N__32765\,
            I => \N__32739\
        );

    \I__7010\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32728\
        );

    \I__7009\ : InMux
    port map (
            O => \N__32761\,
            I => \N__32728\
        );

    \I__7008\ : InMux
    port map (
            O => \N__32760\,
            I => \N__32728\
        );

    \I__7007\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32728\
        );

    \I__7006\ : InMux
    port map (
            O => \N__32758\,
            I => \N__32728\
        );

    \I__7005\ : Span12Mux_v
    port map (
            O => \N__32755\,
            I => \N__32725\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__32750\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7003\ : LocalMux
    port map (
            O => \N__32747\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__32742\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__32739\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__32728\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__6999\ : Odrv12
    port map (
            O => \N__32725\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__6998\ : InMux
    port map (
            O => \N__32712\,
            I => \N__32709\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__32709\,
            I => \VPP_VDDQ.count_4_6\
        );

    \I__6996\ : InMux
    port map (
            O => \N__32706\,
            I => \N__32703\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__32703\,
            I => \N__32700\
        );

    \I__6994\ : Odrv12
    port map (
            O => \N__32700\,
            I => \DSW_PWRGD.DSW_PWROK_0\
        );

    \I__6993\ : IoInMux
    port map (
            O => \N__32697\,
            I => \N__32694\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__32694\,
            I => \N__32691\
        );

    \I__6991\ : IoSpan4Mux
    port map (
            O => \N__32691\,
            I => \N__32688\
        );

    \I__6990\ : Sp12to4
    port map (
            O => \N__32688\,
            I => \N__32685\
        );

    \I__6989\ : Span12Mux_s6_h
    port map (
            O => \N__32685\,
            I => \N__32682\
        );

    \I__6988\ : Odrv12
    port map (
            O => \N__32682\,
            I => dsw_pwrok
        );

    \I__6987\ : InMux
    port map (
            O => \N__32679\,
            I => \N__32676\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__32676\,
            I => \N__32673\
        );

    \I__6985\ : Span4Mux_v
    port map (
            O => \N__32673\,
            I => \N__32670\
        );

    \I__6984\ : Odrv4
    port map (
            O => \N__32670\,
            I => v5s_ok
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__32667\,
            I => \dsw_pwrok_cascade_\
        );

    \I__6982\ : IoInMux
    port map (
            O => \N__32664\,
            I => \N__32661\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32658\
        );

    \I__6980\ : IoSpan4Mux
    port map (
            O => \N__32658\,
            I => \N__32655\
        );

    \I__6979\ : Sp12to4
    port map (
            O => \N__32655\,
            I => \N__32652\
        );

    \I__6978\ : Odrv12
    port map (
            O => \N__32652\,
            I => vccin_en
        );

    \I__6977\ : CascadeMux
    port map (
            O => \N__32649\,
            I => \N__32640\
        );

    \I__6976\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32632\
        );

    \I__6975\ : InMux
    port map (
            O => \N__32647\,
            I => \N__32623\
        );

    \I__6974\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32623\
        );

    \I__6973\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32623\
        );

    \I__6972\ : InMux
    port map (
            O => \N__32644\,
            I => \N__32618\
        );

    \I__6971\ : InMux
    port map (
            O => \N__32643\,
            I => \N__32618\
        );

    \I__6970\ : InMux
    port map (
            O => \N__32640\,
            I => \N__32615\
        );

    \I__6969\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32610\
        );

    \I__6968\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32610\
        );

    \I__6967\ : CascadeMux
    port map (
            O => \N__32637\,
            I => \N__32607\
        );

    \I__6966\ : CascadeMux
    port map (
            O => \N__32636\,
            I => \N__32604\
        );

    \I__6965\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32599\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32596\
        );

    \I__6963\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32589\
        );

    \I__6962\ : InMux
    port map (
            O => \N__32630\,
            I => \N__32589\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__32623\,
            I => \N__32580\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__32618\,
            I => \N__32580\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__32615\,
            I => \N__32580\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__32610\,
            I => \N__32580\
        );

    \I__6957\ : InMux
    port map (
            O => \N__32607\,
            I => \N__32573\
        );

    \I__6956\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32573\
        );

    \I__6955\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32573\
        );

    \I__6954\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32566\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__32599\,
            I => \N__32563\
        );

    \I__6952\ : Span4Mux_v
    port map (
            O => \N__32596\,
            I => \N__32560\
        );

    \I__6951\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32554\
        );

    \I__6950\ : InMux
    port map (
            O => \N__32594\,
            I => \N__32554\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32549\
        );

    \I__6948\ : Span4Mux_v
    port map (
            O => \N__32580\,
            I => \N__32549\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__32573\,
            I => \N__32546\
        );

    \I__6946\ : InMux
    port map (
            O => \N__32572\,
            I => \N__32539\
        );

    \I__6945\ : InMux
    port map (
            O => \N__32571\,
            I => \N__32539\
        );

    \I__6944\ : InMux
    port map (
            O => \N__32570\,
            I => \N__32539\
        );

    \I__6943\ : InMux
    port map (
            O => \N__32569\,
            I => \N__32536\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32531\
        );

    \I__6941\ : Span12Mux_s11_h
    port map (
            O => \N__32563\,
            I => \N__32531\
        );

    \I__6940\ : Span4Mux_h
    port map (
            O => \N__32560\,
            I => \N__32528\
        );

    \I__6939\ : IoInMux
    port map (
            O => \N__32559\,
            I => \N__32525\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__32554\,
            I => \N__32518\
        );

    \I__6937\ : Span4Mux_h
    port map (
            O => \N__32549\,
            I => \N__32518\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__32546\,
            I => \N__32518\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__32539\,
            I => \N__32513\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__32536\,
            I => \N__32513\
        );

    \I__6933\ : Odrv12
    port map (
            O => \N__32531\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6932\ : Odrv4
    port map (
            O => \N__32528\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__32525\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__32518\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__32513\,
            I => \VPP_VDDQ_delayed_vddq_pwrgd_en\
        );

    \I__6928\ : CascadeMux
    port map (
            O => \N__32502\,
            I => \N__32497\
        );

    \I__6927\ : InMux
    port map (
            O => \N__32501\,
            I => \N__32488\
        );

    \I__6926\ : InMux
    port map (
            O => \N__32500\,
            I => \N__32488\
        );

    \I__6925\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32477\
        );

    \I__6924\ : InMux
    port map (
            O => \N__32496\,
            I => \N__32477\
        );

    \I__6923\ : InMux
    port map (
            O => \N__32495\,
            I => \N__32477\
        );

    \I__6922\ : InMux
    port map (
            O => \N__32494\,
            I => \N__32477\
        );

    \I__6921\ : InMux
    port map (
            O => \N__32493\,
            I => \N__32477\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__32488\,
            I => \N__32474\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__32477\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__6918\ : Odrv4
    port map (
            O => \N__32474\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__6917\ : CascadeMux
    port map (
            O => \N__32469\,
            I => \N__32466\
        );

    \I__6916\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32460\
        );

    \I__6915\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32460\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__32460\,
            I => \N__32451\
        );

    \I__6913\ : InMux
    port map (
            O => \N__32459\,
            I => \N__32448\
        );

    \I__6912\ : InMux
    port map (
            O => \N__32458\,
            I => \N__32437\
        );

    \I__6911\ : InMux
    port map (
            O => \N__32457\,
            I => \N__32437\
        );

    \I__6910\ : InMux
    port map (
            O => \N__32456\,
            I => \N__32437\
        );

    \I__6909\ : InMux
    port map (
            O => \N__32455\,
            I => \N__32437\
        );

    \I__6908\ : InMux
    port map (
            O => \N__32454\,
            I => \N__32437\
        );

    \I__6907\ : Span4Mux_v
    port map (
            O => \N__32451\,
            I => \N__32434\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32429\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__32437\,
            I => \N__32429\
        );

    \I__6904\ : Span4Mux_h
    port map (
            O => \N__32434\,
            I => \N__32424\
        );

    \I__6903\ : Span4Mux_v
    port map (
            O => \N__32429\,
            I => \N__32424\
        );

    \I__6902\ : Span4Mux_v
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__6901\ : Span4Mux_h
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__6900\ : Odrv4
    port map (
            O => \N__32418\,
            I => v33dsw_ok
        );

    \I__6899\ : InMux
    port map (
            O => \N__32415\,
            I => \N__32407\
        );

    \I__6898\ : InMux
    port map (
            O => \N__32414\,
            I => \N__32407\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__32413\,
            I => \N__32404\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__32412\,
            I => \N__32399\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__32407\,
            I => \N__32395\
        );

    \I__6894\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32384\
        );

    \I__6893\ : InMux
    port map (
            O => \N__32403\,
            I => \N__32384\
        );

    \I__6892\ : InMux
    port map (
            O => \N__32402\,
            I => \N__32384\
        );

    \I__6891\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32384\
        );

    \I__6890\ : InMux
    port map (
            O => \N__32398\,
            I => \N__32384\
        );

    \I__6889\ : Odrv12
    port map (
            O => \N__32395\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__32384\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__6887\ : InMux
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__32376\,
            I => \DSW_PWRGD.curr_state_RNI3E27Z0Z_0\
        );

    \I__6885\ : InMux
    port map (
            O => \N__32373\,
            I => \N__32370\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__6883\ : Span4Mux_v
    port map (
            O => \N__32367\,
            I => \N__32364\
        );

    \I__6882\ : Span4Mux_v
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__6881\ : Odrv4
    port map (
            O => \N__32361\,
            I => v33s_ok
        );

    \I__6880\ : InMux
    port map (
            O => \N__32358\,
            I => \N__32355\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__32355\,
            I => \N__32352\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__32352\,
            I => \N__32349\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__32349\,
            I => vccst_cpu_ok
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__32346\,
            I => \N__32343\
        );

    \I__6875\ : InMux
    port map (
            O => \N__32343\,
            I => \N__32340\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__32340\,
            I => \N__32337\
        );

    \I__6873\ : Span4Mux_v
    port map (
            O => \N__32337\,
            I => \N__32328\
        );

    \I__6872\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32317\
        );

    \I__6871\ : InMux
    port map (
            O => \N__32335\,
            I => \N__32317\
        );

    \I__6870\ : InMux
    port map (
            O => \N__32334\,
            I => \N__32317\
        );

    \I__6869\ : InMux
    port map (
            O => \N__32333\,
            I => \N__32317\
        );

    \I__6868\ : InMux
    port map (
            O => \N__32332\,
            I => \N__32317\
        );

    \I__6867\ : IoInMux
    port map (
            O => \N__32331\,
            I => \N__32313\
        );

    \I__6866\ : Span4Mux_h
    port map (
            O => \N__32328\,
            I => \N__32310\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__32317\,
            I => \N__32305\
        );

    \I__6864\ : CascadeMux
    port map (
            O => \N__32316\,
            I => \N__32302\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__32313\,
            I => \N__32297\
        );

    \I__6862\ : Span4Mux_h
    port map (
            O => \N__32310\,
            I => \N__32293\
        );

    \I__6861\ : InMux
    port map (
            O => \N__32309\,
            I => \N__32288\
        );

    \I__6860\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32288\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__32305\,
            I => \N__32284\
        );

    \I__6858\ : InMux
    port map (
            O => \N__32302\,
            I => \N__32275\
        );

    \I__6857\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32275\
        );

    \I__6856\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32272\
        );

    \I__6855\ : IoSpan4Mux
    port map (
            O => \N__32297\,
            I => \N__32269\
        );

    \I__6854\ : IoInMux
    port map (
            O => \N__32296\,
            I => \N__32266\
        );

    \I__6853\ : Sp12to4
    port map (
            O => \N__32293\,
            I => \N__32261\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__32288\,
            I => \N__32261\
        );

    \I__6851\ : InMux
    port map (
            O => \N__32287\,
            I => \N__32258\
        );

    \I__6850\ : Span4Mux_v
    port map (
            O => \N__32284\,
            I => \N__32255\
        );

    \I__6849\ : InMux
    port map (
            O => \N__32283\,
            I => \N__32246\
        );

    \I__6848\ : InMux
    port map (
            O => \N__32282\,
            I => \N__32246\
        );

    \I__6847\ : InMux
    port map (
            O => \N__32281\,
            I => \N__32246\
        );

    \I__6846\ : InMux
    port map (
            O => \N__32280\,
            I => \N__32246\
        );

    \I__6845\ : LocalMux
    port map (
            O => \N__32275\,
            I => \N__32241\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__32272\,
            I => \N__32241\
        );

    \I__6843\ : Odrv4
    port map (
            O => \N__32269\,
            I => v5s_enn
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__32266\,
            I => v5s_enn
        );

    \I__6841\ : Odrv12
    port map (
            O => \N__32261\,
            I => v5s_enn
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__32258\,
            I => v5s_enn
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__32255\,
            I => v5s_enn
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__32246\,
            I => v5s_enn
        );

    \I__6837\ : Odrv12
    port map (
            O => \N__32241\,
            I => v5s_enn
        );

    \I__6836\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__32223\,
            I => \N__32217\
        );

    \I__6834\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32212\
        );

    \I__6833\ : InMux
    port map (
            O => \N__32221\,
            I => \N__32212\
        );

    \I__6832\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32208\
        );

    \I__6831\ : Span4Mux_v
    port map (
            O => \N__32217\,
            I => \N__32205\
        );

    \I__6830\ : LocalMux
    port map (
            O => \N__32212\,
            I => \N__32202\
        );

    \I__6829\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32199\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__32208\,
            I => \N__32196\
        );

    \I__6827\ : Span4Mux_h
    port map (
            O => \N__32205\,
            I => \N__32193\
        );

    \I__6826\ : Span4Mux_v
    port map (
            O => \N__32202\,
            I => \N__32188\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__32199\,
            I => \N__32188\
        );

    \I__6824\ : Span12Mux_v
    port map (
            O => \N__32196\,
            I => \N__32185\
        );

    \I__6823\ : Span4Mux_v
    port map (
            O => \N__32193\,
            I => \N__32180\
        );

    \I__6822\ : Span4Mux_v
    port map (
            O => \N__32188\,
            I => \N__32180\
        );

    \I__6821\ : Odrv12
    port map (
            O => \N__32185\,
            I => \N_392\
        );

    \I__6820\ : Odrv4
    port map (
            O => \N__32180\,
            I => \N_392\
        );

    \I__6819\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32172\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__32172\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_3\
        );

    \I__6817\ : InMux
    port map (
            O => \N__32169\,
            I => \N__32166\
        );

    \I__6816\ : LocalMux
    port map (
            O => \N__32166\,
            I => \VPP_VDDQ.count_4_14\
        );

    \I__6815\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__32160\,
            I => \VPP_VDDQ.count_4_5\
        );

    \I__6813\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32154\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__32154\,
            I => \VPP_VDDQ.count_4_15\
        );

    \I__6811\ : InMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__32148\,
            I => \VPP_VDDQ.un13_clk_100khz_9\
        );

    \I__6809\ : InMux
    port map (
            O => \N__32145\,
            I => \N__32142\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__32142\,
            I => \VPP_VDDQ.count_4_0\
        );

    \I__6807\ : CascadeMux
    port map (
            O => \N__32139\,
            I => \VPP_VDDQ.count_rst_5_cascade_\
        );

    \I__6806\ : CascadeMux
    port map (
            O => \N__32136\,
            I => \VPP_VDDQ.countZ0Z_0_cascade_\
        );

    \I__6805\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32130\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__32130\,
            I => \VPP_VDDQ.count_4_1\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__32127\,
            I => \VPP_VDDQ.countZ0Z_1_cascade_\
        );

    \I__6802\ : InMux
    port map (
            O => \N__32124\,
            I => \N__32121\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__32121\,
            I => \VPP_VDDQ.count_rst_6\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__32118\,
            I => \N__32113\
        );

    \I__6799\ : InMux
    port map (
            O => \N__32117\,
            I => \N__32108\
        );

    \I__6798\ : InMux
    port map (
            O => \N__32116\,
            I => \N__32103\
        );

    \I__6797\ : InMux
    port map (
            O => \N__32113\,
            I => \N__32103\
        );

    \I__6796\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32098\
        );

    \I__6795\ : InMux
    port map (
            O => \N__32111\,
            I => \N__32098\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__32108\,
            I => \N__32095\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32092\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__32098\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__6791\ : Odrv4
    port map (
            O => \N__32095\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__32092\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__6789\ : CascadeMux
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__6788\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32079\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__32079\,
            I => \N__32076\
        );

    \I__6786\ : Span4Mux_v
    port map (
            O => \N__32076\,
            I => \N__32070\
        );

    \I__6785\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32067\
        );

    \I__6784\ : InMux
    port map (
            O => \N__32074\,
            I => \N__32062\
        );

    \I__6783\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32062\
        );

    \I__6782\ : Odrv4
    port map (
            O => \N__32070\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__32067\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__32062\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__6779\ : InMux
    port map (
            O => \N__32055\,
            I => \N__32051\
        );

    \I__6778\ : CascadeMux
    port map (
            O => \N__32054\,
            I => \N__32048\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__32051\,
            I => \N__32043\
        );

    \I__6776\ : InMux
    port map (
            O => \N__32048\,
            I => \N__32036\
        );

    \I__6775\ : InMux
    port map (
            O => \N__32047\,
            I => \N__32036\
        );

    \I__6774\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32036\
        );

    \I__6773\ : Span4Mux_s2_h
    port map (
            O => \N__32043\,
            I => \N__32033\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__32036\,
            I => \N__32030\
        );

    \I__6771\ : Span4Mux_v
    port map (
            O => \N__32033\,
            I => \N__32027\
        );

    \I__6770\ : Span4Mux_v
    port map (
            O => \N__32030\,
            I => \N__32024\
        );

    \I__6769\ : Odrv4
    port map (
            O => \N__32027\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__6768\ : Odrv4
    port map (
            O => \N__32024\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__6767\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__6765\ : Odrv12
    port map (
            O => \N__32013\,
            I => \POWERLED.curr_state_0_0\
        );

    \I__6764\ : InMux
    port map (
            O => \N__32010\,
            I => \N__32007\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__6762\ : Span4Mux_h
    port map (
            O => \N__32004\,
            I => \N__32000\
        );

    \I__6761\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31997\
        );

    \I__6760\ : Odrv4
    port map (
            O => \N__32000\,
            I => \VPP_VDDQ.count_2_rst_9\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__31997\,
            I => \VPP_VDDQ.count_2_rst_9\
        );

    \I__6758\ : InMux
    port map (
            O => \N__31992\,
            I => \N__31989\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31986\
        );

    \I__6756\ : Span4Mux_v
    port map (
            O => \N__31986\,
            I => \N__31983\
        );

    \I__6755\ : Span4Mux_h
    port map (
            O => \N__31983\,
            I => \N__31980\
        );

    \I__6754\ : Odrv4
    port map (
            O => \N__31980\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__6753\ : CEMux
    port map (
            O => \N__31977\,
            I => \N__31972\
        );

    \I__6752\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31966\
        );

    \I__6751\ : InMux
    port map (
            O => \N__31975\,
            I => \N__31960\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__31972\,
            I => \N__31957\
        );

    \I__6749\ : CEMux
    port map (
            O => \N__31971\,
            I => \N__31954\
        );

    \I__6748\ : InMux
    port map (
            O => \N__31970\,
            I => \N__31948\
        );

    \I__6747\ : CEMux
    port map (
            O => \N__31969\,
            I => \N__31948\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__31966\,
            I => \N__31945\
        );

    \I__6745\ : CEMux
    port map (
            O => \N__31965\,
            I => \N__31942\
        );

    \I__6744\ : InMux
    port map (
            O => \N__31964\,
            I => \N__31937\
        );

    \I__6743\ : InMux
    port map (
            O => \N__31963\,
            I => \N__31937\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__31960\,
            I => \N__31929\
        );

    \I__6741\ : Span4Mux_h
    port map (
            O => \N__31957\,
            I => \N__31929\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__31954\,
            I => \N__31929\
        );

    \I__6739\ : CEMux
    port map (
            O => \N__31953\,
            I => \N__31926\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__31948\,
            I => \N__31910\
        );

    \I__6737\ : Span4Mux_h
    port map (
            O => \N__31945\,
            I => \N__31903\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__31942\,
            I => \N__31903\
        );

    \I__6735\ : LocalMux
    port map (
            O => \N__31937\,
            I => \N__31903\
        );

    \I__6734\ : CEMux
    port map (
            O => \N__31936\,
            I => \N__31900\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__31929\,
            I => \N__31895\
        );

    \I__6732\ : LocalMux
    port map (
            O => \N__31926\,
            I => \N__31895\
        );

    \I__6731\ : InMux
    port map (
            O => \N__31925\,
            I => \N__31888\
        );

    \I__6730\ : InMux
    port map (
            O => \N__31924\,
            I => \N__31888\
        );

    \I__6729\ : InMux
    port map (
            O => \N__31923\,
            I => \N__31888\
        );

    \I__6728\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31878\
        );

    \I__6727\ : InMux
    port map (
            O => \N__31921\,
            I => \N__31878\
        );

    \I__6726\ : InMux
    port map (
            O => \N__31920\,
            I => \N__31878\
        );

    \I__6725\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31867\
        );

    \I__6724\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31867\
        );

    \I__6723\ : InMux
    port map (
            O => \N__31917\,
            I => \N__31867\
        );

    \I__6722\ : InMux
    port map (
            O => \N__31916\,
            I => \N__31867\
        );

    \I__6721\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31867\
        );

    \I__6720\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31862\
        );

    \I__6719\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31862\
        );

    \I__6718\ : Span4Mux_v
    port map (
            O => \N__31910\,
            I => \N__31857\
        );

    \I__6717\ : Span4Mux_v
    port map (
            O => \N__31903\,
            I => \N__31857\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__31900\,
            I => \N__31850\
        );

    \I__6715\ : Span4Mux_s0_v
    port map (
            O => \N__31895\,
            I => \N__31850\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31850\
        );

    \I__6713\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31843\
        );

    \I__6712\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31843\
        );

    \I__6711\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31843\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__31878\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__31867\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__31862\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__6707\ : Odrv4
    port map (
            O => \N__31857\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__6706\ : Odrv4
    port map (
            O => \N__31850\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__31843\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\
        );

    \I__6704\ : InMux
    port map (
            O => \N__31830\,
            I => \N__31827\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__31827\,
            I => \N__31823\
        );

    \I__6702\ : InMux
    port map (
            O => \N__31826\,
            I => \N__31820\
        );

    \I__6701\ : Span4Mux_v
    port map (
            O => \N__31823\,
            I => \N__31817\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__31820\,
            I => \N__31814\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__31817\,
            I => \N__31811\
        );

    \I__6698\ : Span4Mux_v
    port map (
            O => \N__31814\,
            I => \N__31808\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__31811\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__6696\ : Odrv4
    port map (
            O => \N__31808\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__6695\ : InMux
    port map (
            O => \N__31803\,
            I => \N__31797\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__31802\,
            I => \N__31794\
        );

    \I__6693\ : InMux
    port map (
            O => \N__31801\,
            I => \N__31789\
        );

    \I__6692\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31789\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__31797\,
            I => \N__31786\
        );

    \I__6690\ : InMux
    port map (
            O => \N__31794\,
            I => \N__31783\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__31789\,
            I => \N__31780\
        );

    \I__6688\ : Span4Mux_s3_h
    port map (
            O => \N__31786\,
            I => \N__31777\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__31783\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__6686\ : Odrv4
    port map (
            O => \N__31780\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__6685\ : Odrv4
    port map (
            O => \N__31777\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__6684\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31766\
        );

    \I__6683\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31763\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31760\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__31763\,
            I => \N__31757\
        );

    \I__6680\ : Span4Mux_v
    port map (
            O => \N__31760\,
            I => \N__31752\
        );

    \I__6679\ : Span4Mux_s2_v
    port map (
            O => \N__31757\,
            I => \N__31752\
        );

    \I__6678\ : Odrv4
    port map (
            O => \N__31752\,
            I => \DSW_PWRGD.un2_count_1_cry_9_THRU_CO\
        );

    \I__6677\ : InMux
    port map (
            O => \N__31749\,
            I => \DSW_PWRGD.un2_count_1_cry_9\
        );

    \I__6676\ : InMux
    port map (
            O => \N__31746\,
            I => \DSW_PWRGD.un2_count_1_cry_10\
        );

    \I__6675\ : InMux
    port map (
            O => \N__31743\,
            I => \DSW_PWRGD.un2_count_1_cry_11\
        );

    \I__6674\ : InMux
    port map (
            O => \N__31740\,
            I => \DSW_PWRGD.un2_count_1_cry_12\
        );

    \I__6673\ : InMux
    port map (
            O => \N__31737\,
            I => \DSW_PWRGD.un2_count_1_cry_13\
        );

    \I__6672\ : InMux
    port map (
            O => \N__31734\,
            I => \DSW_PWRGD.un2_count_1_cry_14\
        );

    \I__6671\ : CascadeMux
    port map (
            O => \N__31731\,
            I => \VPP_VDDQ.un13_clk_100khz_10_cascade_\
        );

    \I__6670\ : CascadeMux
    port map (
            O => \N__31728\,
            I => \VPP_VDDQ.un13_clk_100khz_i_cascade_\
        );

    \I__6669\ : InMux
    port map (
            O => \N__31725\,
            I => \N__31722\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__31722\,
            I => \VPP_VDDQ.un13_clk_100khz_8\
        );

    \I__6667\ : InMux
    port map (
            O => \N__31719\,
            I => \N__31715\
        );

    \I__6666\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31712\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__31715\,
            I => \DSW_PWRGD.un2_count_1_axb_2\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__31712\,
            I => \DSW_PWRGD.un2_count_1_axb_2\
        );

    \I__6663\ : InMux
    port map (
            O => \N__31707\,
            I => \N__31701\
        );

    \I__6662\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31701\
        );

    \I__6661\ : LocalMux
    port map (
            O => \N__31701\,
            I => \DSW_PWRGD.un2_count_1_cry_1_THRU_CO\
        );

    \I__6660\ : InMux
    port map (
            O => \N__31698\,
            I => \DSW_PWRGD.un2_count_1_cry_1\
        );

    \I__6659\ : CascadeMux
    port map (
            O => \N__31695\,
            I => \N__31691\
        );

    \I__6658\ : CascadeMux
    port map (
            O => \N__31694\,
            I => \N__31688\
        );

    \I__6657\ : InMux
    port map (
            O => \N__31691\,
            I => \N__31682\
        );

    \I__6656\ : InMux
    port map (
            O => \N__31688\,
            I => \N__31682\
        );

    \I__6655\ : InMux
    port map (
            O => \N__31687\,
            I => \N__31679\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__31682\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__31679\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__6652\ : InMux
    port map (
            O => \N__31674\,
            I => \N__31668\
        );

    \I__6651\ : InMux
    port map (
            O => \N__31673\,
            I => \N__31668\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__31668\,
            I => \DSW_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__6649\ : InMux
    port map (
            O => \N__31665\,
            I => \DSW_PWRGD.un2_count_1_cry_2\
        );

    \I__6648\ : InMux
    port map (
            O => \N__31662\,
            I => \DSW_PWRGD.un2_count_1_cry_3\
        );

    \I__6647\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31655\
        );

    \I__6646\ : InMux
    port map (
            O => \N__31658\,
            I => \N__31652\
        );

    \I__6645\ : LocalMux
    port map (
            O => \N__31655\,
            I => \N__31649\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__31652\,
            I => \DSW_PWRGD.un2_count_1_axb_5\
        );

    \I__6643\ : Odrv12
    port map (
            O => \N__31649\,
            I => \DSW_PWRGD.un2_count_1_axb_5\
        );

    \I__6642\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31638\
        );

    \I__6641\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31638\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__6639\ : Odrv4
    port map (
            O => \N__31635\,
            I => \DSW_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__6638\ : InMux
    port map (
            O => \N__31632\,
            I => \DSW_PWRGD.un2_count_1_cry_4\
        );

    \I__6637\ : InMux
    port map (
            O => \N__31629\,
            I => \N__31623\
        );

    \I__6636\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31623\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__6634\ : Span12Mux_v
    port map (
            O => \N__31620\,
            I => \N__31617\
        );

    \I__6633\ : Odrv12
    port map (
            O => \N__31617\,
            I => \DSW_PWRGD.count_rst_8\
        );

    \I__6632\ : InMux
    port map (
            O => \N__31614\,
            I => \DSW_PWRGD.un2_count_1_cry_5\
        );

    \I__6631\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31607\
        );

    \I__6630\ : CascadeMux
    port map (
            O => \N__31610\,
            I => \N__31603\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__31607\,
            I => \N__31599\
        );

    \I__6628\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31596\
        );

    \I__6627\ : InMux
    port map (
            O => \N__31603\,
            I => \N__31593\
        );

    \I__6626\ : InMux
    port map (
            O => \N__31602\,
            I => \N__31590\
        );

    \I__6625\ : Span4Mux_s1_v
    port map (
            O => \N__31599\,
            I => \N__31585\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__31596\,
            I => \N__31585\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__31593\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__6622\ : LocalMux
    port map (
            O => \N__31590\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__6621\ : Odrv4
    port map (
            O => \N__31585\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__6620\ : InMux
    port map (
            O => \N__31578\,
            I => \N__31574\
        );

    \I__6619\ : InMux
    port map (
            O => \N__31577\,
            I => \N__31571\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__31574\,
            I => \N__31568\
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31565\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__31568\,
            I => \DSW_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__31565\,
            I => \DSW_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__6614\ : InMux
    port map (
            O => \N__31560\,
            I => \DSW_PWRGD.un2_count_1_cry_6\
        );

    \I__6613\ : InMux
    port map (
            O => \N__31557\,
            I => \N__31554\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__31554\,
            I => \N__31550\
        );

    \I__6611\ : InMux
    port map (
            O => \N__31553\,
            I => \N__31547\
        );

    \I__6610\ : Span4Mux_s3_h
    port map (
            O => \N__31550\,
            I => \N__31544\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__31547\,
            I => \DSW_PWRGD.un2_count_1_axb_8\
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__31544\,
            I => \DSW_PWRGD.un2_count_1_axb_8\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__31539\,
            I => \N__31535\
        );

    \I__6606\ : InMux
    port map (
            O => \N__31538\,
            I => \N__31530\
        );

    \I__6605\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31530\
        );

    \I__6604\ : LocalMux
    port map (
            O => \N__31530\,
            I => \N__31527\
        );

    \I__6603\ : Span4Mux_h
    port map (
            O => \N__31527\,
            I => \N__31524\
        );

    \I__6602\ : Odrv4
    port map (
            O => \N__31524\,
            I => \DSW_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__6601\ : InMux
    port map (
            O => \N__31521\,
            I => \bfn_11_3_0_\
        );

    \I__6600\ : InMux
    port map (
            O => \N__31518\,
            I => \DSW_PWRGD.un2_count_1_cry_8\
        );

    \I__6599\ : InMux
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__31512\,
            I => \DSW_PWRGD.count_rst_12\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__31509\,
            I => \DSW_PWRGD.count_rst_12_cascade_\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__31506\,
            I => \DSW_PWRGD.un2_count_1_axb_2_cascade_\
        );

    \I__6595\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31497\
        );

    \I__6594\ : InMux
    port map (
            O => \N__31502\,
            I => \N__31497\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__31497\,
            I => \DSW_PWRGD.count_1_2\
        );

    \I__6592\ : CascadeMux
    port map (
            O => \N__31494\,
            I => \DSW_PWRGD.count_rst_11_cascade_\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__31491\,
            I => \DSW_PWRGD.countZ0Z_3_cascade_\
        );

    \I__6590\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31485\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__31485\,
            I => \DSW_PWRGD.count_1_3\
        );

    \I__6588\ : InMux
    port map (
            O => \N__31482\,
            I => \N__31479\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__31479\,
            I => \N__31476\
        );

    \I__6586\ : Span4Mux_h
    port map (
            O => \N__31476\,
            I => \N__31473\
        );

    \I__6585\ : Odrv4
    port map (
            O => \N__31473\,
            I => \DSW_PWRGD.count_1_7\
        );

    \I__6584\ : InMux
    port map (
            O => \N__31470\,
            I => \DSW_PWRGD.un2_count_1_cry_0\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__31467\,
            I => \N__31462\
        );

    \I__6582\ : InMux
    port map (
            O => \N__31466\,
            I => \N__31457\
        );

    \I__6581\ : InMux
    port map (
            O => \N__31465\,
            I => \N__31454\
        );

    \I__6580\ : InMux
    port map (
            O => \N__31462\,
            I => \N__31447\
        );

    \I__6579\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31447\
        );

    \I__6578\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31447\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__31457\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__31454\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__31447\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__31440\,
            I => \N__31436\
        );

    \I__6573\ : CascadeMux
    port map (
            O => \N__31439\,
            I => \N__31432\
        );

    \I__6572\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31425\
        );

    \I__6571\ : InMux
    port map (
            O => \N__31435\,
            I => \N__31425\
        );

    \I__6570\ : InMux
    port map (
            O => \N__31432\,
            I => \N__31425\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__31425\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__31422\,
            I => \N__31412\
        );

    \I__6567\ : CascadeMux
    port map (
            O => \N__31421\,
            I => \N__31409\
        );

    \I__6566\ : InMux
    port map (
            O => \N__31420\,
            I => \N__31406\
        );

    \I__6565\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31401\
        );

    \I__6564\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31401\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__31417\,
            I => \N__31397\
        );

    \I__6562\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31388\
        );

    \I__6561\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31388\
        );

    \I__6560\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31388\
        );

    \I__6559\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31388\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__31406\,
            I => \N__31385\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31382\
        );

    \I__6556\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31377\
        );

    \I__6555\ : InMux
    port map (
            O => \N__31397\,
            I => \N__31377\
        );

    \I__6554\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31372\
        );

    \I__6553\ : Span4Mux_s3_v
    port map (
            O => \N__31385\,
            I => \N__31365\
        );

    \I__6552\ : Span4Mux_v
    port map (
            O => \N__31382\,
            I => \N__31365\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__31377\,
            I => \N__31365\
        );

    \I__6550\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31362\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__31375\,
            I => \N__31356\
        );

    \I__6548\ : Span4Mux_s3_v
    port map (
            O => \N__31372\,
            I => \N__31348\
        );

    \I__6547\ : Span4Mux_h
    port map (
            O => \N__31365\,
            I => \N__31348\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__31362\,
            I => \N__31348\
        );

    \I__6545\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31339\
        );

    \I__6544\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31339\
        );

    \I__6543\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31339\
        );

    \I__6542\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31339\
        );

    \I__6541\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31336\
        );

    \I__6540\ : Span4Mux_h
    port map (
            O => \N__31348\,
            I => \N__31333\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__31339\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__31336\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__31333\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6536\ : CascadeMux
    port map (
            O => \N__31326\,
            I => \N__31323\
        );

    \I__6535\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31320\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31317\
        );

    \I__6533\ : Odrv4
    port map (
            O => \N__31317\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__31314\,
            I => \N__31310\
        );

    \I__6531\ : InMux
    port map (
            O => \N__31313\,
            I => \N__31302\
        );

    \I__6530\ : InMux
    port map (
            O => \N__31310\,
            I => \N__31302\
        );

    \I__6529\ : InMux
    port map (
            O => \N__31309\,
            I => \N__31302\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__31302\,
            I => \G_3119\
        );

    \I__6527\ : InMux
    port map (
            O => \N__31299\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__31296\,
            I => \N__31293\
        );

    \I__6525\ : InMux
    port map (
            O => \N__31293\,
            I => \N__31290\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__31290\,
            I => \N__31287\
        );

    \I__6523\ : Span4Mux_v
    port map (
            O => \N__31287\,
            I => \N__31284\
        );

    \I__6522\ : Span4Mux_v
    port map (
            O => \N__31284\,
            I => \N__31281\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__31281\,
            I => \POWERLED.un85_clk_100khz_0\
        );

    \I__6520\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31275\
        );

    \I__6519\ : LocalMux
    port map (
            O => \N__31275\,
            I => \N__31272\
        );

    \I__6518\ : Span4Mux_v
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__31269\,
            I => \DSW_PWRGD.un12_clk_100khz_4\
        );

    \I__6516\ : InMux
    port map (
            O => \N__31266\,
            I => \N__31263\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__31263\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__6514\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31256\
        );

    \I__6513\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31253\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__31256\,
            I => \N__31250\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__31253\,
            I => \N__31245\
        );

    \I__6510\ : Span4Mux_s2_v
    port map (
            O => \N__31250\,
            I => \N__31245\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__31245\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__6508\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31239\
        );

    \I__6507\ : LocalMux
    port map (
            O => \N__31239\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__6506\ : CascadeMux
    port map (
            O => \N__31236\,
            I => \N__31233\
        );

    \I__6505\ : InMux
    port map (
            O => \N__31233\,
            I => \N__31230\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__31230\,
            I => \N__31227\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__31227\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__6502\ : InMux
    port map (
            O => \N__31224\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__31221\,
            I => \N__31218\
        );

    \I__6500\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31215\
        );

    \I__6499\ : LocalMux
    port map (
            O => \N__31215\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__6498\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31209\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__31209\,
            I => \N__31206\
        );

    \I__6496\ : Odrv4
    port map (
            O => \N__31206\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__6495\ : InMux
    port map (
            O => \N__31203\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__6494\ : CascadeMux
    port map (
            O => \N__31200\,
            I => \N__31197\
        );

    \I__6493\ : InMux
    port map (
            O => \N__31197\,
            I => \N__31194\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__31194\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__6490\ : InMux
    port map (
            O => \N__31188\,
            I => \N__31185\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__31185\,
            I => \N__31182\
        );

    \I__6488\ : Odrv4
    port map (
            O => \N__31182\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__6487\ : InMux
    port map (
            O => \N__31179\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__6486\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31173\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__31173\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__6484\ : InMux
    port map (
            O => \N__31170\,
            I => \N__31167\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31164\
        );

    \I__6482\ : Odrv4
    port map (
            O => \N__31164\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__6481\ : InMux
    port map (
            O => \N__31161\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__6480\ : InMux
    port map (
            O => \N__31158\,
            I => \N__31155\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__31155\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__31152\,
            I => \N__31149\
        );

    \I__6477\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31146\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__31146\,
            I => \N__31143\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__31143\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__6474\ : InMux
    port map (
            O => \N__31140\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__6473\ : CascadeMux
    port map (
            O => \N__31137\,
            I => \N__31134\
        );

    \I__6472\ : InMux
    port map (
            O => \N__31134\,
            I => \N__31131\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__31131\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__6470\ : InMux
    port map (
            O => \N__31128\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__6469\ : CascadeMux
    port map (
            O => \N__31125\,
            I => \N__31120\
        );

    \I__6468\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31117\
        );

    \I__6467\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31112\
        );

    \I__6466\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31112\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__31117\,
            I => \N__31107\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__31112\,
            I => \N__31104\
        );

    \I__6463\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31101\
        );

    \I__6462\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31098\
        );

    \I__6461\ : Odrv12
    port map (
            O => \N__31107\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__6460\ : Odrv4
    port map (
            O => \N__31104\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__6459\ : LocalMux
    port map (
            O => \N__31101\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__31098\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__6457\ : CascadeMux
    port map (
            O => \N__31089\,
            I => \N__31086\
        );

    \I__6456\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31083\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__31083\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__6454\ : InMux
    port map (
            O => \N__31080\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__6453\ : InMux
    port map (
            O => \N__31077\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__6452\ : InMux
    port map (
            O => \N__31074\,
            I => \N__31070\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__31073\,
            I => \N__31066\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__31070\,
            I => \N__31061\
        );

    \I__6449\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31058\
        );

    \I__6448\ : InMux
    port map (
            O => \N__31066\,
            I => \N__31051\
        );

    \I__6447\ : InMux
    port map (
            O => \N__31065\,
            I => \N__31051\
        );

    \I__6446\ : InMux
    port map (
            O => \N__31064\,
            I => \N__31051\
        );

    \I__6445\ : Odrv4
    port map (
            O => \N__31061\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__6444\ : LocalMux
    port map (
            O => \N__31058\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__31051\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__6442\ : InMux
    port map (
            O => \N__31044\,
            I => \N__31038\
        );

    \I__6441\ : InMux
    port map (
            O => \N__31043\,
            I => \N__31038\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__31038\,
            I => \N__31035\
        );

    \I__6439\ : Span4Mux_h
    port map (
            O => \N__31035\,
            I => \N__31032\
        );

    \I__6438\ : Odrv4
    port map (
            O => \N__31032\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__6437\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31026\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__31026\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__31023\,
            I => \N__31019\
        );

    \I__6434\ : CascadeMux
    port map (
            O => \N__31022\,
            I => \N__31015\
        );

    \I__6433\ : InMux
    port map (
            O => \N__31019\,
            I => \N__31008\
        );

    \I__6432\ : InMux
    port map (
            O => \N__31018\,
            I => \N__31008\
        );

    \I__6431\ : InMux
    port map (
            O => \N__31015\,
            I => \N__31008\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__31008\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__6429\ : CascadeMux
    port map (
            O => \N__31005\,
            I => \N__31001\
        );

    \I__6428\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30998\
        );

    \I__6427\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30995\
        );

    \I__6426\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30992\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__30995\,
            I => \N__30989\
        );

    \I__6424\ : Odrv4
    port map (
            O => \N__30992\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__6423\ : Odrv4
    port map (
            O => \N__30989\,
            I => \POWERLED.mult1_un47_sum\
        );

    \I__6422\ : CascadeMux
    port map (
            O => \N__30984\,
            I => \N__30981\
        );

    \I__6421\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30978\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__30978\,
            I => \POWERLED.mult1_un47_sum_i\
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__30975\,
            I => \N__30972\
        );

    \I__6418\ : InMux
    port map (
            O => \N__30972\,
            I => \N__30969\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__30969\,
            I => \N__30965\
        );

    \I__6416\ : IoInMux
    port map (
            O => \N__30968\,
            I => \N__30962\
        );

    \I__6415\ : Span4Mux_s2_v
    port map (
            O => \N__30965\,
            I => \N__30959\
        );

    \I__6414\ : LocalMux
    port map (
            O => \N__30962\,
            I => \N__30956\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__30959\,
            I => \N__30953\
        );

    \I__6412\ : Span4Mux_s3_h
    port map (
            O => \N__30956\,
            I => \N__30949\
        );

    \I__6411\ : Span4Mux_v
    port map (
            O => \N__30953\,
            I => \N__30946\
        );

    \I__6410\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30943\
        );

    \I__6409\ : Sp12to4
    port map (
            O => \N__30949\,
            I => \N__30940\
        );

    \I__6408\ : Span4Mux_h
    port map (
            O => \N__30946\,
            I => \N__30935\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__30943\,
            I => \N__30935\
        );

    \I__6406\ : Span12Mux_v
    port map (
            O => \N__30940\,
            I => \N__30932\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__30935\,
            I => \N__30929\
        );

    \I__6404\ : Odrv12
    port map (
            O => \N__30932\,
            I => v33a_ok
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__30929\,
            I => v33a_ok
        );

    \I__6402\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__30921\,
            I => \N__30918\
        );

    \I__6400\ : Span4Mux_v
    port map (
            O => \N__30918\,
            I => \N__30915\
        );

    \I__6399\ : Span4Mux_v
    port map (
            O => \N__30915\,
            I => \N__30912\
        );

    \I__6398\ : Span4Mux_h
    port map (
            O => \N__30912\,
            I => \N__30908\
        );

    \I__6397\ : InMux
    port map (
            O => \N__30911\,
            I => \N__30905\
        );

    \I__6396\ : Span4Mux_v
    port map (
            O => \N__30908\,
            I => \N__30900\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__30905\,
            I => \N__30900\
        );

    \I__6394\ : Odrv4
    port map (
            O => \N__30900\,
            I => slp_susn
        );

    \I__6393\ : IoInMux
    port map (
            O => \N__30897\,
            I => \N__30894\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__30894\,
            I => \N__30891\
        );

    \I__6391\ : Span12Mux_s2_h
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__6390\ : Odrv12
    port map (
            O => \N__30888\,
            I => v1p8a_en
        );

    \I__6389\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30881\
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__30884\,
            I => \N__30878\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__30881\,
            I => \N__30875\
        );

    \I__6386\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30872\
        );

    \I__6385\ : Odrv4
    port map (
            O => \N__30875\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__30872\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__6383\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30864\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__30864\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__6381\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30858\
        );

    \I__6380\ : LocalMux
    port map (
            O => \N__30858\,
            I => \N__30855\
        );

    \I__6379\ : Odrv12
    port map (
            O => \N__30855\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__6378\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30849\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__30849\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__6376\ : InMux
    port map (
            O => \N__30846\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__6375\ : CascadeMux
    port map (
            O => \N__30843\,
            I => \N__30840\
        );

    \I__6374\ : InMux
    port map (
            O => \N__30840\,
            I => \N__30837\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__30837\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__6372\ : InMux
    port map (
            O => \N__30834\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__6371\ : InMux
    port map (
            O => \N__30831\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__30828\,
            I => \N__30823\
        );

    \I__6369\ : InMux
    port map (
            O => \N__30827\,
            I => \N__30818\
        );

    \I__6368\ : InMux
    port map (
            O => \N__30826\,
            I => \N__30815\
        );

    \I__6367\ : InMux
    port map (
            O => \N__30823\,
            I => \N__30808\
        );

    \I__6366\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30808\
        );

    \I__6365\ : InMux
    port map (
            O => \N__30821\,
            I => \N__30808\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__30818\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__30815\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__30808\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__6361\ : CascadeMux
    port map (
            O => \N__30801\,
            I => \N__30797\
        );

    \I__6360\ : CascadeMux
    port map (
            O => \N__30800\,
            I => \N__30793\
        );

    \I__6359\ : InMux
    port map (
            O => \N__30797\,
            I => \N__30786\
        );

    \I__6358\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30786\
        );

    \I__6357\ : InMux
    port map (
            O => \N__30793\,
            I => \N__30786\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__30786\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__30783\,
            I => \N__30780\
        );

    \I__6354\ : InMux
    port map (
            O => \N__30780\,
            I => \N__30777\
        );

    \I__6353\ : LocalMux
    port map (
            O => \N__30777\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__6352\ : InMux
    port map (
            O => \N__30774\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__6351\ : CascadeMux
    port map (
            O => \N__30771\,
            I => \N__30768\
        );

    \I__6350\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30765\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__30765\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__6348\ : InMux
    port map (
            O => \N__30762\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__6347\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__30756\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__6345\ : InMux
    port map (
            O => \N__30753\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__6344\ : InMux
    port map (
            O => \N__30750\,
            I => \N__30747\
        );

    \I__6343\ : LocalMux
    port map (
            O => \N__30747\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__6342\ : InMux
    port map (
            O => \N__30744\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__6341\ : InMux
    port map (
            O => \N__30741\,
            I => \bfn_9_11_0_\
        );

    \I__6340\ : CascadeMux
    port map (
            O => \N__30738\,
            I => \N__30734\
        );

    \I__6339\ : CascadeMux
    port map (
            O => \N__30737\,
            I => \N__30731\
        );

    \I__6338\ : InMux
    port map (
            O => \N__30734\,
            I => \N__30725\
        );

    \I__6337\ : InMux
    port map (
            O => \N__30731\,
            I => \N__30720\
        );

    \I__6336\ : InMux
    port map (
            O => \N__30730\,
            I => \N__30720\
        );

    \I__6335\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30717\
        );

    \I__6334\ : InMux
    port map (
            O => \N__30728\,
            I => \N__30714\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__30725\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__30720\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__30717\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__30714\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__6329\ : CascadeMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__6328\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__6327\ : LocalMux
    port map (
            O => \N__30699\,
            I => \POWERLED.mult1_un89_sum_i_8\
        );

    \I__6326\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__30693\,
            I => \POWERLED.mult1_un68_sum_i_8\
        );

    \I__6324\ : InMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__6323\ : LocalMux
    port map (
            O => \N__30687\,
            I => \POWERLED.mult1_un75_sum_i_8\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__30684\,
            I => \N__30681\
        );

    \I__6321\ : InMux
    port map (
            O => \N__30681\,
            I => \N__30678\
        );

    \I__6320\ : LocalMux
    port map (
            O => \N__30678\,
            I => \POWERLED.mult1_un82_sum_i_8\
        );

    \I__6319\ : CascadeMux
    port map (
            O => \N__30675\,
            I => \N__30672\
        );

    \I__6318\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30669\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__30669\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__6316\ : InMux
    port map (
            O => \N__30666\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__6315\ : CascadeMux
    port map (
            O => \N__30663\,
            I => \N__30660\
        );

    \I__6314\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30657\
        );

    \I__6313\ : LocalMux
    port map (
            O => \N__30657\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__6312\ : InMux
    port map (
            O => \N__30654\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__6311\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30648\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__30648\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__6309\ : InMux
    port map (
            O => \N__30645\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__6308\ : InMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__6306\ : Span4Mux_v
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__30633\,
            I => \POWERLED.mult1_un103_sum_i_8\
        );

    \I__6304\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__6302\ : Span12Mux_s11_v
    port map (
            O => \N__30624\,
            I => \N__30619\
        );

    \I__6301\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30616\
        );

    \I__6300\ : InMux
    port map (
            O => \N__30622\,
            I => \N__30613\
        );

    \I__6299\ : Odrv12
    port map (
            O => \N__30619\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__30616\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__30613\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__6296\ : CascadeMux
    port map (
            O => \N__30606\,
            I => \N__30603\
        );

    \I__6295\ : InMux
    port map (
            O => \N__30603\,
            I => \N__30600\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__30600\,
            I => \POWERLED.N_6486_i\
        );

    \I__6293\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30592\
        );

    \I__6292\ : CascadeMux
    port map (
            O => \N__30596\,
            I => \N__30589\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__30595\,
            I => \N__30586\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__30592\,
            I => \N__30583\
        );

    \I__6289\ : InMux
    port map (
            O => \N__30589\,
            I => \N__30578\
        );

    \I__6288\ : InMux
    port map (
            O => \N__30586\,
            I => \N__30578\
        );

    \I__6287\ : Odrv12
    port map (
            O => \N__30583\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__30578\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__6285\ : InMux
    port map (
            O => \N__30573\,
            I => \N__30570\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__30570\,
            I => \POWERLED.N_6487_i\
        );

    \I__6283\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30564\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__30564\,
            I => \N__30560\
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__30563\,
            I => \N__30557\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__30560\,
            I => \N__30553\
        );

    \I__6279\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30548\
        );

    \I__6278\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30548\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__30553\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__30548\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__6275\ : InMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__30540\,
            I => \POWERLED.N_6488_i\
        );

    \I__6273\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__30534\,
            I => \N__30531\
        );

    \I__6271\ : Span4Mux_v
    port map (
            O => \N__30531\,
            I => \N__30526\
        );

    \I__6270\ : InMux
    port map (
            O => \N__30530\,
            I => \N__30521\
        );

    \I__6269\ : InMux
    port map (
            O => \N__30529\,
            I => \N__30521\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__30526\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__30521\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__6266\ : InMux
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__30513\,
            I => \POWERLED.N_6489_i\
        );

    \I__6264\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30507\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__30507\,
            I => \N__30504\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__30504\,
            I => \N__30499\
        );

    \I__6261\ : InMux
    port map (
            O => \N__30503\,
            I => \N__30494\
        );

    \I__6260\ : InMux
    port map (
            O => \N__30502\,
            I => \N__30494\
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__30499\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__30494\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__6256\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__30483\,
            I => \POWERLED.N_6490_i\
        );

    \I__6254\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30476\
        );

    \I__6253\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30472\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__30476\,
            I => \N__30469\
        );

    \I__6251\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30466\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__30472\,
            I => \N__30463\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__30469\,
            I => \N__30458\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__30466\,
            I => \N__30458\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__30463\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__30458\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__6245\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__6244\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__30447\,
            I => \POWERLED.N_6491_i\
        );

    \I__6242\ : InMux
    port map (
            O => \N__30444\,
            I => \N__30441\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__6240\ : Span4Mux_v
    port map (
            O => \N__30438\,
            I => \N__30434\
        );

    \I__6239\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30431\
        );

    \I__6238\ : Span4Mux_v
    port map (
            O => \N__30434\,
            I => \N__30427\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__30431\,
            I => \N__30424\
        );

    \I__6236\ : InMux
    port map (
            O => \N__30430\,
            I => \N__30421\
        );

    \I__6235\ : Odrv4
    port map (
            O => \N__30427\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__6234\ : Odrv4
    port map (
            O => \N__30424\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__6233\ : LocalMux
    port map (
            O => \N__30421\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__6232\ : CascadeMux
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__6231\ : InMux
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__30408\,
            I => \POWERLED.N_6492_i\
        );

    \I__6229\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30401\
        );

    \I__6228\ : CascadeMux
    port map (
            O => \N__30404\,
            I => \N__30397\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__30401\,
            I => \N__30394\
        );

    \I__6226\ : InMux
    port map (
            O => \N__30400\,
            I => \N__30391\
        );

    \I__6225\ : InMux
    port map (
            O => \N__30397\,
            I => \N__30388\
        );

    \I__6224\ : Odrv12
    port map (
            O => \N__30394\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__30391\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__30388\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__6220\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30375\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__30375\,
            I => \POWERLED.N_6478_i\
        );

    \I__6218\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30367\
        );

    \I__6217\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30364\
        );

    \I__6216\ : InMux
    port map (
            O => \N__30370\,
            I => \N__30361\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__30367\,
            I => \N__30358\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__30364\,
            I => \N__30353\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__30361\,
            I => \N__30353\
        );

    \I__6212\ : Odrv4
    port map (
            O => \N__30358\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__30353\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__6210\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__30345\,
            I => \POWERLED.N_6479_i\
        );

    \I__6208\ : InMux
    port map (
            O => \N__30342\,
            I => \N__30337\
        );

    \I__6207\ : InMux
    port map (
            O => \N__30341\,
            I => \N__30334\
        );

    \I__6206\ : CascadeMux
    port map (
            O => \N__30340\,
            I => \N__30331\
        );

    \I__6205\ : LocalMux
    port map (
            O => \N__30337\,
            I => \N__30328\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__30334\,
            I => \N__30325\
        );

    \I__6203\ : InMux
    port map (
            O => \N__30331\,
            I => \N__30322\
        );

    \I__6202\ : Span4Mux_v
    port map (
            O => \N__30328\,
            I => \N__30319\
        );

    \I__6201\ : Span4Mux_v
    port map (
            O => \N__30325\,
            I => \N__30316\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__30322\,
            I => \N__30313\
        );

    \I__6199\ : Odrv4
    port map (
            O => \N__30319\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__30316\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__30313\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__30306\,
            I => \N__30303\
        );

    \I__6195\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30300\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__30300\,
            I => \POWERLED.N_6480_i\
        );

    \I__6193\ : InMux
    port map (
            O => \N__30297\,
            I => \N__30292\
        );

    \I__6192\ : InMux
    port map (
            O => \N__30296\,
            I => \N__30289\
        );

    \I__6191\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30286\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30283\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__30289\,
            I => \N__30280\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__30286\,
            I => \N__30275\
        );

    \I__6187\ : Span4Mux_h
    port map (
            O => \N__30283\,
            I => \N__30275\
        );

    \I__6186\ : Odrv4
    port map (
            O => \N__30280\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__6185\ : Odrv4
    port map (
            O => \N__30275\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__6184\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__30267\,
            I => \POWERLED.N_6481_i\
        );

    \I__6182\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30257\
        );

    \I__6180\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30253\
        );

    \I__6179\ : Span4Mux_v
    port map (
            O => \N__30257\,
            I => \N__30250\
        );

    \I__6178\ : InMux
    port map (
            O => \N__30256\,
            I => \N__30247\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__30253\,
            I => \N__30244\
        );

    \I__6176\ : Odrv4
    port map (
            O => \N__30250\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__30247\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__6174\ : Odrv4
    port map (
            O => \N__30244\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__6173\ : InMux
    port map (
            O => \N__30237\,
            I => \N__30234\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__30234\,
            I => \POWERLED.N_6482_i\
        );

    \I__6171\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30228\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__30228\,
            I => \N__30224\
        );

    \I__6169\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30220\
        );

    \I__6168\ : Span4Mux_v
    port map (
            O => \N__30224\,
            I => \N__30217\
        );

    \I__6167\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30214\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__30220\,
            I => \N__30211\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__30217\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__30214\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__6163\ : Odrv4
    port map (
            O => \N__30211\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__6162\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30201\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__30201\,
            I => \POWERLED.N_6483_i\
        );

    \I__6160\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30195\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__30195\,
            I => \N__30192\
        );

    \I__6158\ : Span4Mux_v
    port map (
            O => \N__30192\,
            I => \N__30187\
        );

    \I__6157\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30184\
        );

    \I__6156\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30181\
        );

    \I__6155\ : Odrv4
    port map (
            O => \N__30187\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__30184\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__30181\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__6152\ : CascadeMux
    port map (
            O => \N__30174\,
            I => \N__30171\
        );

    \I__6151\ : InMux
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__30168\,
            I => \N__30165\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__30165\,
            I => \N__30162\
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__30162\,
            I => \POWERLED.un85_clk_100khz_7\
        );

    \I__6147\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__6146\ : LocalMux
    port map (
            O => \N__30156\,
            I => \POWERLED.N_6484_i\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__30153\,
            I => \N__30150\
        );

    \I__6144\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__30147\,
            I => \N__30144\
        );

    \I__6142\ : Span4Mux_v
    port map (
            O => \N__30144\,
            I => \N__30141\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__30141\,
            I => \POWERLED.un85_clk_100khz_8\
        );

    \I__6140\ : InMux
    port map (
            O => \N__30138\,
            I => \N__30135\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__30135\,
            I => \N__30132\
        );

    \I__6138\ : Span4Mux_v
    port map (
            O => \N__30132\,
            I => \N__30129\
        );

    \I__6137\ : Span4Mux_v
    port map (
            O => \N__30129\,
            I => \N__30124\
        );

    \I__6136\ : InMux
    port map (
            O => \N__30128\,
            I => \N__30121\
        );

    \I__6135\ : InMux
    port map (
            O => \N__30127\,
            I => \N__30118\
        );

    \I__6134\ : Odrv4
    port map (
            O => \N__30124\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__30121\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__30118\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__6131\ : InMux
    port map (
            O => \N__30111\,
            I => \N__30108\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__30108\,
            I => \POWERLED.N_6485_i\
        );

    \I__6129\ : InMux
    port map (
            O => \N__30105\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__6128\ : InMux
    port map (
            O => \N__30102\,
            I => \N__30099\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__30099\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__6126\ : InMux
    port map (
            O => \N__30096\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__30093\,
            I => \N__30090\
        );

    \I__6124\ : InMux
    port map (
            O => \N__30090\,
            I => \N__30087\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__30087\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__6122\ : InMux
    port map (
            O => \N__30084\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__6121\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30078\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__30078\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__6119\ : InMux
    port map (
            O => \N__30075\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__6118\ : CascadeMux
    port map (
            O => \N__30072\,
            I => \N__30069\
        );

    \I__6117\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30066\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__30066\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__6115\ : InMux
    port map (
            O => \N__30063\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__6114\ : InMux
    port map (
            O => \N__30060\,
            I => \N__30057\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__30057\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__6112\ : InMux
    port map (
            O => \N__30054\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__30051\,
            I => \N__30048\
        );

    \I__6110\ : InMux
    port map (
            O => \N__30048\,
            I => \N__30037\
        );

    \I__6109\ : InMux
    port map (
            O => \N__30047\,
            I => \N__30037\
        );

    \I__6108\ : InMux
    port map (
            O => \N__30046\,
            I => \N__30037\
        );

    \I__6107\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30034\
        );

    \I__6106\ : InMux
    port map (
            O => \N__30044\,
            I => \N__30031\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__30037\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__30034\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__30031\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__30024\,
            I => \N__30020\
        );

    \I__6101\ : InMux
    port map (
            O => \N__30023\,
            I => \N__30012\
        );

    \I__6100\ : InMux
    port map (
            O => \N__30020\,
            I => \N__30012\
        );

    \I__6099\ : InMux
    port map (
            O => \N__30019\,
            I => \N__30012\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__30012\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__6097\ : InMux
    port map (
            O => \N__30009\,
            I => \N__30005\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__30008\,
            I => \N__29999\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__30005\,
            I => \N__29995\
        );

    \I__6094\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29992\
        );

    \I__6093\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29989\
        );

    \I__6092\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29982\
        );

    \I__6091\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29982\
        );

    \I__6090\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29982\
        );

    \I__6089\ : Odrv12
    port map (
            O => \N__29995\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__29992\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__29989\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__29982\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__6085\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29970\
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__29970\,
            I => \POWERLED.un1_count_cry_0_i\
        );

    \I__6083\ : CascadeMux
    port map (
            O => \N__29967\,
            I => \N__29964\
        );

    \I__6082\ : InMux
    port map (
            O => \N__29964\,
            I => \N__29958\
        );

    \I__6081\ : InMux
    port map (
            O => \N__29963\,
            I => \N__29958\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__29958\,
            I => \POWERLED.count_1_2\
        );

    \I__6079\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29952\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__29952\,
            I => \POWERLED.count_0_2\
        );

    \I__6077\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29946\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__29946\,
            I => \DSW_PWRGD.count_1_6\
        );

    \I__6075\ : InMux
    port map (
            O => \N__29943\,
            I => \N__29940\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29937\
        );

    \I__6073\ : Span12Mux_s8_h
    port map (
            O => \N__29937\,
            I => \N__29934\
        );

    \I__6072\ : Odrv12
    port map (
            O => \N__29934\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__6071\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29928\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__29928\,
            I => \N__29924\
        );

    \I__6069\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29921\
        );

    \I__6068\ : Span4Mux_v
    port map (
            O => \N__29924\,
            I => \N__29918\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__29921\,
            I => \N__29915\
        );

    \I__6066\ : Span4Mux_h
    port map (
            O => \N__29918\,
            I => \N__29912\
        );

    \I__6065\ : Span4Mux_h
    port map (
            O => \N__29915\,
            I => \N__29909\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__29912\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__6063\ : Odrv4
    port map (
            O => \N__29909\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__6062\ : CEMux
    port map (
            O => \N__29904\,
            I => \N__29901\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__29901\,
            I => \N__29898\
        );

    \I__6060\ : Span4Mux_s2_v
    port map (
            O => \N__29898\,
            I => \N__29891\
        );

    \I__6059\ : CEMux
    port map (
            O => \N__29897\,
            I => \N__29888\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__29896\,
            I => \N__29883\
        );

    \I__6057\ : InMux
    port map (
            O => \N__29895\,
            I => \N__29880\
        );

    \I__6056\ : CEMux
    port map (
            O => \N__29894\,
            I => \N__29862\
        );

    \I__6055\ : Span4Mux_s2_h
    port map (
            O => \N__29891\,
            I => \N__29857\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__29888\,
            I => \N__29857\
        );

    \I__6053\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29850\
        );

    \I__6052\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29850\
        );

    \I__6051\ : InMux
    port map (
            O => \N__29883\,
            I => \N__29850\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29847\
        );

    \I__6049\ : CEMux
    port map (
            O => \N__29879\,
            I => \N__29844\
        );

    \I__6048\ : CEMux
    port map (
            O => \N__29878\,
            I => \N__29841\
        );

    \I__6047\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29834\
        );

    \I__6046\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29834\
        );

    \I__6045\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29834\
        );

    \I__6044\ : CEMux
    port map (
            O => \N__29874\,
            I => \N__29827\
        );

    \I__6043\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29814\
        );

    \I__6042\ : CEMux
    port map (
            O => \N__29872\,
            I => \N__29814\
        );

    \I__6041\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29814\
        );

    \I__6040\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29814\
        );

    \I__6039\ : InMux
    port map (
            O => \N__29869\,
            I => \N__29814\
        );

    \I__6038\ : InMux
    port map (
            O => \N__29868\,
            I => \N__29814\
        );

    \I__6037\ : InMux
    port map (
            O => \N__29867\,
            I => \N__29807\
        );

    \I__6036\ : InMux
    port map (
            O => \N__29866\,
            I => \N__29807\
        );

    \I__6035\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29807\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__29862\,
            I => \N__29804\
        );

    \I__6033\ : Span4Mux_h
    port map (
            O => \N__29857\,
            I => \N__29799\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__29850\,
            I => \N__29799\
        );

    \I__6031\ : Span4Mux_h
    port map (
            O => \N__29847\,
            I => \N__29796\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__29844\,
            I => \N__29789\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__29841\,
            I => \N__29789\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__29834\,
            I => \N__29789\
        );

    \I__6027\ : InMux
    port map (
            O => \N__29833\,
            I => \N__29780\
        );

    \I__6026\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29780\
        );

    \I__6025\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29780\
        );

    \I__6024\ : InMux
    port map (
            O => \N__29830\,
            I => \N__29780\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__29827\,
            I => \N__29774\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__29814\,
            I => \N__29769\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__29807\,
            I => \N__29769\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__29804\,
            I => \N__29766\
        );

    \I__6019\ : Span4Mux_s2_v
    port map (
            O => \N__29799\,
            I => \N__29761\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__29796\,
            I => \N__29761\
        );

    \I__6017\ : Span4Mux_s2_v
    port map (
            O => \N__29789\,
            I => \N__29756\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__29780\,
            I => \N__29756\
        );

    \I__6015\ : InMux
    port map (
            O => \N__29779\,
            I => \N__29749\
        );

    \I__6014\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29749\
        );

    \I__6013\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29749\
        );

    \I__6012\ : Span4Mux_h
    port map (
            O => \N__29774\,
            I => \N__29744\
        );

    \I__6011\ : Span4Mux_s3_h
    port map (
            O => \N__29769\,
            I => \N__29744\
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__29766\,
            I => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__29761\,
            I => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__29756\,
            I => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__29749\,
            I => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\
        );

    \I__6006\ : Odrv4
    port map (
            O => \N__29744\,
            I => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\
        );

    \I__6005\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29730\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__29730\,
            I => \N__29726\
        );

    \I__6003\ : InMux
    port map (
            O => \N__29729\,
            I => \N__29723\
        );

    \I__6002\ : Span4Mux_s3_v
    port map (
            O => \N__29726\,
            I => \N__29718\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__29723\,
            I => \N__29718\
        );

    \I__6000\ : Span4Mux_h
    port map (
            O => \N__29718\,
            I => \N__29715\
        );

    \I__5999\ : Span4Mux_h
    port map (
            O => \N__29715\,
            I => \N__29712\
        );

    \I__5998\ : Odrv4
    port map (
            O => \N__29712\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__5997\ : InMux
    port map (
            O => \N__29709\,
            I => \N__29706\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__29706\,
            I => \N__29703\
        );

    \I__5995\ : Span4Mux_v
    port map (
            O => \N__29703\,
            I => \N__29700\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__29700\,
            I => \POWERLED.count_0_4\
        );

    \I__5993\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29693\
        );

    \I__5992\ : InMux
    port map (
            O => \N__29696\,
            I => \N__29690\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__29693\,
            I => \N__29687\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__29690\,
            I => \POWERLED.count_1_4\
        );

    \I__5989\ : Odrv4
    port map (
            O => \N__29687\,
            I => \POWERLED.count_1_4\
        );

    \I__5988\ : CascadeMux
    port map (
            O => \N__29682\,
            I => \POWERLED.curr_stateZ0Z_0_cascade_\
        );

    \I__5987\ : CascadeMux
    port map (
            O => \N__29679\,
            I => \POWERLED.count_0_sqmuxa_i_cascade_\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \POWERLED.count_1_0_cascade_\
        );

    \I__5985\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \POWERLED.count_1_1_cascade_\
        );

    \I__5984\ : CascadeMux
    port map (
            O => \N__29670\,
            I => \POWERLED.countZ0Z_1_cascade_\
        );

    \I__5983\ : InMux
    port map (
            O => \N__29667\,
            I => \N__29664\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__29664\,
            I => \POWERLED.count_0_1\
        );

    \I__5981\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29642\
        );

    \I__5980\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29637\
        );

    \I__5979\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29637\
        );

    \I__5978\ : InMux
    port map (
            O => \N__29658\,
            I => \N__29628\
        );

    \I__5977\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29628\
        );

    \I__5976\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29628\
        );

    \I__5975\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29628\
        );

    \I__5974\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29621\
        );

    \I__5973\ : InMux
    port map (
            O => \N__29653\,
            I => \N__29621\
        );

    \I__5972\ : InMux
    port map (
            O => \N__29652\,
            I => \N__29621\
        );

    \I__5971\ : InMux
    port map (
            O => \N__29651\,
            I => \N__29614\
        );

    \I__5970\ : InMux
    port map (
            O => \N__29650\,
            I => \N__29614\
        );

    \I__5969\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29614\
        );

    \I__5968\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29605\
        );

    \I__5967\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29605\
        );

    \I__5966\ : InMux
    port map (
            O => \N__29646\,
            I => \N__29605\
        );

    \I__5965\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29605\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__29642\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__29637\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__29628\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__29621\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__29614\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__29605\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__5958\ : InMux
    port map (
            O => \N__29592\,
            I => \N__29589\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__29589\,
            I => \POWERLED.count_0_0\
        );

    \I__5956\ : CascadeMux
    port map (
            O => \N__29586\,
            I => \N__29583\
        );

    \I__5955\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29577\
        );

    \I__5954\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29577\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__29577\,
            I => \POWERLED.count_1_10\
        );

    \I__5952\ : InMux
    port map (
            O => \N__29574\,
            I => \N__29571\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__29571\,
            I => \POWERLED.count_0_10\
        );

    \I__5950\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29565\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__29565\,
            I => \DSW_PWRGD.count_rst_6\
        );

    \I__5948\ : CascadeMux
    port map (
            O => \N__29562\,
            I => \DSW_PWRGD.un2_count_1_axb_8_cascade_\
        );

    \I__5947\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29553\
        );

    \I__5946\ : InMux
    port map (
            O => \N__29558\,
            I => \N__29553\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__29553\,
            I => \DSW_PWRGD.count_1_8\
        );

    \I__5944\ : InMux
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__29547\,
            I => \DSW_PWRGD.un12_clk_100khz_13\
        );

    \I__5942\ : CascadeMux
    port map (
            O => \N__29544\,
            I => \DSW_PWRGD.N_1_i_cascade_\
        );

    \I__5941\ : InMux
    port map (
            O => \N__29541\,
            I => \N__29538\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__5939\ : Odrv4
    port map (
            O => \N__29535\,
            I => \DSW_PWRGD.count_1_10\
        );

    \I__5938\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \POWERLED.g0_i_o3_0_cascade_\
        );

    \I__5937\ : SRMux
    port map (
            O => \N__29529\,
            I => \N__29526\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__29520\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__5933\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29511\
        );

    \I__5932\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29511\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__29511\,
            I => \POWERLED.N_8\
        );

    \I__5930\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29502\
        );

    \I__5929\ : InMux
    port map (
            O => \N__29507\,
            I => \N__29502\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__29502\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__5927\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29496\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__29496\,
            I => \POWERLED.g0_i_o3_0\
        );

    \I__5925\ : IoInMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__29490\,
            I => \N__29487\
        );

    \I__5923\ : Span4Mux_s1_v
    port map (
            O => \N__29487\,
            I => \N__29484\
        );

    \I__5922\ : Sp12to4
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__5921\ : Span12Mux_s8_h
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__5920\ : Odrv12
    port map (
            O => \N__29478\,
            I => pwrbtn_led
        );

    \I__5919\ : CascadeMux
    port map (
            O => \N__29475\,
            I => \POWERLED.curr_state_3_0_cascade_\
        );

    \I__5918\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29466\
        );

    \I__5917\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29466\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__29466\,
            I => \DSW_PWRGD.count_1_5\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__29463\,
            I => \DSW_PWRGD.count_rst_4_cascade_\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__5913\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29451\
        );

    \I__5912\ : InMux
    port map (
            O => \N__29456\,
            I => \N__29451\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__29451\,
            I => \N__29448\
        );

    \I__5910\ : Span4Mux_v
    port map (
            O => \N__29448\,
            I => \N__29445\
        );

    \I__5909\ : Span4Mux_h
    port map (
            O => \N__29445\,
            I => \N__29441\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__29444\,
            I => \N__29438\
        );

    \I__5907\ : Span4Mux_h
    port map (
            O => \N__29441\,
            I => \N__29434\
        );

    \I__5906\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29429\
        );

    \I__5905\ : InMux
    port map (
            O => \N__29437\,
            I => \N__29429\
        );

    \I__5904\ : Span4Mux_v
    port map (
            O => \N__29434\,
            I => \N__29424\
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__29429\,
            I => \N__29424\
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__29424\,
            I => \VPP_VDDQ.N_3160_i\
        );

    \I__5901\ : CascadeMux
    port map (
            O => \N__29421\,
            I => \DSW_PWRGD.count_rst_6_cascade_\
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__29418\,
            I => \DSW_PWRGD.un12_clk_100khz_6_cascade_\
        );

    \I__5899\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__5897\ : Odrv12
    port map (
            O => \N__29409\,
            I => \DSW_PWRGD.un12_clk_100khz_5\
        );

    \I__5896\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29403\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__29403\,
            I => \N__29399\
        );

    \I__5894\ : InMux
    port map (
            O => \N__29402\,
            I => \N__29396\
        );

    \I__5893\ : Span4Mux_h
    port map (
            O => \N__29399\,
            I => \N__29393\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__29396\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__5891\ : Odrv4
    port map (
            O => \N__29393\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__5890\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29385\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__29385\,
            I => \N__29381\
        );

    \I__5888\ : InMux
    port map (
            O => \N__29384\,
            I => \N__29378\
        );

    \I__5887\ : Span4Mux_h
    port map (
            O => \N__29381\,
            I => \N__29375\
        );

    \I__5886\ : LocalMux
    port map (
            O => \N__29378\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__5885\ : Odrv4
    port map (
            O => \N__29375\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__29370\,
            I => \N__29367\
        );

    \I__5883\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29364\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__29364\,
            I => \N__29360\
        );

    \I__5881\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29357\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__29360\,
            I => \N__29354\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__29357\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__5878\ : Odrv4
    port map (
            O => \N__29354\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__5877\ : InMux
    port map (
            O => \N__29349\,
            I => \N__29346\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__29346\,
            I => \N__29342\
        );

    \I__5875\ : InMux
    port map (
            O => \N__29345\,
            I => \N__29339\
        );

    \I__5874\ : Span4Mux_v
    port map (
            O => \N__29342\,
            I => \N__29336\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__29339\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__5872\ : Odrv4
    port map (
            O => \N__29336\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__5870\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29325\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__29325\,
            I => \N__29322\
        );

    \I__5868\ : Odrv12
    port map (
            O => \N__29322\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__5867\ : CascadeMux
    port map (
            O => \N__29319\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\
        );

    \I__5866\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29310\
        );

    \I__5865\ : InMux
    port map (
            O => \N__29315\,
            I => \N__29310\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__5863\ : Span4Mux_h
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__5862\ : Span4Mux_h
    port map (
            O => \N__29304\,
            I => \N__29300\
        );

    \I__5861\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29297\
        );

    \I__5860\ : Sp12to4
    port map (
            O => \N__29300\,
            I => \N__29294\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__29297\,
            I => \VPP_VDDQ.N_3140_i\
        );

    \I__5858\ : Odrv12
    port map (
            O => \N__29294\,
            I => \VPP_VDDQ.N_3140_i\
        );

    \I__5857\ : InMux
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__29286\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__5855\ : InMux
    port map (
            O => \N__29283\,
            I => \N__29277\
        );

    \I__5854\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29277\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__29277\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__5852\ : InMux
    port map (
            O => \N__29274\,
            I => \N__29265\
        );

    \I__5851\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29265\
        );

    \I__5850\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29262\
        );

    \I__5849\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29257\
        );

    \I__5848\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29257\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__29265\,
            I => \N__29254\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29251\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29248\
        );

    \I__5844\ : Span4Mux_s3_v
    port map (
            O => \N__29254\,
            I => \N__29245\
        );

    \I__5843\ : Span4Mux_v
    port map (
            O => \N__29251\,
            I => \N__29242\
        );

    \I__5842\ : Sp12to4
    port map (
            O => \N__29248\,
            I => \N__29239\
        );

    \I__5841\ : Sp12to4
    port map (
            O => \N__29245\,
            I => \N__29236\
        );

    \I__5840\ : Span4Mux_v
    port map (
            O => \N__29242\,
            I => \N__29233\
        );

    \I__5839\ : Span12Mux_v
    port map (
            O => \N__29239\,
            I => \N__29230\
        );

    \I__5838\ : Span12Mux_v
    port map (
            O => \N__29236\,
            I => \N__29227\
        );

    \I__5837\ : Span4Mux_h
    port map (
            O => \N__29233\,
            I => \N__29224\
        );

    \I__5836\ : Odrv12
    port map (
            O => \N__29230\,
            I => vddq_ok
        );

    \I__5835\ : Odrv12
    port map (
            O => \N__29227\,
            I => vddq_ok
        );

    \I__5834\ : Odrv4
    port map (
            O => \N__29224\,
            I => vddq_ok
        );

    \I__5833\ : CascadeMux
    port map (
            O => \N__29217\,
            I => \N__29214\
        );

    \I__5832\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29208\
        );

    \I__5831\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29208\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__29208\,
            I => \N__29203\
        );

    \I__5829\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29198\
        );

    \I__5828\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29198\
        );

    \I__5827\ : Odrv12
    port map (
            O => \N__29203\,
            I => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__29198\,
            I => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\
        );

    \I__5825\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29189\
        );

    \I__5824\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29186\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__29186\,
            I => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\
        );

    \I__5821\ : Odrv4
    port map (
            O => \N__29183\,
            I => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\
        );

    \I__5820\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29175\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__29175\,
            I => \VPP_VDDQ.curr_state_2_0_1\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__29172\,
            I => \DSW_PWRGD.count_rst_7_cascade_\
        );

    \I__5817\ : CascadeMux
    port map (
            O => \N__29169\,
            I => \DSW_PWRGD.un2_count_1_axb_5_cascade_\
        );

    \I__5816\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__29163\,
            I => \DSW_PWRGD.count_rst_9\
        );

    \I__5814\ : CascadeMux
    port map (
            O => \N__29160\,
            I => \DSW_PWRGD.count_rst_9_cascade_\
        );

    \I__5813\ : InMux
    port map (
            O => \N__29157\,
            I => \N__29153\
        );

    \I__5812\ : CascadeMux
    port map (
            O => \N__29156\,
            I => \N__29148\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__29153\,
            I => \N__29138\
        );

    \I__5810\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29133\
        );

    \I__5809\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29133\
        );

    \I__5808\ : InMux
    port map (
            O => \N__29148\,
            I => \N__29130\
        );

    \I__5807\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29125\
        );

    \I__5806\ : InMux
    port map (
            O => \N__29146\,
            I => \N__29125\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__29145\,
            I => \N__29113\
        );

    \I__5804\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29105\
        );

    \I__5803\ : InMux
    port map (
            O => \N__29143\,
            I => \N__29105\
        );

    \I__5802\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29105\
        );

    \I__5801\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29102\
        );

    \I__5800\ : Span4Mux_v
    port map (
            O => \N__29138\,
            I => \N__29092\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__29133\,
            I => \N__29092\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__29130\,
            I => \N__29092\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__29125\,
            I => \N__29092\
        );

    \I__5796\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29088\
        );

    \I__5795\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29083\
        );

    \I__5794\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29083\
        );

    \I__5793\ : InMux
    port map (
            O => \N__29121\,
            I => \N__29075\
        );

    \I__5792\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29075\
        );

    \I__5791\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29075\
        );

    \I__5790\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29068\
        );

    \I__5789\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29068\
        );

    \I__5788\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29068\
        );

    \I__5787\ : InMux
    port map (
            O => \N__29113\,
            I => \N__29063\
        );

    \I__5786\ : InMux
    port map (
            O => \N__29112\,
            I => \N__29063\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29058\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__29102\,
            I => \N__29058\
        );

    \I__5783\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29055\
        );

    \I__5782\ : IoSpan4Mux
    port map (
            O => \N__29092\,
            I => \N__29052\
        );

    \I__5781\ : InMux
    port map (
            O => \N__29091\,
            I => \N__29049\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__29088\,
            I => \N__29041\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__29083\,
            I => \N__29041\
        );

    \I__5778\ : InMux
    port map (
            O => \N__29082\,
            I => \N__29038\
        );

    \I__5777\ : LocalMux
    port map (
            O => \N__29075\,
            I => \N__29031\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29031\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29031\
        );

    \I__5774\ : Span4Mux_s3_v
    port map (
            O => \N__29058\,
            I => \N__29028\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__29055\,
            I => \N__29023\
        );

    \I__5772\ : IoSpan4Mux
    port map (
            O => \N__29052\,
            I => \N__29023\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__29020\
        );

    \I__5770\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29013\
        );

    \I__5769\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29013\
        );

    \I__5768\ : InMux
    port map (
            O => \N__29046\,
            I => \N__29013\
        );

    \I__5767\ : Span12Mux_s6_v
    port map (
            O => \N__29041\,
            I => \N__29010\
        );

    \I__5766\ : LocalMux
    port map (
            O => \N__29038\,
            I => \N__28997\
        );

    \I__5765\ : Span4Mux_s3_v
    port map (
            O => \N__29031\,
            I => \N__28997\
        );

    \I__5764\ : Span4Mux_h
    port map (
            O => \N__29028\,
            I => \N__28997\
        );

    \I__5763\ : Span4Mux_s1_h
    port map (
            O => \N__29023\,
            I => \N__28997\
        );

    \I__5762\ : Span4Mux_h
    port map (
            O => \N__29020\,
            I => \N__28997\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__29013\,
            I => \N__28997\
        );

    \I__5760\ : Odrv12
    port map (
            O => \N__29010\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5759\ : Odrv4
    port map (
            O => \N__28997\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__28992\,
            I => \POWERLED.un1_i3_mux_cascade_\
        );

    \I__5757\ : InMux
    port map (
            O => \N__28989\,
            I => \N__28986\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__28986\,
            I => \POWERLED.d_i3_mux\
        );

    \I__5755\ : InMux
    port map (
            O => \N__28983\,
            I => \N__28980\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__28980\,
            I => \N__28977\
        );

    \I__5753\ : Span4Mux_v
    port map (
            O => \N__28977\,
            I => \N__28974\
        );

    \I__5752\ : Odrv4
    port map (
            O => \N__28974\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_5\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__28971\,
            I => \N__28963\
        );

    \I__5750\ : CascadeMux
    port map (
            O => \N__28970\,
            I => \N__28960\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__28969\,
            I => \N__28956\
        );

    \I__5748\ : InMux
    port map (
            O => \N__28968\,
            I => \N__28951\
        );

    \I__5747\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28951\
        );

    \I__5746\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28948\
        );

    \I__5745\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28945\
        );

    \I__5744\ : InMux
    port map (
            O => \N__28960\,
            I => \N__28942\
        );

    \I__5743\ : InMux
    port map (
            O => \N__28959\,
            I => \N__28937\
        );

    \I__5742\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28937\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__28951\,
            I => \N__28934\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__28948\,
            I => \N__28931\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28924\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__28942\,
            I => \N__28921\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__28937\,
            I => \N__28916\
        );

    \I__5736\ : Span4Mux_s3_v
    port map (
            O => \N__28934\,
            I => \N__28916\
        );

    \I__5735\ : Span4Mux_s3_v
    port map (
            O => \N__28931\,
            I => \N__28913\
        );

    \I__5734\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28908\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28908\
        );

    \I__5732\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28905\
        );

    \I__5731\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28902\
        );

    \I__5730\ : Span4Mux_v
    port map (
            O => \N__28924\,
            I => \N__28895\
        );

    \I__5729\ : Span4Mux_h
    port map (
            O => \N__28921\,
            I => \N__28895\
        );

    \I__5728\ : Span4Mux_h
    port map (
            O => \N__28916\,
            I => \N__28895\
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__28913\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__28908\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__28905\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__28902\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__28895\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__5722\ : CascadeMux
    port map (
            O => \N__28884\,
            I => \N__28881\
        );

    \I__5721\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28878\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28875\
        );

    \I__5719\ : Span4Mux_h
    port map (
            O => \N__28875\,
            I => \N__28872\
        );

    \I__5718\ : Odrv4
    port map (
            O => \N__28872\,
            I => \POWERLED.dutycycle_RNIZ0Z_5\
        );

    \I__5717\ : CascadeMux
    port map (
            O => \N__28869\,
            I => \N__28860\
        );

    \I__5716\ : CascadeMux
    port map (
            O => \N__28868\,
            I => \N__28857\
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__28867\,
            I => \N__28851\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__28866\,
            I => \N__28848\
        );

    \I__5713\ : CascadeMux
    port map (
            O => \N__28865\,
            I => \N__28843\
        );

    \I__5712\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28833\
        );

    \I__5711\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28833\
        );

    \I__5710\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28828\
        );

    \I__5709\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28823\
        );

    \I__5708\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28823\
        );

    \I__5707\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28820\
        );

    \I__5706\ : InMux
    port map (
            O => \N__28854\,
            I => \N__28817\
        );

    \I__5705\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28814\
        );

    \I__5704\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28811\
        );

    \I__5703\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28806\
        );

    \I__5702\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28806\
        );

    \I__5701\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28803\
        );

    \I__5700\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28796\
        );

    \I__5699\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28796\
        );

    \I__5698\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28796\
        );

    \I__5697\ : InMux
    port map (
            O => \N__28839\,
            I => \N__28791\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__28838\,
            I => \N__28788\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__28833\,
            I => \N__28782\
        );

    \I__5694\ : InMux
    port map (
            O => \N__28832\,
            I => \N__28777\
        );

    \I__5693\ : InMux
    port map (
            O => \N__28831\,
            I => \N__28777\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__28828\,
            I => \N__28772\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__28823\,
            I => \N__28772\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__28820\,
            I => \N__28769\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__28817\,
            I => \N__28766\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__28814\,
            I => \N__28763\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__28811\,
            I => \N__28756\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__28806\,
            I => \N__28756\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28756\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__28796\,
            I => \N__28753\
        );

    \I__5683\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28750\
        );

    \I__5682\ : CascadeMux
    port map (
            O => \N__28794\,
            I => \N__28747\
        );

    \I__5681\ : LocalMux
    port map (
            O => \N__28791\,
            I => \N__28744\
        );

    \I__5680\ : InMux
    port map (
            O => \N__28788\,
            I => \N__28741\
        );

    \I__5679\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28734\
        );

    \I__5678\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28734\
        );

    \I__5677\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28734\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__28782\,
            I => \N__28727\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28727\
        );

    \I__5674\ : Span4Mux_h
    port map (
            O => \N__28772\,
            I => \N__28727\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__28769\,
            I => \N__28720\
        );

    \I__5672\ : Span4Mux_s3_h
    port map (
            O => \N__28766\,
            I => \N__28720\
        );

    \I__5671\ : Span4Mux_s3_h
    port map (
            O => \N__28763\,
            I => \N__28720\
        );

    \I__5670\ : Span4Mux_h
    port map (
            O => \N__28756\,
            I => \N__28713\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__28753\,
            I => \N__28713\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__28750\,
            I => \N__28713\
        );

    \I__5667\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28710\
        );

    \I__5666\ : Odrv4
    port map (
            O => \N__28744\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__28741\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__28734\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__28727\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5662\ : Odrv4
    port map (
            O => \N__28720\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__28713\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__28710\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__5659\ : CascadeMux
    port map (
            O => \N__28695\,
            I => \N__28691\
        );

    \I__5658\ : InMux
    port map (
            O => \N__28694\,
            I => \N__28685\
        );

    \I__5657\ : InMux
    port map (
            O => \N__28691\,
            I => \N__28682\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__28690\,
            I => \N__28679\
        );

    \I__5655\ : InMux
    port map (
            O => \N__28689\,
            I => \N__28671\
        );

    \I__5654\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28668\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__28685\,
            I => \N__28663\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28663\
        );

    \I__5651\ : InMux
    port map (
            O => \N__28679\,
            I => \N__28660\
        );

    \I__5650\ : InMux
    port map (
            O => \N__28678\,
            I => \N__28651\
        );

    \I__5649\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28651\
        );

    \I__5648\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28651\
        );

    \I__5647\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28651\
        );

    \I__5646\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28646\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__28671\,
            I => \N__28643\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28636\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__28663\,
            I => \N__28636\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__28660\,
            I => \N__28636\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28633\
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__28650\,
            I => \N__28628\
        );

    \I__5639\ : InMux
    port map (
            O => \N__28649\,
            I => \N__28625\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28622\
        );

    \I__5637\ : Span4Mux_v
    port map (
            O => \N__28643\,
            I => \N__28617\
        );

    \I__5636\ : Span4Mux_v
    port map (
            O => \N__28636\,
            I => \N__28617\
        );

    \I__5635\ : Span4Mux_v
    port map (
            O => \N__28633\,
            I => \N__28614\
        );

    \I__5634\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28609\
        );

    \I__5633\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28609\
        );

    \I__5632\ : InMux
    port map (
            O => \N__28628\,
            I => \N__28606\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__28625\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5630\ : Odrv4
    port map (
            O => \N__28622\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5629\ : Odrv4
    port map (
            O => \N__28617\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__28614\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__28609\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__28606\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__28593\,
            I => \N__28583\
        );

    \I__5624\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28575\
        );

    \I__5623\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28575\
        );

    \I__5622\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28575\
        );

    \I__5621\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28570\
        );

    \I__5620\ : InMux
    port map (
            O => \N__28588\,
            I => \N__28566\
        );

    \I__5619\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28563\
        );

    \I__5618\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28553\
        );

    \I__5617\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28553\
        );

    \I__5616\ : InMux
    port map (
            O => \N__28582\,
            I => \N__28553\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__28575\,
            I => \N__28550\
        );

    \I__5614\ : CascadeMux
    port map (
            O => \N__28574\,
            I => \N__28547\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__28573\,
            I => \N__28544\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__28570\,
            I => \N__28541\
        );

    \I__5611\ : CascadeMux
    port map (
            O => \N__28569\,
            I => \N__28538\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28535\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__28563\,
            I => \N__28532\
        );

    \I__5608\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28525\
        );

    \I__5607\ : InMux
    port map (
            O => \N__28561\,
            I => \N__28525\
        );

    \I__5606\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28525\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__28553\,
            I => \N__28522\
        );

    \I__5604\ : Span4Mux_v
    port map (
            O => \N__28550\,
            I => \N__28519\
        );

    \I__5603\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28516\
        );

    \I__5602\ : InMux
    port map (
            O => \N__28544\,
            I => \N__28513\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__28541\,
            I => \N__28510\
        );

    \I__5600\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28507\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__28535\,
            I => \N__28494\
        );

    \I__5598\ : Span4Mux_h
    port map (
            O => \N__28532\,
            I => \N__28494\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__28525\,
            I => \N__28494\
        );

    \I__5596\ : Span4Mux_h
    port map (
            O => \N__28522\,
            I => \N__28494\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__28519\,
            I => \N__28494\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__28516\,
            I => \N__28494\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__28513\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__28510\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__28507\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__28494\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__5588\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28479\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__28479\,
            I => \N__28475\
        );

    \I__5586\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28472\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__28475\,
            I => \N__28469\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__28472\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_3\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__28469\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_3\
        );

    \I__5582\ : CascadeMux
    port map (
            O => \N__28464\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__5581\ : CascadeMux
    port map (
            O => \N__28461\,
            I => \VPP_VDDQ.N_3140_i_cascade_\
        );

    \I__5580\ : InMux
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__28455\,
            I => \VPP_VDDQ.m4_0\
        );

    \I__5578\ : CascadeMux
    port map (
            O => \N__28452\,
            I => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0_cascade_\
        );

    \I__5577\ : CascadeMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__5576\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28443\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__28443\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__5574\ : InMux
    port map (
            O => \N__28440\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__5573\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__28434\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__5571\ : InMux
    port map (
            O => \N__28431\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__5570\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28425\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__28425\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__5568\ : InMux
    port map (
            O => \N__28422\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__28419\,
            I => \N__28416\
        );

    \I__5566\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28413\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__28413\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__5564\ : InMux
    port map (
            O => \N__28410\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__28407\,
            I => \N__28403\
        );

    \I__5562\ : InMux
    port map (
            O => \N__28406\,
            I => \N__28398\
        );

    \I__5561\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28391\
        );

    \I__5560\ : InMux
    port map (
            O => \N__28402\,
            I => \N__28391\
        );

    \I__5559\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28391\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__28398\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__28391\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__5556\ : CascadeMux
    port map (
            O => \N__28386\,
            I => \N__28382\
        );

    \I__5555\ : CascadeMux
    port map (
            O => \N__28385\,
            I => \N__28378\
        );

    \I__5554\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28371\
        );

    \I__5553\ : InMux
    port map (
            O => \N__28381\,
            I => \N__28371\
        );

    \I__5552\ : InMux
    port map (
            O => \N__28378\,
            I => \N__28371\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__28371\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__5550\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__28365\,
            I => \N__28361\
        );

    \I__5548\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28358\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__28361\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__28358\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__5545\ : CascadeMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__5544\ : InMux
    port map (
            O => \N__28350\,
            I => \N__28347\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__28347\,
            I => \POWERLED.un1_dutycycle_53_axb_3_1_0\
        );

    \I__5542\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__28341\,
            I => \N__28338\
        );

    \I__5540\ : Odrv4
    port map (
            O => \N__28338\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__5539\ : CascadeMux
    port map (
            O => \N__28335\,
            I => \N__28332\
        );

    \I__5538\ : InMux
    port map (
            O => \N__28332\,
            I => \N__28329\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__28329\,
            I => \N__28324\
        );

    \I__5536\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28321\
        );

    \I__5535\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28318\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__28324\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__28321\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__28318\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__5531\ : InMux
    port map (
            O => \N__28311\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__28308\,
            I => \N__28305\
        );

    \I__5529\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28302\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__28302\,
            I => \N__28299\
        );

    \I__5527\ : Odrv4
    port map (
            O => \N__28299\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__5526\ : InMux
    port map (
            O => \N__28296\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__5525\ : InMux
    port map (
            O => \N__28293\,
            I => \N__28288\
        );

    \I__5524\ : InMux
    port map (
            O => \N__28292\,
            I => \N__28285\
        );

    \I__5523\ : InMux
    port map (
            O => \N__28291\,
            I => \N__28282\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__28288\,
            I => \N__28275\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__28285\,
            I => \N__28275\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28275\
        );

    \I__5519\ : Odrv12
    port map (
            O => \N__28275\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__28272\,
            I => \N__28269\
        );

    \I__5517\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__28266\,
            I => \N__28263\
        );

    \I__5515\ : Odrv4
    port map (
            O => \N__28263\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__5514\ : InMux
    port map (
            O => \N__28260\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__5513\ : InMux
    port map (
            O => \N__28257\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__5512\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28247\
        );

    \I__5510\ : InMux
    port map (
            O => \N__28250\,
            I => \N__28244\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__28247\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__28244\,
            I => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__5507\ : CascadeMux
    port map (
            O => \N__28239\,
            I => \N__28235\
        );

    \I__5506\ : InMux
    port map (
            O => \N__28238\,
            I => \N__28232\
        );

    \I__5505\ : InMux
    port map (
            O => \N__28235\,
            I => \N__28229\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__28232\,
            I => \N__28226\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__28229\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__28226\,
            I => \POWERLED.mult1_un40_sum_i_5\
        );

    \I__5501\ : InMux
    port map (
            O => \N__28221\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__5500\ : InMux
    port map (
            O => \N__28218\,
            I => \N__28211\
        );

    \I__5499\ : InMux
    port map (
            O => \N__28217\,
            I => \N__28211\
        );

    \I__5498\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28208\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__28211\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__28208\,
            I => \POWERLED.mult1_un47_sum_s_6\
        );

    \I__5495\ : CascadeMux
    port map (
            O => \N__28203\,
            I => \N__28200\
        );

    \I__5494\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__28197\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__5492\ : InMux
    port map (
            O => \N__28194\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__5491\ : CascadeMux
    port map (
            O => \N__28191\,
            I => \N__28188\
        );

    \I__5490\ : InMux
    port map (
            O => \N__28188\,
            I => \N__28185\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__28185\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__5488\ : InMux
    port map (
            O => \N__28182\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__5487\ : InMux
    port map (
            O => \N__28179\,
            I => \N__28173\
        );

    \I__5486\ : InMux
    port map (
            O => \N__28178\,
            I => \N__28173\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__5484\ : Span4Mux_h
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__5483\ : Span4Mux_v
    port map (
            O => \N__28167\,
            I => \N__28164\
        );

    \I__5482\ : Odrv4
    port map (
            O => \N__28164\,
            I => \POWERLED.count_off_1_7\
        );

    \I__5481\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28158\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__28158\,
            I => \POWERLED.count_off_0_7\
        );

    \I__5479\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28152\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__28152\,
            I => \N__28148\
        );

    \I__5477\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28145\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__28148\,
            I => \N__28140\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__28145\,
            I => \N__28140\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__28140\,
            I => \N__28137\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__28134\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__5471\ : InMux
    port map (
            O => \N__28131\,
            I => \N__28125\
        );

    \I__5470\ : InMux
    port map (
            O => \N__28130\,
            I => \N__28125\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__5468\ : Span12Mux_s7_h
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__5467\ : Odrv12
    port map (
            O => \N__28119\,
            I => \POWERLED.count_off_1_8\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__28116\,
            I => \N__28113\
        );

    \I__5465\ : InMux
    port map (
            O => \N__28113\,
            I => \N__28110\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__28110\,
            I => \POWERLED.count_off_0_8\
        );

    \I__5463\ : CEMux
    port map (
            O => \N__28107\,
            I => \N__28100\
        );

    \I__5462\ : InMux
    port map (
            O => \N__28106\,
            I => \N__28090\
        );

    \I__5461\ : InMux
    port map (
            O => \N__28105\,
            I => \N__28090\
        );

    \I__5460\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28090\
        );

    \I__5459\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28090\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__28100\,
            I => \N__28077\
        );

    \I__5457\ : CEMux
    port map (
            O => \N__28099\,
            I => \N__28074\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__28090\,
            I => \N__28071\
        );

    \I__5455\ : CEMux
    port map (
            O => \N__28089\,
            I => \N__28065\
        );

    \I__5454\ : CascadeMux
    port map (
            O => \N__28088\,
            I => \N__28062\
        );

    \I__5453\ : CEMux
    port map (
            O => \N__28087\,
            I => \N__28059\
        );

    \I__5452\ : CEMux
    port map (
            O => \N__28086\,
            I => \N__28056\
        );

    \I__5451\ : CEMux
    port map (
            O => \N__28085\,
            I => \N__28053\
        );

    \I__5450\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28050\
        );

    \I__5449\ : InMux
    port map (
            O => \N__28083\,
            I => \N__28045\
        );

    \I__5448\ : InMux
    port map (
            O => \N__28082\,
            I => \N__28045\
        );

    \I__5447\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28036\
        );

    \I__5446\ : CEMux
    port map (
            O => \N__28080\,
            I => \N__28036\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__28077\,
            I => \N__28033\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__28074\,
            I => \N__28028\
        );

    \I__5443\ : Span4Mux_v
    port map (
            O => \N__28071\,
            I => \N__28028\
        );

    \I__5442\ : InMux
    port map (
            O => \N__28070\,
            I => \N__28021\
        );

    \I__5441\ : InMux
    port map (
            O => \N__28069\,
            I => \N__28021\
        );

    \I__5440\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28021\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__28065\,
            I => \N__28018\
        );

    \I__5438\ : InMux
    port map (
            O => \N__28062\,
            I => \N__28015\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__28059\,
            I => \N__28004\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__28056\,
            I => \N__28004\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__28053\,
            I => \N__28004\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__28050\,
            I => \N__28004\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__28045\,
            I => \N__28004\
        );

    \I__5432\ : InMux
    port map (
            O => \N__28044\,
            I => \N__27999\
        );

    \I__5431\ : InMux
    port map (
            O => \N__28043\,
            I => \N__27999\
        );

    \I__5430\ : InMux
    port map (
            O => \N__28042\,
            I => \N__27996\
        );

    \I__5429\ : InMux
    port map (
            O => \N__28041\,
            I => \N__27993\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__27984\
        );

    \I__5427\ : Sp12to4
    port map (
            O => \N__28033\,
            I => \N__27984\
        );

    \I__5426\ : Sp12to4
    port map (
            O => \N__28028\,
            I => \N__27984\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__28021\,
            I => \N__27984\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__28018\,
            I => \N__27981\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__28015\,
            I => \N__27974\
        );

    \I__5422\ : Span4Mux_v
    port map (
            O => \N__28004\,
            I => \N__27974\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__27999\,
            I => \N__27974\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__27996\,
            I => \N__27969\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27969\
        );

    \I__5418\ : Span12Mux_s11_h
    port map (
            O => \N__27984\,
            I => \N__27966\
        );

    \I__5417\ : Span4Mux_h
    port map (
            O => \N__27981\,
            I => \N__27961\
        );

    \I__5416\ : Span4Mux_h
    port map (
            O => \N__27974\,
            I => \N__27961\
        );

    \I__5415\ : Span12Mux_s5_v
    port map (
            O => \N__27969\,
            I => \N__27958\
        );

    \I__5414\ : Odrv12
    port map (
            O => \N__27966\,
            I => \POWERLED.dutycycle_RNIBADV5Z0Z_0\
        );

    \I__5413\ : Odrv4
    port map (
            O => \N__27961\,
            I => \POWERLED.dutycycle_RNIBADV5Z0Z_0\
        );

    \I__5412\ : Odrv12
    port map (
            O => \N__27958\,
            I => \POWERLED.dutycycle_RNIBADV5Z0Z_0\
        );

    \I__5411\ : CascadeMux
    port map (
            O => \N__27951\,
            I => \N__27947\
        );

    \I__5410\ : InMux
    port map (
            O => \N__27950\,
            I => \N__27944\
        );

    \I__5409\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27941\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__27944\,
            I => \N__27938\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__27941\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__5406\ : Odrv4
    port map (
            O => \N__27938\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__5405\ : CascadeMux
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__5404\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27927\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__27927\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__5402\ : InMux
    port map (
            O => \N__27924\,
            I => \N__27918\
        );

    \I__5401\ : InMux
    port map (
            O => \N__27923\,
            I => \N__27915\
        );

    \I__5400\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27910\
        );

    \I__5399\ : InMux
    port map (
            O => \N__27921\,
            I => \N__27910\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__27918\,
            I => \N__27907\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__27915\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__27910\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__27907\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__27900\,
            I => \N__27897\
        );

    \I__5393\ : InMux
    port map (
            O => \N__27897\,
            I => \N__27890\
        );

    \I__5392\ : InMux
    port map (
            O => \N__27896\,
            I => \N__27890\
        );

    \I__5391\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27887\
        );

    \I__5390\ : LocalMux
    port map (
            O => \N__27890\,
            I => \N__27884\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__27887\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__5388\ : Odrv4
    port map (
            O => \N__27884\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__27879\,
            I => \N__27876\
        );

    \I__5386\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27873\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__27873\,
            I => \POWERLED.mult1_un47_sum_s_4_sf\
        );

    \I__5384\ : InMux
    port map (
            O => \N__27870\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__5383\ : CascadeMux
    port map (
            O => \N__27867\,
            I => \N__27863\
        );

    \I__5382\ : CascadeMux
    port map (
            O => \N__27866\,
            I => \N__27859\
        );

    \I__5381\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27852\
        );

    \I__5380\ : InMux
    port map (
            O => \N__27862\,
            I => \N__27852\
        );

    \I__5379\ : InMux
    port map (
            O => \N__27859\,
            I => \N__27852\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__27852\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__27849\,
            I => \N__27846\
        );

    \I__5376\ : InMux
    port map (
            O => \N__27846\,
            I => \N__27843\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__27843\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__5374\ : InMux
    port map (
            O => \N__27840\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__5373\ : InMux
    port map (
            O => \N__27837\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__5372\ : InMux
    port map (
            O => \N__27834\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__5371\ : InMux
    port map (
            O => \N__27831\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__5370\ : InMux
    port map (
            O => \N__27828\,
            I => \N__27824\
        );

    \I__5369\ : InMux
    port map (
            O => \N__27827\,
            I => \N__27821\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__27824\,
            I => \N__27818\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__27821\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__5366\ : Odrv4
    port map (
            O => \N__27818\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__27813\,
            I => \N__27810\
        );

    \I__5364\ : InMux
    port map (
            O => \N__27810\,
            I => \N__27807\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__27807\,
            I => \N__27804\
        );

    \I__5362\ : Odrv12
    port map (
            O => \N__27804\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__27801\,
            I => \N__27797\
        );

    \I__5360\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27794\
        );

    \I__5359\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27791\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__27794\,
            I => \N__27788\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__27791\,
            I => \N__27785\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__27788\,
            I => \N__27782\
        );

    \I__5355\ : Span4Mux_h
    port map (
            O => \N__27785\,
            I => \N__27779\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__27782\,
            I => \N__27776\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__27779\,
            I => \N__27773\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__27776\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__5351\ : Odrv4
    port map (
            O => \N__27773\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__5350\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27765\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__27765\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__5348\ : InMux
    port map (
            O => \N__27762\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__5347\ : InMux
    port map (
            O => \N__27759\,
            I => \N__27755\
        );

    \I__5346\ : CascadeMux
    port map (
            O => \N__27758\,
            I => \N__27752\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27746\
        );

    \I__5344\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27739\
        );

    \I__5343\ : InMux
    port map (
            O => \N__27751\,
            I => \N__27739\
        );

    \I__5342\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27739\
        );

    \I__5341\ : InMux
    port map (
            O => \N__27749\,
            I => \N__27736\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__27746\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__27739\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__27736\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__5337\ : CascadeMux
    port map (
            O => \N__27729\,
            I => \N__27725\
        );

    \I__5336\ : InMux
    port map (
            O => \N__27728\,
            I => \N__27717\
        );

    \I__5335\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27717\
        );

    \I__5334\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27717\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__27717\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__5332\ : InMux
    port map (
            O => \N__27714\,
            I => \N__27711\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__27711\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__5330\ : InMux
    port map (
            O => \N__27708\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__5329\ : InMux
    port map (
            O => \N__27705\,
            I => \N__27702\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__27702\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__5327\ : InMux
    port map (
            O => \N__27699\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__5326\ : InMux
    port map (
            O => \N__27696\,
            I => \N__27693\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__27693\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__5324\ : InMux
    port map (
            O => \N__27690\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__27687\,
            I => \N__27684\
        );

    \I__5322\ : InMux
    port map (
            O => \N__27684\,
            I => \N__27681\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__27681\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__5320\ : InMux
    port map (
            O => \N__27678\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__5319\ : InMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__27672\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__5317\ : InMux
    port map (
            O => \N__27669\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__5316\ : InMux
    port map (
            O => \N__27666\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__5315\ : InMux
    port map (
            O => \N__27663\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__27660\,
            I => \N__27656\
        );

    \I__5313\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27650\
        );

    \I__5312\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27643\
        );

    \I__5311\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27643\
        );

    \I__5310\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27643\
        );

    \I__5309\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27640\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__27650\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__27643\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__27640\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__27633\,
            I => \N__27629\
        );

    \I__5304\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27621\
        );

    \I__5303\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27621\
        );

    \I__5302\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27621\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__27621\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__5300\ : InMux
    port map (
            O => \N__27618\,
            I => \N__27615\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__27615\,
            I => \N__27611\
        );

    \I__5298\ : InMux
    port map (
            O => \N__27614\,
            I => \N__27608\
        );

    \I__5297\ : Span4Mux_v
    port map (
            O => \N__27611\,
            I => \N__27605\
        );

    \I__5296\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27602\
        );

    \I__5295\ : Odrv4
    port map (
            O => \N__27605\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__5294\ : Odrv4
    port map (
            O => \N__27602\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__5293\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27594\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__27594\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__5291\ : InMux
    port map (
            O => \N__27591\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__5290\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27585\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__27585\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__5288\ : CascadeMux
    port map (
            O => \N__27582\,
            I => \N__27579\
        );

    \I__5287\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27576\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__27576\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__5285\ : InMux
    port map (
            O => \N__27573\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__27570\,
            I => \N__27567\
        );

    \I__5283\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27564\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__27564\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__5281\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27558\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__27558\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__5279\ : InMux
    port map (
            O => \N__27555\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__5278\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27549\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__27549\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__27546\,
            I => \N__27543\
        );

    \I__5275\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27540\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__27540\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__5273\ : InMux
    port map (
            O => \N__27537\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__5272\ : CascadeMux
    port map (
            O => \N__27534\,
            I => \N__27531\
        );

    \I__5271\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27528\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__27525\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__5268\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27519\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__27519\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__5266\ : InMux
    port map (
            O => \N__27516\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__5265\ : InMux
    port map (
            O => \N__27513\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__5264\ : InMux
    port map (
            O => \N__27510\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__5263\ : CascadeMux
    port map (
            O => \N__27507\,
            I => \N__27503\
        );

    \I__5262\ : InMux
    port map (
            O => \N__27506\,
            I => \N__27495\
        );

    \I__5261\ : InMux
    port map (
            O => \N__27503\,
            I => \N__27495\
        );

    \I__5260\ : InMux
    port map (
            O => \N__27502\,
            I => \N__27495\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__27495\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__5258\ : InMux
    port map (
            O => \N__27492\,
            I => \N__27489\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__27489\,
            I => \N__27485\
        );

    \I__5256\ : InMux
    port map (
            O => \N__27488\,
            I => \N__27482\
        );

    \I__5255\ : Span4Mux_h
    port map (
            O => \N__27485\,
            I => \N__27479\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__27482\,
            I => \N__27476\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__27479\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__5252\ : Odrv12
    port map (
            O => \N__27476\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__27471\,
            I => \N__27468\
        );

    \I__5250\ : InMux
    port map (
            O => \N__27468\,
            I => \N__27465\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__27465\,
            I => \N__27462\
        );

    \I__5248\ : Span4Mux_v
    port map (
            O => \N__27462\,
            I => \N__27459\
        );

    \I__5247\ : Odrv4
    port map (
            O => \N__27459\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__5246\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__27453\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__5244\ : InMux
    port map (
            O => \N__27450\,
            I => \POWERLED.mult1_un110_sum_cry_2_c\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__27447\,
            I => \N__27444\
        );

    \I__5242\ : InMux
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__27441\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__5240\ : InMux
    port map (
            O => \N__27438\,
            I => \POWERLED.mult1_un110_sum_cry_3_c\
        );

    \I__5239\ : InMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__27432\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__5237\ : InMux
    port map (
            O => \N__27429\,
            I => \POWERLED.mult1_un110_sum_cry_4_c\
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__27426\,
            I => \N__27423\
        );

    \I__5235\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27420\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__27420\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__5233\ : InMux
    port map (
            O => \N__27417\,
            I => \POWERLED.mult1_un110_sum_cry_5_c\
        );

    \I__5232\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__27411\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__5230\ : InMux
    port map (
            O => \N__27408\,
            I => \POWERLED.mult1_un110_sum_cry_6_c\
        );

    \I__5229\ : InMux
    port map (
            O => \N__27405\,
            I => \N__27402\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__27402\,
            I => \DSW_PWRGD.curr_state_3_0\
        );

    \I__5227\ : CascadeMux
    port map (
            O => \N__27399\,
            I => \DSW_PWRGD.curr_state_7_0_cascade_\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__27396\,
            I => \DSW_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__27393\,
            I => \N__27390\
        );

    \I__5224\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27387\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__27387\,
            I => \N__27384\
        );

    \I__5222\ : Odrv4
    port map (
            O => \N__27384\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__5221\ : InMux
    port map (
            O => \N__27381\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__5220\ : InMux
    port map (
            O => \N__27378\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__5219\ : InMux
    port map (
            O => \N__27375\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__5218\ : InMux
    port map (
            O => \N__27372\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__5217\ : InMux
    port map (
            O => \N__27369\,
            I => \N__27363\
        );

    \I__5216\ : InMux
    port map (
            O => \N__27368\,
            I => \N__27363\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__27363\,
            I => \POWERLED.count_1_12\
        );

    \I__5214\ : InMux
    port map (
            O => \N__27360\,
            I => \POWERLED.un1_count_cry_11\
        );

    \I__5213\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27353\
        );

    \I__5212\ : InMux
    port map (
            O => \N__27356\,
            I => \N__27350\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__27353\,
            I => \POWERLED.count_1_13\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__27350\,
            I => \POWERLED.count_1_13\
        );

    \I__5209\ : InMux
    port map (
            O => \N__27345\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__5208\ : InMux
    port map (
            O => \N__27342\,
            I => \N__27336\
        );

    \I__5207\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27336\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__27336\,
            I => \POWERLED.count_1_14\
        );

    \I__5205\ : InMux
    port map (
            O => \N__27333\,
            I => \POWERLED.un1_count_cry_13\
        );

    \I__5204\ : InMux
    port map (
            O => \N__27330\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__5203\ : CascadeMux
    port map (
            O => \N__27327\,
            I => \N__27324\
        );

    \I__5202\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27318\
        );

    \I__5201\ : InMux
    port map (
            O => \N__27323\,
            I => \N__27318\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__27318\,
            I => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\
        );

    \I__5199\ : InMux
    port map (
            O => \N__27315\,
            I => \N__27312\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__27312\,
            I => \N__27309\
        );

    \I__5197\ : Odrv12
    port map (
            O => \N__27309\,
            I => \POWERLED.un79_clk_100khzlto15_5\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__27306\,
            I => \DSW_PWRGD.curr_state_7_1_cascade_\
        );

    \I__5195\ : InMux
    port map (
            O => \N__27303\,
            I => \N__27300\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__27300\,
            I => \DSW_PWRGD.curr_state_2_1\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__27297\,
            I => \DSW_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__5192\ : InMux
    port map (
            O => \N__27294\,
            I => \POWERLED.un1_count_cry_3\
        );

    \I__5191\ : CascadeMux
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__5190\ : InMux
    port map (
            O => \N__27288\,
            I => \N__27282\
        );

    \I__5189\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27282\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__27282\,
            I => \POWERLED.count_1_5\
        );

    \I__5187\ : InMux
    port map (
            O => \N__27279\,
            I => \POWERLED.un1_count_cry_4\
        );

    \I__5186\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27272\
        );

    \I__5185\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27269\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__27272\,
            I => \POWERLED.count_1_6\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__27269\,
            I => \POWERLED.count_1_6\
        );

    \I__5182\ : InMux
    port map (
            O => \N__27264\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__27261\,
            I => \N__27257\
        );

    \I__5180\ : InMux
    port map (
            O => \N__27260\,
            I => \N__27252\
        );

    \I__5179\ : InMux
    port map (
            O => \N__27257\,
            I => \N__27252\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__27252\,
            I => \POWERLED.count_1_7\
        );

    \I__5177\ : InMux
    port map (
            O => \N__27249\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__5175\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27237\
        );

    \I__5174\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27237\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__27237\,
            I => \POWERLED.count_1_8\
        );

    \I__5172\ : InMux
    port map (
            O => \N__27234\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__27231\,
            I => \N__27228\
        );

    \I__5170\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27222\
        );

    \I__5169\ : InMux
    port map (
            O => \N__27227\,
            I => \N__27222\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__27222\,
            I => \POWERLED.count_1_9\
        );

    \I__5167\ : InMux
    port map (
            O => \N__27219\,
            I => \bfn_8_6_0_\
        );

    \I__5166\ : InMux
    port map (
            O => \N__27216\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__5165\ : InMux
    port map (
            O => \N__27213\,
            I => \N__27207\
        );

    \I__5164\ : InMux
    port map (
            O => \N__27212\,
            I => \N__27207\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__27207\,
            I => \POWERLED.count_1_11\
        );

    \I__5162\ : InMux
    port map (
            O => \N__27204\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__5161\ : CascadeMux
    port map (
            O => \N__27201\,
            I => \POWERLED.un79_clk_100khzlt6_cascade_\
        );

    \I__5160\ : CascadeMux
    port map (
            O => \N__27198\,
            I => \POWERLED.un79_clk_100khzlto15_7_cascade_\
        );

    \I__5159\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__27192\,
            I => \POWERLED.un79_clk_100khzlto15_3\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__27189\,
            I => \POWERLED.count_RNIZ0Z_8_cascade_\
        );

    \I__5156\ : InMux
    port map (
            O => \N__27186\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__27183\,
            I => \N__27179\
        );

    \I__5154\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27174\
        );

    \I__5153\ : InMux
    port map (
            O => \N__27179\,
            I => \N__27174\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__27174\,
            I => \N__27171\
        );

    \I__5151\ : Odrv4
    port map (
            O => \N__27171\,
            I => \POWERLED.count_1_3\
        );

    \I__5150\ : InMux
    port map (
            O => \N__27168\,
            I => \POWERLED.un1_count_cry_2\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__27165\,
            I => \HDA_STRAP.curr_stateZ0Z_0_cascade_\
        );

    \I__5148\ : InMux
    port map (
            O => \N__27162\,
            I => \N__27159\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__27159\,
            I => \N__27156\
        );

    \I__5146\ : Odrv12
    port map (
            O => \N__27156\,
            I => \HDA_STRAP.N_51\
        );

    \I__5145\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27150\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__27150\,
            I => \HDA_STRAP.N_53\
        );

    \I__5143\ : IoInMux
    port map (
            O => \N__27147\,
            I => \N__27144\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__27144\,
            I => \N__27141\
        );

    \I__5141\ : IoSpan4Mux
    port map (
            O => \N__27141\,
            I => \N__27138\
        );

    \I__5140\ : Span4Mux_s1_v
    port map (
            O => \N__27138\,
            I => \N__27135\
        );

    \I__5139\ : Sp12to4
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__5138\ : Odrv12
    port map (
            O => \N__27132\,
            I => \HDA_STRAP.count_enZ0\
        );

    \I__5137\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27126\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__27126\,
            I => \N__27122\
        );

    \I__5135\ : InMux
    port map (
            O => \N__27125\,
            I => \N__27119\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__27122\,
            I => \N__27116\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__27119\,
            I => \N__27113\
        );

    \I__5132\ : Span4Mux_v
    port map (
            O => \N__27116\,
            I => \N__27110\
        );

    \I__5131\ : Span4Mux_s3_v
    port map (
            O => \N__27113\,
            I => \N__27107\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__27110\,
            I => \N__27104\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__27107\,
            I => \N__27101\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__27104\,
            I => \HDA_STRAP.N_3252_i\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__27101\,
            I => \HDA_STRAP.N_3252_i\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__27096\,
            I => \N_414_cascade_\
        );

    \I__5125\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27083\
        );

    \I__5124\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27083\
        );

    \I__5123\ : InMux
    port map (
            O => \N__27091\,
            I => \N__27083\
        );

    \I__5122\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27080\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27077\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__27080\,
            I => \HDA_STRAP.N_285\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__27077\,
            I => \HDA_STRAP.N_285\
        );

    \I__5118\ : InMux
    port map (
            O => \N__27072\,
            I => \N__27069\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__27069\,
            I => \N__27066\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__27066\,
            I => \N__27061\
        );

    \I__5115\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27056\
        );

    \I__5114\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27056\
        );

    \I__5113\ : Span4Mux_v
    port map (
            O => \N__27061\,
            I => \N__27053\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__27056\,
            I => \N__27050\
        );

    \I__5111\ : Span4Mux_v
    port map (
            O => \N__27053\,
            I => \N__27047\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__27050\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__5109\ : Odrv4
    port map (
            O => \N__27047\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__5108\ : InMux
    port map (
            O => \N__27042\,
            I => \N__27038\
        );

    \I__5107\ : InMux
    port map (
            O => \N__27041\,
            I => \N__27035\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27028\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__27035\,
            I => \N__27028\
        );

    \I__5104\ : InMux
    port map (
            O => \N__27034\,
            I => \N__27023\
        );

    \I__5103\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27023\
        );

    \I__5102\ : Odrv12
    port map (
            O => \N__27028\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__27023\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__5099\ : InMux
    port map (
            O => \N__27015\,
            I => \N__27012\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__27012\,
            I => \N__27009\
        );

    \I__5097\ : Odrv4
    port map (
            O => \N__27009\,
            I => gpio_fpga_soc_1
        );

    \I__5096\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26998\
        );

    \I__5095\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26998\
        );

    \I__5094\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26993\
        );

    \I__5093\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26993\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26990\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__26993\,
            I => \N__26984\
        );

    \I__5090\ : Span4Mux_s1_v
    port map (
            O => \N__26990\,
            I => \N__26981\
        );

    \I__5089\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26974\
        );

    \I__5088\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26974\
        );

    \I__5087\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26974\
        );

    \I__5086\ : Span4Mux_h
    port map (
            O => \N__26984\,
            I => \N__26971\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__26981\,
            I => \N_227\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N_227\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__26971\,
            I => \N_227\
        );

    \I__5082\ : InMux
    port map (
            O => \N__26964\,
            I => \N__26961\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__26961\,
            I => \HDA_STRAP.m6_i_0\
        );

    \I__5080\ : CascadeMux
    port map (
            O => \N__26958\,
            I => \HDA_STRAP.m6_i_0_cascade_\
        );

    \I__5079\ : CascadeMux
    port map (
            O => \N__26955\,
            I => \N__26952\
        );

    \I__5078\ : InMux
    port map (
            O => \N__26952\,
            I => \N__26943\
        );

    \I__5077\ : InMux
    port map (
            O => \N__26951\,
            I => \N__26943\
        );

    \I__5076\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26943\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__26943\,
            I => \N_414\
        );

    \I__5074\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26937\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__26937\,
            I => \HDA_STRAP.curr_state_4_0\
        );

    \I__5072\ : CascadeMux
    port map (
            O => \N__26934\,
            I => \N__26927\
        );

    \I__5071\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26924\
        );

    \I__5070\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26917\
        );

    \I__5069\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26917\
        );

    \I__5068\ : InMux
    port map (
            O => \N__26930\,
            I => \N__26917\
        );

    \I__5067\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26914\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__26924\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__26917\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__26914\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__5063\ : InMux
    port map (
            O => \N__26907\,
            I => \N__26904\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__26904\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__26901\,
            I => \VPP_VDDQ.count_2Z0Z_8_cascade_\
        );

    \I__5060\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26895\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__26895\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__5058\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26886\
        );

    \I__5057\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26886\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__26886\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\
        );

    \I__5055\ : CascadeMux
    port map (
            O => \N__26883\,
            I => \VPP_VDDQ.count_2_rst_3_cascade_\
        );

    \I__5054\ : InMux
    port map (
            O => \N__26880\,
            I => \N__26877\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26874\
        );

    \I__5052\ : Span4Mux_h
    port map (
            O => \N__26874\,
            I => \N__26871\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__26871\,
            I => \VPP_VDDQ.un29_clk_100khz_12\
        );

    \I__5050\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__26865\,
            I => \N__26862\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__26862\,
            I => \VPP_VDDQ.un29_clk_100khz_11\
        );

    \I__5047\ : CascadeMux
    port map (
            O => \N__26859\,
            I => \VPP_VDDQ.un29_clk_100khz_5_cascade_\
        );

    \I__5046\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__26853\,
            I => \VPP_VDDQ.un29_clk_100khz_4\
        );

    \I__5044\ : CascadeMux
    port map (
            O => \N__26850\,
            I => \N__26846\
        );

    \I__5043\ : InMux
    port map (
            O => \N__26849\,
            I => \N__26842\
        );

    \I__5042\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26839\
        );

    \I__5041\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26836\
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__26842\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__26839\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__26836\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__5037\ : InMux
    port map (
            O => \N__26829\,
            I => \N__26823\
        );

    \I__5036\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26823\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__26823\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\
        );

    \I__5034\ : CascadeMux
    port map (
            O => \N__26820\,
            I => \VPP_VDDQ.N_1_i_cascade_\
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__26817\,
            I => \N__26808\
        );

    \I__5032\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26797\
        );

    \I__5031\ : CascadeMux
    port map (
            O => \N__26815\,
            I => \N__26786\
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__26814\,
            I => \N__26778\
        );

    \I__5029\ : SRMux
    port map (
            O => \N__26813\,
            I => \N__26764\
        );

    \I__5028\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26764\
        );

    \I__5027\ : InMux
    port map (
            O => \N__26811\,
            I => \N__26764\
        );

    \I__5026\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26764\
        );

    \I__5025\ : InMux
    port map (
            O => \N__26807\,
            I => \N__26764\
        );

    \I__5024\ : SRMux
    port map (
            O => \N__26806\,
            I => \N__26760\
        );

    \I__5023\ : SRMux
    port map (
            O => \N__26805\,
            I => \N__26749\
        );

    \I__5022\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26749\
        );

    \I__5021\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26749\
        );

    \I__5020\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26749\
        );

    \I__5019\ : InMux
    port map (
            O => \N__26801\,
            I => \N__26749\
        );

    \I__5018\ : SRMux
    port map (
            O => \N__26800\,
            I => \N__26746\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__26797\,
            I => \N__26743\
        );

    \I__5016\ : InMux
    port map (
            O => \N__26796\,
            I => \N__26734\
        );

    \I__5015\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26734\
        );

    \I__5014\ : InMux
    port map (
            O => \N__26794\,
            I => \N__26734\
        );

    \I__5013\ : InMux
    port map (
            O => \N__26793\,
            I => \N__26734\
        );

    \I__5012\ : SRMux
    port map (
            O => \N__26792\,
            I => \N__26731\
        );

    \I__5011\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26728\
        );

    \I__5010\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26725\
        );

    \I__5009\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26718\
        );

    \I__5008\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26718\
        );

    \I__5007\ : InMux
    port map (
            O => \N__26785\,
            I => \N__26718\
        );

    \I__5006\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26713\
        );

    \I__5005\ : InMux
    port map (
            O => \N__26783\,
            I => \N__26713\
        );

    \I__5004\ : SRMux
    port map (
            O => \N__26782\,
            I => \N__26710\
        );

    \I__5003\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26701\
        );

    \I__5002\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26701\
        );

    \I__5001\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26701\
        );

    \I__5000\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26701\
        );

    \I__4999\ : InMux
    port map (
            O => \N__26775\,
            I => \N__26698\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__26764\,
            I => \N__26695\
        );

    \I__4997\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26692\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__26760\,
            I => \N__26687\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__26749\,
            I => \N__26687\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__26746\,
            I => \N__26680\
        );

    \I__4993\ : Span4Mux_s2_v
    port map (
            O => \N__26743\,
            I => \N__26680\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__26734\,
            I => \N__26680\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26677\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__26728\,
            I => \N__26674\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__26725\,
            I => \N__26671\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26666\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__26713\,
            I => \N__26666\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__26710\,
            I => \N__26655\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__26701\,
            I => \N__26655\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__26698\,
            I => \N__26655\
        );

    \I__4983\ : Span4Mux_s1_v
    port map (
            O => \N__26695\,
            I => \N__26655\
        );

    \I__4982\ : LocalMux
    port map (
            O => \N__26692\,
            I => \N__26655\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__26687\,
            I => \N__26652\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__26680\,
            I => \N__26649\
        );

    \I__4979\ : Span4Mux_s1_v
    port map (
            O => \N__26677\,
            I => \N__26644\
        );

    \I__4978\ : Span4Mux_s1_v
    port map (
            O => \N__26674\,
            I => \N__26644\
        );

    \I__4977\ : Span4Mux_s1_v
    port map (
            O => \N__26671\,
            I => \N__26637\
        );

    \I__4976\ : Span4Mux_h
    port map (
            O => \N__26666\,
            I => \N__26637\
        );

    \I__4975\ : Span4Mux_h
    port map (
            O => \N__26655\,
            I => \N__26637\
        );

    \I__4974\ : Span4Mux_v
    port map (
            O => \N__26652\,
            I => \N__26634\
        );

    \I__4973\ : Span4Mux_v
    port map (
            O => \N__26649\,
            I => \N__26631\
        );

    \I__4972\ : Span4Mux_v
    port map (
            O => \N__26644\,
            I => \N__26628\
        );

    \I__4971\ : Span4Mux_v
    port map (
            O => \N__26637\,
            I => \N__26625\
        );

    \I__4970\ : Span4Mux_v
    port map (
            O => \N__26634\,
            I => \N__26622\
        );

    \I__4969\ : Span4Mux_h
    port map (
            O => \N__26631\,
            I => \N__26619\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__26628\,
            I => \N__26616\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__26625\,
            I => \N__26613\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__26622\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__4965\ : Odrv4
    port map (
            O => \N__26619\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__26616\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__26613\,
            I => \VPP_VDDQ.count_2_0_sqmuxa\
        );

    \I__4962\ : InMux
    port map (
            O => \N__26604\,
            I => \N__26601\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__26601\,
            I => \VPP_VDDQ.count_2_rst_0\
        );

    \I__4960\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26592\
        );

    \I__4959\ : InMux
    port map (
            O => \N__26597\,
            I => \N__26592\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__26592\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__4957\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26586\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__26586\,
            I => \VPP_VDDQ.count_2_rst_3\
        );

    \I__4955\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26576\
        );

    \I__4954\ : InMux
    port map (
            O => \N__26582\,
            I => \N__26576\
        );

    \I__4953\ : InMux
    port map (
            O => \N__26581\,
            I => \N__26573\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__26576\,
            I => \VPP_VDDQ.un1_count_2_1_axb_5\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__26573\,
            I => \VPP_VDDQ.un1_count_2_1_axb_5\
        );

    \I__4950\ : CascadeMux
    port map (
            O => \N__26568\,
            I => \N__26562\
        );

    \I__4949\ : CascadeMux
    port map (
            O => \N__26567\,
            I => \N__26556\
        );

    \I__4948\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26550\
        );

    \I__4947\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26545\
        );

    \I__4946\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26545\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__26561\,
            I => \N__26540\
        );

    \I__4944\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26535\
        );

    \I__4943\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26530\
        );

    \I__4942\ : InMux
    port map (
            O => \N__26556\,
            I => \N__26530\
        );

    \I__4941\ : InMux
    port map (
            O => \N__26555\,
            I => \N__26523\
        );

    \I__4940\ : InMux
    port map (
            O => \N__26554\,
            I => \N__26523\
        );

    \I__4939\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26523\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__26550\,
            I => \N__26518\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__26545\,
            I => \N__26518\
        );

    \I__4936\ : InMux
    port map (
            O => \N__26544\,
            I => \N__26511\
        );

    \I__4935\ : InMux
    port map (
            O => \N__26543\,
            I => \N__26511\
        );

    \I__4934\ : InMux
    port map (
            O => \N__26540\,
            I => \N__26511\
        );

    \I__4933\ : CascadeMux
    port map (
            O => \N__26539\,
            I => \N__26508\
        );

    \I__4932\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26505\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__26535\,
            I => \N__26500\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__26530\,
            I => \N__26500\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__26523\,
            I => \N__26495\
        );

    \I__4928\ : Span4Mux_s2_v
    port map (
            O => \N__26518\,
            I => \N__26495\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__26511\,
            I => \N__26492\
        );

    \I__4926\ : InMux
    port map (
            O => \N__26508\,
            I => \N__26489\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__26505\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__26500\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__26495\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4922\ : Odrv12
    port map (
            O => \N__26492\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__26489\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__4920\ : CascadeMux
    port map (
            O => \N__26478\,
            I => \N__26473\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__26477\,
            I => \N__26467\
        );

    \I__4918\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26464\
        );

    \I__4917\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26461\
        );

    \I__4916\ : InMux
    port map (
            O => \N__26472\,
            I => \N__26458\
        );

    \I__4915\ : CascadeMux
    port map (
            O => \N__26471\,
            I => \N__26455\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__26470\,
            I => \N__26450\
        );

    \I__4913\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26445\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__26464\,
            I => \N__26442\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__26461\,
            I => \N__26437\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__26458\,
            I => \N__26437\
        );

    \I__4909\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26434\
        );

    \I__4908\ : InMux
    port map (
            O => \N__26454\,
            I => \N__26427\
        );

    \I__4907\ : InMux
    port map (
            O => \N__26453\,
            I => \N__26427\
        );

    \I__4906\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26427\
        );

    \I__4905\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26422\
        );

    \I__4904\ : InMux
    port map (
            O => \N__26448\,
            I => \N__26422\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26419\
        );

    \I__4902\ : Span4Mux_s2_h
    port map (
            O => \N__26442\,
            I => \N__26414\
        );

    \I__4901\ : Span4Mux_s2_v
    port map (
            O => \N__26437\,
            I => \N__26414\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__26434\,
            I => \N__26409\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__26427\,
            I => \N__26409\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__26422\,
            I => \N__26406\
        );

    \I__4897\ : Odrv4
    port map (
            O => \N__26419\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_11\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__26414\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_11\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__26409\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_11\
        );

    \I__4894\ : Odrv12
    port map (
            O => \N__26406\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_11\
        );

    \I__4893\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26388\
        );

    \I__4892\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26385\
        );

    \I__4891\ : InMux
    port map (
            O => \N__26395\,
            I => \N__26382\
        );

    \I__4890\ : InMux
    port map (
            O => \N__26394\,
            I => \N__26379\
        );

    \I__4889\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26372\
        );

    \I__4888\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26372\
        );

    \I__4887\ : InMux
    port map (
            O => \N__26391\,
            I => \N__26372\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__26388\,
            I => \N__26364\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__26385\,
            I => \N__26361\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__26382\,
            I => \N__26358\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__26379\,
            I => \N__26352\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__26372\,
            I => \N__26349\
        );

    \I__4881\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26344\
        );

    \I__4880\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26344\
        );

    \I__4879\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26339\
        );

    \I__4878\ : InMux
    port map (
            O => \N__26368\,
            I => \N__26339\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__26367\,
            I => \N__26334\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__26364\,
            I => \N__26327\
        );

    \I__4875\ : Span4Mux_h
    port map (
            O => \N__26361\,
            I => \N__26327\
        );

    \I__4874\ : Span4Mux_s1_v
    port map (
            O => \N__26358\,
            I => \N__26327\
        );

    \I__4873\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26324\
        );

    \I__4872\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26319\
        );

    \I__4871\ : InMux
    port map (
            O => \N__26355\,
            I => \N__26319\
        );

    \I__4870\ : Span4Mux_s1_v
    port map (
            O => \N__26352\,
            I => \N__26310\
        );

    \I__4869\ : Span4Mux_s1_v
    port map (
            O => \N__26349\,
            I => \N__26310\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__26344\,
            I => \N__26310\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26310\
        );

    \I__4866\ : InMux
    port map (
            O => \N__26338\,
            I => \N__26305\
        );

    \I__4865\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26305\
        );

    \I__4864\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26302\
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__26327\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__26324\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__26319\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__26310\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__26305\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__26302\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__4857\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26286\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__26286\,
            I => \POWERLED.un1_m2_2_0\
        );

    \I__4855\ : CascadeMux
    port map (
            O => \N__26283\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2_cascade_\
        );

    \I__4854\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26277\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__26277\,
            I => \VPP_VDDQ.count_2_rst_6\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__26274\,
            I => \VPP_VDDQ.count_2_rst_6_cascade_\
        );

    \I__4851\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26267\
        );

    \I__4850\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26264\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__26267\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__26264\,
            I => \VPP_VDDQ.un1_count_2_1_axb_2\
        );

    \I__4847\ : InMux
    port map (
            O => \N__26259\,
            I => \N__26253\
        );

    \I__4846\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26253\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__26253\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\
        );

    \I__4844\ : InMux
    port map (
            O => \N__26250\,
            I => \N__26244\
        );

    \I__4843\ : InMux
    port map (
            O => \N__26249\,
            I => \N__26244\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__26244\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__26241\,
            I => \VPP_VDDQ.count_2_rst_5_cascade_\
        );

    \I__4840\ : InMux
    port map (
            O => \N__26238\,
            I => \N__26231\
        );

    \I__4839\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26231\
        );

    \I__4838\ : InMux
    port map (
            O => \N__26236\,
            I => \N__26228\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__26231\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__26228\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__4835\ : InMux
    port map (
            O => \N__26223\,
            I => \N__26217\
        );

    \I__4834\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26217\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__26217\,
            I => \N__26214\
        );

    \I__4832\ : Odrv4
    port map (
            O => \N__26214\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__26211\,
            I => \VPP_VDDQ.count_2Z0Z_3_cascade_\
        );

    \I__4830\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26205\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__26205\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__4828\ : CascadeMux
    port map (
            O => \N__26202\,
            I => \POWERLED.dutycycle_RNIZ0Z_1_cascade_\
        );

    \I__4827\ : InMux
    port map (
            O => \N__26199\,
            I => \N__26196\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__26196\,
            I => \N__26193\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__26193\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_2\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__26190\,
            I => \N__26184\
        );

    \I__4823\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26179\
        );

    \I__4822\ : CascadeMux
    port map (
            O => \N__26188\,
            I => \N__26173\
        );

    \I__4821\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26165\
        );

    \I__4820\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26165\
        );

    \I__4819\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26165\
        );

    \I__4818\ : CascadeMux
    port map (
            O => \N__26182\,
            I => \N__26160\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__26179\,
            I => \N__26157\
        );

    \I__4816\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26154\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__26177\,
            I => \N__26150\
        );

    \I__4814\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26139\
        );

    \I__4813\ : InMux
    port map (
            O => \N__26173\,
            I => \N__26139\
        );

    \I__4812\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26139\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__26165\,
            I => \N__26136\
        );

    \I__4810\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26131\
        );

    \I__4809\ : InMux
    port map (
            O => \N__26163\,
            I => \N__26131\
        );

    \I__4808\ : InMux
    port map (
            O => \N__26160\,
            I => \N__26128\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__26157\,
            I => \N__26123\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__26154\,
            I => \N__26123\
        );

    \I__4805\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26116\
        );

    \I__4804\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26116\
        );

    \I__4803\ : InMux
    port map (
            O => \N__26149\,
            I => \N__26116\
        );

    \I__4802\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26109\
        );

    \I__4801\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26109\
        );

    \I__4800\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26109\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__26139\,
            I => \N__26100\
        );

    \I__4798\ : Sp12to4
    port map (
            O => \N__26136\,
            I => \N__26100\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26100\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__26128\,
            I => \N__26100\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__26123\,
            I => \N__26093\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__26116\,
            I => \N__26093\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__26109\,
            I => \N__26093\
        );

    \I__4792\ : Span12Mux_s3_v
    port map (
            O => \N__26100\,
            I => \N__26090\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__26093\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__4790\ : Odrv12
    port map (
            O => \N__26090\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__26085\,
            I => \N__26082\
        );

    \I__4788\ : InMux
    port map (
            O => \N__26082\,
            I => \N__26079\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__4786\ : Span4Mux_h
    port map (
            O => \N__26076\,
            I => \N__26073\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__26073\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_8\
        );

    \I__4784\ : CascadeMux
    port map (
            O => \N__26070\,
            I => \N__26067\
        );

    \I__4783\ : InMux
    port map (
            O => \N__26067\,
            I => \N__26064\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__26064\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_13\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__4780\ : InMux
    port map (
            O => \N__26058\,
            I => \N__26055\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__26055\,
            I => \N__26052\
        );

    \I__4778\ : Odrv12
    port map (
            O => \N__26052\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_7\
        );

    \I__4777\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26046\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__26046\,
            I => \N__26043\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__26043\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__4774\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26037\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__26037\,
            I => \N__26034\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__26034\,
            I => \POWERLED.un1_dutycycle_53_axb_11\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__26031\,
            I => \N__26028\
        );

    \I__4770\ : InMux
    port map (
            O => \N__26028\,
            I => \N__26025\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__26025\,
            I => \N__26022\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__26022\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_14\
        );

    \I__4767\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26016\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__26016\,
            I => \N__26013\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__26013\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_15\
        );

    \I__4764\ : InMux
    port map (
            O => \N__26010\,
            I => \N__26007\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__26007\,
            I => \N__26004\
        );

    \I__4762\ : Span4Mux_s1_v
    port map (
            O => \N__26004\,
            I => \N__25999\
        );

    \I__4761\ : InMux
    port map (
            O => \N__26003\,
            I => \N__25996\
        );

    \I__4760\ : InMux
    port map (
            O => \N__26002\,
            I => \N__25993\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__25999\,
            I => \POWERLED.un1_dutycycle_53_44_d_1_a0_0\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__25996\,
            I => \POWERLED.un1_dutycycle_53_44_d_1_a0_0\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__25993\,
            I => \POWERLED.un1_dutycycle_53_44_d_1_a0_0\
        );

    \I__4756\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25983\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25978\
        );

    \I__4754\ : CascadeMux
    port map (
            O => \N__25982\,
            I => \N__25974\
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__25981\,
            I => \N__25967\
        );

    \I__4752\ : Span4Mux_v
    port map (
            O => \N__25978\,
            I => \N__25964\
        );

    \I__4751\ : InMux
    port map (
            O => \N__25977\,
            I => \N__25961\
        );

    \I__4750\ : InMux
    port map (
            O => \N__25974\,
            I => \N__25956\
        );

    \I__4749\ : InMux
    port map (
            O => \N__25973\,
            I => \N__25956\
        );

    \I__4748\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25951\
        );

    \I__4747\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25951\
        );

    \I__4746\ : InMux
    port map (
            O => \N__25970\,
            I => \N__25948\
        );

    \I__4745\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25945\
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__25964\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__25961\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__25956\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__25951\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__25948\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__25945\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__25932\,
            I => \N__25926\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__25931\,
            I => \N__25922\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__25930\,
            I => \N__25919\
        );

    \I__4735\ : InMux
    port map (
            O => \N__25929\,
            I => \N__25913\
        );

    \I__4734\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25910\
        );

    \I__4733\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25907\
        );

    \I__4732\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25904\
        );

    \I__4731\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25899\
        );

    \I__4730\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25899\
        );

    \I__4729\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25894\
        );

    \I__4728\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25894\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__25913\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__25910\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__25907\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__25904\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__25899\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__25894\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4721\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25878\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__25878\,
            I => \N__25875\
        );

    \I__4719\ : Span4Mux_s3_h
    port map (
            O => \N__25875\,
            I => \N__25871\
        );

    \I__4718\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25868\
        );

    \I__4717\ : Odrv4
    port map (
            O => \N__25871\,
            I => \POWERLED.N_361\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__25868\,
            I => \POWERLED.N_361\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__25863\,
            I => \N__25857\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__25862\,
            I => \N__25853\
        );

    \I__4713\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25849\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__25860\,
            I => \N__25845\
        );

    \I__4711\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25841\
        );

    \I__4710\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25838\
        );

    \I__4709\ : InMux
    port map (
            O => \N__25853\,
            I => \N__25833\
        );

    \I__4708\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25833\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__25849\,
            I => \N__25830\
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__25848\,
            I => \N__25825\
        );

    \I__4705\ : InMux
    port map (
            O => \N__25845\,
            I => \N__25822\
        );

    \I__4704\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25819\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25816\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__25838\,
            I => \N__25811\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__25833\,
            I => \N__25811\
        );

    \I__4700\ : Span4Mux_h
    port map (
            O => \N__25830\,
            I => \N__25808\
        );

    \I__4699\ : InMux
    port map (
            O => \N__25829\,
            I => \N__25803\
        );

    \I__4698\ : InMux
    port map (
            O => \N__25828\,
            I => \N__25803\
        );

    \I__4697\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25800\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__25822\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__25819\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__25816\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__25811\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4692\ : Odrv4
    port map (
            O => \N__25808\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__25803\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__25800\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9\
        );

    \I__4689\ : CascadeMux
    port map (
            O => \N__25785\,
            I => \POWERLED.un2_count_clk_17_0_a2_1_4_cascade_\
        );

    \I__4688\ : CascadeMux
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__4687\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25773\
        );

    \I__4686\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25773\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__25773\,
            I => \N__25770\
        );

    \I__4684\ : Span4Mux_s2_h
    port map (
            O => \N__25770\,
            I => \N__25767\
        );

    \I__4683\ : Span4Mux_h
    port map (
            O => \N__25767\,
            I => \N__25764\
        );

    \I__4682\ : Odrv4
    port map (
            O => \N__25764\,
            I => \POWERLED.N_369\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__25761\,
            I => \N__25755\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__25760\,
            I => \N__25748\
        );

    \I__4679\ : InMux
    port map (
            O => \N__25759\,
            I => \N__25736\
        );

    \I__4678\ : InMux
    port map (
            O => \N__25758\,
            I => \N__25736\
        );

    \I__4677\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25736\
        );

    \I__4676\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25736\
        );

    \I__4675\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25736\
        );

    \I__4674\ : InMux
    port map (
            O => \N__25752\,
            I => \N__25733\
        );

    \I__4673\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25730\
        );

    \I__4672\ : InMux
    port map (
            O => \N__25748\,
            I => \N__25725\
        );

    \I__4671\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25725\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__25736\,
            I => \N__25722\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__25733\,
            I => \N__25719\
        );

    \I__4668\ : InMux
    port map (
            O => \N__25730\,
            I => \N__25716\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__25725\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4666\ : Odrv4
    port map (
            O => \N__25722\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4665\ : Odrv4
    port map (
            O => \N__25719\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__25716\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__25707\,
            I => \N__25703\
        );

    \I__4662\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25698\
        );

    \I__4661\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25698\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__25698\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_8\
        );

    \I__4659\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25692\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__25692\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__4657\ : InMux
    port map (
            O => \N__25689\,
            I => \POWERLED.un1_dutycycle_53_cry_9\
        );

    \I__4656\ : InMux
    port map (
            O => \N__25686\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__25683\,
            I => \N__25680\
        );

    \I__4654\ : InMux
    port map (
            O => \N__25680\,
            I => \N__25677\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__25677\,
            I => \POWERLED.dutycycle_RNIZ0Z_15\
        );

    \I__4652\ : InMux
    port map (
            O => \N__25674\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__4651\ : InMux
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__25665\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_13\
        );

    \I__4648\ : InMux
    port map (
            O => \N__25662\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__4647\ : InMux
    port map (
            O => \N__25659\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__4646\ : InMux
    port map (
            O => \N__25656\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__4645\ : InMux
    port map (
            O => \N__25653\,
            I => \bfn_7_15_0_\
        );

    \I__4644\ : InMux
    port map (
            O => \N__25650\,
            I => \POWERLED.CO2\
        );

    \I__4643\ : InMux
    port map (
            O => \N__25647\,
            I => \N__25642\
        );

    \I__4642\ : InMux
    port map (
            O => \N__25646\,
            I => \N__25637\
        );

    \I__4641\ : InMux
    port map (
            O => \N__25645\,
            I => \N__25637\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__25642\,
            I => \N__25634\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__25637\,
            I => \N__25629\
        );

    \I__4638\ : Span12Mux_s10_h
    port map (
            O => \N__25634\,
            I => \N__25626\
        );

    \I__4637\ : InMux
    port map (
            O => \N__25633\,
            I => \N__25621\
        );

    \I__4636\ : InMux
    port map (
            O => \N__25632\,
            I => \N__25621\
        );

    \I__4635\ : Odrv4
    port map (
            O => \N__25629\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_5\
        );

    \I__4634\ : Odrv12
    port map (
            O => \N__25626\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_5\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__25621\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_5\
        );

    \I__4632\ : InMux
    port map (
            O => \N__25614\,
            I => \POWERLED.un1_dutycycle_53_cry_1_cZ0\
        );

    \I__4631\ : InMux
    port map (
            O => \N__25611\,
            I => \POWERLED.un1_dutycycle_53_cry_2_cZ0\
        );

    \I__4630\ : InMux
    port map (
            O => \N__25608\,
            I => \POWERLED.un1_dutycycle_53_cry_3_cZ0\
        );

    \I__4629\ : InMux
    port map (
            O => \N__25605\,
            I => \N__25602\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__25602\,
            I => \N__25599\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__25596\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_5\
        );

    \I__4625\ : InMux
    port map (
            O => \N__25593\,
            I => \POWERLED.un1_dutycycle_53_cry_4\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__4623\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25584\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__4621\ : Odrv12
    port map (
            O => \N__25581\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5\
        );

    \I__4620\ : InMux
    port map (
            O => \N__25578\,
            I => \POWERLED.un1_dutycycle_53_cry_5\
        );

    \I__4619\ : CascadeMux
    port map (
            O => \N__25575\,
            I => \N__25572\
        );

    \I__4618\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25566\
        );

    \I__4616\ : Span4Mux_h
    port map (
            O => \N__25566\,
            I => \N__25563\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__25563\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_10\
        );

    \I__4614\ : InMux
    port map (
            O => \N__25560\,
            I => \POWERLED.un1_dutycycle_53_cry_6\
        );

    \I__4613\ : InMux
    port map (
            O => \N__25557\,
            I => \N__25551\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__25556\,
            I => \N__25548\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__25555\,
            I => \N__25545\
        );

    \I__4610\ : InMux
    port map (
            O => \N__25554\,
            I => \N__25540\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__25551\,
            I => \N__25537\
        );

    \I__4608\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25534\
        );

    \I__4607\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25529\
        );

    \I__4606\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25529\
        );

    \I__4605\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25524\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__25540\,
            I => \N__25521\
        );

    \I__4603\ : Span4Mux_h
    port map (
            O => \N__25537\,
            I => \N__25516\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__25534\,
            I => \N__25516\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__25529\,
            I => \N__25513\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__25528\,
            I => \N__25510\
        );

    \I__4599\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25507\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__25524\,
            I => \N__25502\
        );

    \I__4597\ : Span4Mux_s2_v
    port map (
            O => \N__25521\,
            I => \N__25502\
        );

    \I__4596\ : Span4Mux_s1_v
    port map (
            O => \N__25516\,
            I => \N__25497\
        );

    \I__4595\ : Span4Mux_h
    port map (
            O => \N__25513\,
            I => \N__25497\
        );

    \I__4594\ : InMux
    port map (
            O => \N__25510\,
            I => \N__25494\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__25507\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__25502\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__25497\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__25494\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__25485\,
            I => \N__25482\
        );

    \I__4588\ : InMux
    port map (
            O => \N__25482\,
            I => \N__25479\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__4586\ : Span4Mux_h
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__4585\ : Span4Mux_h
    port map (
            O => \N__25473\,
            I => \N__25470\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__25470\,
            I => \POWERLED.dutycycle_RNIZ0Z_11\
        );

    \I__4583\ : InMux
    port map (
            O => \N__25467\,
            I => \bfn_7_14_0_\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__25464\,
            I => \N__25461\
        );

    \I__4581\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__4579\ : Span4Mux_h
    port map (
            O => \N__25455\,
            I => \N__25452\
        );

    \I__4578\ : Span4Mux_h
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__25449\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_12\
        );

    \I__4576\ : InMux
    port map (
            O => \N__25446\,
            I => \POWERLED.un1_dutycycle_53_cry_8\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__25443\,
            I => \N__25438\
        );

    \I__4574\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25432\
        );

    \I__4573\ : InMux
    port map (
            O => \N__25441\,
            I => \N__25432\
        );

    \I__4572\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25427\
        );

    \I__4571\ : InMux
    port map (
            O => \N__25437\,
            I => \N__25427\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__25432\,
            I => \N__25422\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__25427\,
            I => \N__25419\
        );

    \I__4568\ : InMux
    port map (
            O => \N__25426\,
            I => \N__25416\
        );

    \I__4567\ : InMux
    port map (
            O => \N__25425\,
            I => \N__25413\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__25422\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__25419\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__25416\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__25413\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__25404\,
            I => \N__25401\
        );

    \I__4561\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25381\
        );

    \I__4560\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25381\
        );

    \I__4559\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25372\
        );

    \I__4558\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25372\
        );

    \I__4557\ : InMux
    port map (
            O => \N__25397\,
            I => \N__25372\
        );

    \I__4556\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25363\
        );

    \I__4555\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25363\
        );

    \I__4554\ : InMux
    port map (
            O => \N__25394\,
            I => \N__25363\
        );

    \I__4553\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25363\
        );

    \I__4552\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25356\
        );

    \I__4551\ : InMux
    port map (
            O => \N__25391\,
            I => \N__25356\
        );

    \I__4550\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25356\
        );

    \I__4549\ : InMux
    port map (
            O => \N__25389\,
            I => \N__25347\
        );

    \I__4548\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25347\
        );

    \I__4547\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25347\
        );

    \I__4546\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25347\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__25381\,
            I => \N__25344\
        );

    \I__4544\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25339\
        );

    \I__4543\ : InMux
    port map (
            O => \N__25379\,
            I => \N__25339\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__25372\,
            I => \N__25330\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__25363\,
            I => \N__25330\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__25356\,
            I => \N__25330\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25330\
        );

    \I__4538\ : Span4Mux_v
    port map (
            O => \N__25344\,
            I => \N__25327\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__25339\,
            I => \POWERLED.func_state_RNI43L44_0_0\
        );

    \I__4536\ : Odrv12
    port map (
            O => \N__25330\,
            I => \POWERLED.func_state_RNI43L44_0_0\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__25327\,
            I => \POWERLED.func_state_RNI43L44_0_0\
        );

    \I__4534\ : InMux
    port map (
            O => \N__25320\,
            I => \N__25317\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__25317\,
            I => \N__25314\
        );

    \I__4532\ : Odrv4
    port map (
            O => \N__25314\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__4531\ : CascadeMux
    port map (
            O => \N__25311\,
            I => \N__25305\
        );

    \I__4530\ : CEMux
    port map (
            O => \N__25310\,
            I => \N__25299\
        );

    \I__4529\ : CEMux
    port map (
            O => \N__25309\,
            I => \N__25296\
        );

    \I__4528\ : InMux
    port map (
            O => \N__25308\,
            I => \N__25286\
        );

    \I__4527\ : InMux
    port map (
            O => \N__25305\,
            I => \N__25286\
        );

    \I__4526\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25286\
        );

    \I__4525\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25286\
        );

    \I__4524\ : CEMux
    port map (
            O => \N__25302\,
            I => \N__25280\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__25299\,
            I => \N__25274\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__25296\,
            I => \N__25274\
        );

    \I__4521\ : CEMux
    port map (
            O => \N__25295\,
            I => \N__25271\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25268\
        );

    \I__4519\ : CEMux
    port map (
            O => \N__25285\,
            I => \N__25261\
        );

    \I__4518\ : InMux
    port map (
            O => \N__25284\,
            I => \N__25261\
        );

    \I__4517\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25261\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__25280\,
            I => \N__25258\
        );

    \I__4515\ : CascadeMux
    port map (
            O => \N__25279\,
            I => \N__25255\
        );

    \I__4514\ : Span4Mux_v
    port map (
            O => \N__25274\,
            I => \N__25247\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25247\
        );

    \I__4512\ : Span4Mux_v
    port map (
            O => \N__25268\,
            I => \N__25239\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__25261\,
            I => \N__25239\
        );

    \I__4510\ : Span4Mux_h
    port map (
            O => \N__25258\,
            I => \N__25231\
        );

    \I__4509\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25224\
        );

    \I__4508\ : InMux
    port map (
            O => \N__25254\,
            I => \N__25224\
        );

    \I__4507\ : InMux
    port map (
            O => \N__25253\,
            I => \N__25224\
        );

    \I__4506\ : CEMux
    port map (
            O => \N__25252\,
            I => \N__25221\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__25247\,
            I => \N__25218\
        );

    \I__4504\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25211\
        );

    \I__4503\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25211\
        );

    \I__4502\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25211\
        );

    \I__4501\ : Span4Mux_h
    port map (
            O => \N__25239\,
            I => \N__25208\
        );

    \I__4500\ : CEMux
    port map (
            O => \N__25238\,
            I => \N__25197\
        );

    \I__4499\ : InMux
    port map (
            O => \N__25237\,
            I => \N__25197\
        );

    \I__4498\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25197\
        );

    \I__4497\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25197\
        );

    \I__4496\ : InMux
    port map (
            O => \N__25234\,
            I => \N__25197\
        );

    \I__4495\ : Span4Mux_s3_h
    port map (
            O => \N__25231\,
            I => \N__25192\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__25224\,
            I => \N__25192\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__25221\,
            I => \POWERLED.count_clk_en\
        );

    \I__4492\ : Odrv4
    port map (
            O => \N__25218\,
            I => \POWERLED.count_clk_en\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__25211\,
            I => \POWERLED.count_clk_en\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__25208\,
            I => \POWERLED.count_clk_en\
        );

    \I__4489\ : LocalMux
    port map (
            O => \N__25197\,
            I => \POWERLED.count_clk_en\
        );

    \I__4488\ : Odrv4
    port map (
            O => \N__25192\,
            I => \POWERLED.count_clk_en\
        );

    \I__4487\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25172\
        );

    \I__4486\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25167\
        );

    \I__4485\ : InMux
    port map (
            O => \N__25177\,
            I => \N__25167\
        );

    \I__4484\ : InMux
    port map (
            O => \N__25176\,
            I => \N__25164\
        );

    \I__4483\ : CascadeMux
    port map (
            O => \N__25175\,
            I => \N__25161\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__25172\,
            I => \N__25155\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__25167\,
            I => \N__25155\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__25164\,
            I => \N__25152\
        );

    \I__4479\ : InMux
    port map (
            O => \N__25161\,
            I => \N__25149\
        );

    \I__4478\ : InMux
    port map (
            O => \N__25160\,
            I => \N__25146\
        );

    \I__4477\ : Span4Mux_s2_v
    port map (
            O => \N__25155\,
            I => \N__25139\
        );

    \I__4476\ : Span4Mux_s1_h
    port map (
            O => \N__25152\,
            I => \N__25139\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__25149\,
            I => \N__25139\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__25146\,
            I => \N__25135\
        );

    \I__4473\ : Span4Mux_h
    port map (
            O => \N__25139\,
            I => \N__25132\
        );

    \I__4472\ : InMux
    port map (
            O => \N__25138\,
            I => \N__25129\
        );

    \I__4471\ : Odrv12
    port map (
            O => \N__25135\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__4470\ : Odrv4
    port map (
            O => \N__25132\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__25129\,
            I => \POWERLED.count_clk_RNIZ0Z_6\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__25122\,
            I => \N__25115\
        );

    \I__4467\ : CascadeMux
    port map (
            O => \N__25121\,
            I => \N__25110\
        );

    \I__4466\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25102\
        );

    \I__4465\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25099\
        );

    \I__4464\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25096\
        );

    \I__4463\ : InMux
    port map (
            O => \N__25115\,
            I => \N__25089\
        );

    \I__4462\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25089\
        );

    \I__4461\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25089\
        );

    \I__4460\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25086\
        );

    \I__4459\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25081\
        );

    \I__4458\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25081\
        );

    \I__4457\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25078\
        );

    \I__4456\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25075\
        );

    \I__4455\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25071\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__25102\,
            I => \N__25068\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25065\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__25096\,
            I => \N__25062\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25055\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__25086\,
            I => \N__25055\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__25081\,
            I => \N__25055\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__25078\,
            I => \N__25050\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__25075\,
            I => \N__25050\
        );

    \I__4446\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25047\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__25071\,
            I => \N__25044\
        );

    \I__4444\ : Span4Mux_s2_h
    port map (
            O => \N__25068\,
            I => \N__25037\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__25065\,
            I => \N__25037\
        );

    \I__4442\ : Span4Mux_v
    port map (
            O => \N__25062\,
            I => \N__25037\
        );

    \I__4441\ : Span4Mux_v
    port map (
            O => \N__25055\,
            I => \N__25030\
        );

    \I__4440\ : Span4Mux_v
    port map (
            O => \N__25050\,
            I => \N__25030\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__25047\,
            I => \N__25030\
        );

    \I__4438\ : Odrv4
    port map (
            O => \N__25044\,
            I => \POWERLED.N_175\
        );

    \I__4437\ : Odrv4
    port map (
            O => \N__25037\,
            I => \POWERLED.N_175\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__25030\,
            I => \POWERLED.N_175\
        );

    \I__4435\ : InMux
    port map (
            O => \N__25023\,
            I => \N__25008\
        );

    \I__4434\ : InMux
    port map (
            O => \N__25022\,
            I => \N__25008\
        );

    \I__4433\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25008\
        );

    \I__4432\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25008\
        );

    \I__4431\ : CascadeMux
    port map (
            O => \N__25019\,
            I => \N__25000\
        );

    \I__4430\ : CascadeMux
    port map (
            O => \N__25018\,
            I => \N__24995\
        );

    \I__4429\ : InMux
    port map (
            O => \N__25017\,
            I => \N__24992\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__25008\,
            I => \N__24989\
        );

    \I__4427\ : InMux
    port map (
            O => \N__25007\,
            I => \N__24982\
        );

    \I__4426\ : InMux
    port map (
            O => \N__25006\,
            I => \N__24982\
        );

    \I__4425\ : InMux
    port map (
            O => \N__25005\,
            I => \N__24982\
        );

    \I__4424\ : InMux
    port map (
            O => \N__25004\,
            I => \N__24969\
        );

    \I__4423\ : InMux
    port map (
            O => \N__25003\,
            I => \N__24969\
        );

    \I__4422\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24969\
        );

    \I__4421\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24969\
        );

    \I__4420\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24969\
        );

    \I__4419\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24969\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__24992\,
            I => \N__24966\
        );

    \I__4417\ : Span4Mux_v
    port map (
            O => \N__24989\,
            I => \N__24963\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__24982\,
            I => \N__24958\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__24969\,
            I => \N__24958\
        );

    \I__4414\ : Span4Mux_v
    port map (
            O => \N__24966\,
            I => \N__24951\
        );

    \I__4413\ : Span4Mux_h
    port map (
            O => \N__24963\,
            I => \N__24951\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__24958\,
            I => \N__24951\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__24951\,
            I => \POWERLED.N_175_i\
        );

    \I__4410\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24942\
        );

    \I__4409\ : InMux
    port map (
            O => \N__24947\,
            I => \N__24937\
        );

    \I__4408\ : InMux
    port map (
            O => \N__24946\,
            I => \N__24937\
        );

    \I__4407\ : InMux
    port map (
            O => \N__24945\,
            I => \N__24932\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__24942\,
            I => \N__24927\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__24937\,
            I => \N__24927\
        );

    \I__4404\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24924\
        );

    \I__4403\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24921\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__24932\,
            I => \N__24918\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__24927\,
            I => \N__24915\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__24924\,
            I => \N__24912\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__24921\,
            I => \N__24909\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__24918\,
            I => \N__24906\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__24915\,
            I => \N__24901\
        );

    \I__4396\ : Span4Mux_h
    port map (
            O => \N__24912\,
            I => \N__24901\
        );

    \I__4395\ : Span4Mux_s2_v
    port map (
            O => \N__24909\,
            I => \N__24896\
        );

    \I__4394\ : Span4Mux_v
    port map (
            O => \N__24906\,
            I => \N__24896\
        );

    \I__4393\ : Span4Mux_h
    port map (
            O => \N__24901\,
            I => \N__24893\
        );

    \I__4392\ : Odrv4
    port map (
            O => \N__24896\,
            I => \POWERLED.N_428\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__24893\,
            I => \POWERLED.N_428\
        );

    \I__4390\ : InMux
    port map (
            O => \N__24888\,
            I => \N__24882\
        );

    \I__4389\ : InMux
    port map (
            O => \N__24887\,
            I => \N__24882\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__24882\,
            I => \N__24879\
        );

    \I__4387\ : Span4Mux_s3_h
    port map (
            O => \N__24879\,
            I => \N__24873\
        );

    \I__4386\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24866\
        );

    \I__4385\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24866\
        );

    \I__4384\ : InMux
    port map (
            O => \N__24876\,
            I => \N__24866\
        );

    \I__4383\ : Span4Mux_h
    port map (
            O => \N__24873\,
            I => \N__24863\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__24866\,
            I => \N__24860\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__24863\,
            I => \POWERLED.func_state_RNI_5Z0Z_0\
        );

    \I__4380\ : Odrv4
    port map (
            O => \N__24860\,
            I => \POWERLED.func_state_RNI_5Z0Z_0\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__4378\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__24849\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_0\
        );

    \I__4376\ : InMux
    port map (
            O => \N__24846\,
            I => \POWERLED.un1_dutycycle_53_cry_0_cZ0\
        );

    \I__4375\ : InMux
    port map (
            O => \N__24843\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__4374\ : InMux
    port map (
            O => \N__24840\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__4373\ : InMux
    port map (
            O => \N__24837\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__4372\ : InMux
    port map (
            O => \N__24834\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__4371\ : InMux
    port map (
            O => \N__24831\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__4370\ : InMux
    port map (
            O => \N__24828\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__24825\,
            I => \N__24822\
        );

    \I__4368\ : InMux
    port map (
            O => \N__24822\,
            I => \N__24813\
        );

    \I__4367\ : InMux
    port map (
            O => \N__24821\,
            I => \N__24813\
        );

    \I__4366\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24813\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__24813\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__4364\ : InMux
    port map (
            O => \N__24810\,
            I => \N__24805\
        );

    \I__4363\ : InMux
    port map (
            O => \N__24809\,
            I => \N__24802\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__24808\,
            I => \N__24797\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__24805\,
            I => \N__24794\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__24802\,
            I => \N__24791\
        );

    \I__4359\ : InMux
    port map (
            O => \N__24801\,
            I => \N__24786\
        );

    \I__4358\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24786\
        );

    \I__4357\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24783\
        );

    \I__4356\ : Odrv12
    port map (
            O => \N__24794\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__24791\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__24786\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__24783\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__4352\ : InMux
    port map (
            O => \N__24774\,
            I => \N__24771\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__24771\,
            I => \N__24768\
        );

    \I__4350\ : Odrv12
    port map (
            O => \N__24768\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__4349\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24762\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__24762\,
            I => \N__24759\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__24759\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__24756\,
            I => \N__24752\
        );

    \I__4345\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24749\
        );

    \I__4344\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24746\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__24749\,
            I => \N__24741\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24741\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__24741\,
            I => \N__24737\
        );

    \I__4340\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24734\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__24737\,
            I => \POWERLED.N_193\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__24734\,
            I => \POWERLED.N_193\
        );

    \I__4337\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24725\
        );

    \I__4336\ : InMux
    port map (
            O => \N__24728\,
            I => \N__24722\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__24725\,
            I => \N__24717\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__24722\,
            I => \N__24717\
        );

    \I__4333\ : Odrv4
    port map (
            O => \N__24717\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__4332\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24708\
        );

    \I__4331\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24708\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__24708\,
            I => \POWERLED.N_178\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__24705\,
            I => \POWERLED.count_clkZ0Z_9_cascade_\
        );

    \I__4328\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24695\
        );

    \I__4327\ : InMux
    port map (
            O => \N__24701\,
            I => \N__24695\
        );

    \I__4326\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24692\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__24695\,
            I => \POWERLED.N_385\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__24692\,
            I => \POWERLED.N_385\
        );

    \I__4323\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24681\
        );

    \I__4322\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24678\
        );

    \I__4321\ : InMux
    port map (
            O => \N__24685\,
            I => \N__24673\
        );

    \I__4320\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24673\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__24681\,
            I => \N__24668\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__24678\,
            I => \N__24668\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24664\
        );

    \I__4316\ : Span4Mux_v
    port map (
            O => \N__24668\,
            I => \N__24661\
        );

    \I__4315\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24658\
        );

    \I__4314\ : Odrv4
    port map (
            O => \N__24664\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__24661\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__24658\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__24651\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__24648\,
            I => \N__24643\
        );

    \I__4309\ : InMux
    port map (
            O => \N__24647\,
            I => \N__24640\
        );

    \I__4308\ : InMux
    port map (
            O => \N__24646\,
            I => \N__24635\
        );

    \I__4307\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24635\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__24640\,
            I => \N__24632\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__24635\,
            I => \N__24629\
        );

    \I__4304\ : Span4Mux_v
    port map (
            O => \N__24632\,
            I => \N__24626\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__24629\,
            I => \N__24623\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__24626\,
            I => \POWERLED.count_clk_RNI_0Z0Z_1\
        );

    \I__4301\ : Odrv4
    port map (
            O => \N__24623\,
            I => \POWERLED.count_clk_RNI_0Z0Z_1\
        );

    \I__4300\ : InMux
    port map (
            O => \N__24618\,
            I => \N__24615\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__24615\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__4298\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24606\
        );

    \I__4297\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24606\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__24606\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__4295\ : CascadeMux
    port map (
            O => \N__24603\,
            I => \N__24599\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__24602\,
            I => \N__24595\
        );

    \I__4293\ : InMux
    port map (
            O => \N__24599\,
            I => \N__24590\
        );

    \I__4292\ : InMux
    port map (
            O => \N__24598\,
            I => \N__24590\
        );

    \I__4291\ : InMux
    port map (
            O => \N__24595\,
            I => \N__24587\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__24590\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__24587\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__4288\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24576\
        );

    \I__4287\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24576\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__24576\,
            I => \POWERLED.count_clk_1_9\
        );

    \I__4285\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24570\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__24570\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__4283\ : CascadeMux
    port map (
            O => \N__24567\,
            I => \N__24564\
        );

    \I__4282\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24561\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__24561\,
            I => \N__24558\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__24555\,
            I => \POWERLED.count_clk_RNIZ0Z_0\
        );

    \I__4278\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24545\
        );

    \I__4277\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24545\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__24550\,
            I => \N__24542\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__24545\,
            I => \N__24539\
        );

    \I__4274\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24536\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__24539\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__24536\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__24531\,
            I => \N__24527\
        );

    \I__4270\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24522\
        );

    \I__4269\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24522\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__24522\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__4267\ : InMux
    port map (
            O => \N__24519\,
            I => \N__24516\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__24516\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__4265\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24510\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__24510\,
            I => \N__24507\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__24507\,
            I => \N__24504\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__24504\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__4261\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__24492\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_4\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__24489\,
            I => \POWERLED.count_clkZ0Z_15_cascade_\
        );

    \I__4256\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24483\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__24483\,
            I => \POWERLED.count_clk_0_14\
        );

    \I__4254\ : InMux
    port map (
            O => \N__24480\,
            I => \N__24474\
        );

    \I__4253\ : InMux
    port map (
            O => \N__24479\,
            I => \N__24474\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__24474\,
            I => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\
        );

    \I__4251\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24467\
        );

    \I__4250\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24464\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__24467\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__24464\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__4247\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24455\
        );

    \I__4246\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24452\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__24455\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__24452\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__4243\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24444\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__24444\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__4241\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24438\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__24438\,
            I => \POWERLED.count_0_11\
        );

    \I__4239\ : InMux
    port map (
            O => \N__24435\,
            I => \N__24432\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__24432\,
            I => \POWERLED.count_0_3\
        );

    \I__4237\ : InMux
    port map (
            O => \N__24429\,
            I => \N__24426\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__24426\,
            I => \POWERLED.count_0_12\
        );

    \I__4235\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__24420\,
            I => \POWERLED.count_0_13\
        );

    \I__4233\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24413\
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__24416\,
            I => \N__24410\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__24413\,
            I => \N__24406\
        );

    \I__4230\ : InMux
    port map (
            O => \N__24410\,
            I => \N__24403\
        );

    \I__4229\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24400\
        );

    \I__4228\ : Span4Mux_v
    port map (
            O => \N__24406\,
            I => \N__24397\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__24403\,
            I => \PCH_PWRGD.N_424\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__24400\,
            I => \PCH_PWRGD.N_424\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__24397\,
            I => \PCH_PWRGD.N_424\
        );

    \I__4224\ : SRMux
    port map (
            O => \N__24390\,
            I => \N__24383\
        );

    \I__4223\ : SRMux
    port map (
            O => \N__24389\,
            I => \N__24380\
        );

    \I__4222\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24373\
        );

    \I__4221\ : SRMux
    port map (
            O => \N__24387\,
            I => \N__24373\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__24386\,
            I => \N__24365\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__24383\,
            I => \N__24354\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__24380\,
            I => \N__24350\
        );

    \I__4217\ : SRMux
    port map (
            O => \N__24379\,
            I => \N__24347\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__24378\,
            I => \N__24341\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__24373\,
            I => \N__24332\
        );

    \I__4214\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24329\
        );

    \I__4213\ : SRMux
    port map (
            O => \N__24371\,
            I => \N__24326\
        );

    \I__4212\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24321\
        );

    \I__4211\ : InMux
    port map (
            O => \N__24369\,
            I => \N__24321\
        );

    \I__4210\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24318\
        );

    \I__4209\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24309\
        );

    \I__4208\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24309\
        );

    \I__4207\ : InMux
    port map (
            O => \N__24363\,
            I => \N__24309\
        );

    \I__4206\ : InMux
    port map (
            O => \N__24362\,
            I => \N__24309\
        );

    \I__4205\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24306\
        );

    \I__4204\ : InMux
    port map (
            O => \N__24360\,
            I => \N__24297\
        );

    \I__4203\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24297\
        );

    \I__4202\ : InMux
    port map (
            O => \N__24358\,
            I => \N__24297\
        );

    \I__4201\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24297\
        );

    \I__4200\ : Span4Mux_s3_h
    port map (
            O => \N__24354\,
            I => \N__24292\
        );

    \I__4199\ : SRMux
    port map (
            O => \N__24353\,
            I => \N__24289\
        );

    \I__4198\ : Span4Mux_s3_v
    port map (
            O => \N__24350\,
            I => \N__24286\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24283\
        );

    \I__4196\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24280\
        );

    \I__4195\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24273\
        );

    \I__4194\ : InMux
    port map (
            O => \N__24344\,
            I => \N__24273\
        );

    \I__4193\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24273\
        );

    \I__4192\ : InMux
    port map (
            O => \N__24340\,
            I => \N__24264\
        );

    \I__4191\ : InMux
    port map (
            O => \N__24339\,
            I => \N__24264\
        );

    \I__4190\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24264\
        );

    \I__4189\ : InMux
    port map (
            O => \N__24337\,
            I => \N__24264\
        );

    \I__4188\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24259\
        );

    \I__4187\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24259\
        );

    \I__4186\ : Span4Mux_s2_v
    port map (
            O => \N__24332\,
            I => \N__24254\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__24329\,
            I => \N__24254\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__24326\,
            I => \N__24249\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__24321\,
            I => \N__24249\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__24318\,
            I => \N__24242\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__24309\,
            I => \N__24242\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__24306\,
            I => \N__24242\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__24297\,
            I => \N__24239\
        );

    \I__4178\ : SRMux
    port map (
            O => \N__24296\,
            I => \N__24234\
        );

    \I__4177\ : InMux
    port map (
            O => \N__24295\,
            I => \N__24234\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__24292\,
            I => \N__24229\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__24289\,
            I => \N__24229\
        );

    \I__4174\ : Sp12to4
    port map (
            O => \N__24286\,
            I => \N__24226\
        );

    \I__4173\ : Sp12to4
    port map (
            O => \N__24283\,
            I => \N__24215\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__24280\,
            I => \N__24215\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24215\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__24264\,
            I => \N__24215\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24215\
        );

    \I__4168\ : Span4Mux_v
    port map (
            O => \N__24254\,
            I => \N__24204\
        );

    \I__4167\ : Span4Mux_s2_h
    port map (
            O => \N__24249\,
            I => \N__24204\
        );

    \I__4166\ : Span4Mux_s2_v
    port map (
            O => \N__24242\,
            I => \N__24204\
        );

    \I__4165\ : Span4Mux_v
    port map (
            O => \N__24239\,
            I => \N__24204\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__24234\,
            I => \N__24204\
        );

    \I__4163\ : Sp12to4
    port map (
            O => \N__24229\,
            I => \N__24197\
        );

    \I__4162\ : Span12Mux_s10_v
    port map (
            O => \N__24226\,
            I => \N__24197\
        );

    \I__4161\ : Span12Mux_s5_v
    port map (
            O => \N__24215\,
            I => \N__24197\
        );

    \I__4160\ : Span4Mux_h
    port map (
            O => \N__24204\,
            I => \N__24194\
        );

    \I__4159\ : Odrv12
    port map (
            O => \N__24197\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4158\ : Odrv4
    port map (
            O => \N__24194\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4157\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24186\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__24186\,
            I => \POWERLED.count_0_5\
        );

    \I__4155\ : InMux
    port map (
            O => \N__24183\,
            I => \N__24180\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__24180\,
            I => \POWERLED.count_0_14\
        );

    \I__4153\ : InMux
    port map (
            O => \N__24177\,
            I => \N__24174\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__24174\,
            I => \N__24171\
        );

    \I__4151\ : Odrv4
    port map (
            O => \N__24171\,
            I => \POWERLED.count_0_6\
        );

    \I__4150\ : InMux
    port map (
            O => \N__24168\,
            I => \N__24165\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__24165\,
            I => \POWERLED.count_0_15\
        );

    \I__4148\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24159\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__24159\,
            I => \POWERLED.count_0_7\
        );

    \I__4146\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24153\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__24153\,
            I => \POWERLED.count_0_8\
        );

    \I__4144\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24147\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__24147\,
            I => \POWERLED.count_0_9\
        );

    \I__4142\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24141\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__24141\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__4140\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24132\
        );

    \I__4139\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24132\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__24132\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\
        );

    \I__4137\ : InMux
    port map (
            O => \N__24129\,
            I => \bfn_7_3_0_\
        );

    \I__4136\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24123\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__24123\,
            I => \N__24120\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__24120\,
            I => \VPP_VDDQ.un1_count_2_1_axb_10\
        );

    \I__4133\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24112\
        );

    \I__4132\ : InMux
    port map (
            O => \N__24116\,
            I => \N__24109\
        );

    \I__4131\ : InMux
    port map (
            O => \N__24115\,
            I => \N__24106\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__24112\,
            I => \N__24101\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__24109\,
            I => \N__24101\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__24106\,
            I => \N__24098\
        );

    \I__4127\ : Span4Mux_s2_v
    port map (
            O => \N__24101\,
            I => \N__24095\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__24098\,
            I => \VPP_VDDQ.count_2_rst_14\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__24095\,
            I => \VPP_VDDQ.count_2_rst_14\
        );

    \I__4124\ : InMux
    port map (
            O => \N__24090\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__4123\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24084\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__24084\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__4121\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24075\
        );

    \I__4120\ : InMux
    port map (
            O => \N__24080\,
            I => \N__24075\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__24075\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__4118\ : InMux
    port map (
            O => \N__24072\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__4117\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24066\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__24066\,
            I => \N__24063\
        );

    \I__4115\ : Span4Mux_h
    port map (
            O => \N__24063\,
            I => \N__24060\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__24060\,
            I => \VPP_VDDQ.un1_count_2_1_axb_12\
        );

    \I__4113\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24052\
        );

    \I__4112\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24047\
        );

    \I__4111\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24047\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__24052\,
            I => \N__24044\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__24047\,
            I => \N__24041\
        );

    \I__4108\ : Span4Mux_s2_v
    port map (
            O => \N__24044\,
            I => \N__24038\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__24041\,
            I => \N__24035\
        );

    \I__4106\ : Odrv4
    port map (
            O => \N__24038\,
            I => \VPP_VDDQ.count_2_rst_12\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__24035\,
            I => \VPP_VDDQ.count_2_rst_12\
        );

    \I__4104\ : InMux
    port map (
            O => \N__24030\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__4103\ : InMux
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__24024\,
            I => \N__24021\
        );

    \I__4101\ : Span4Mux_h
    port map (
            O => \N__24021\,
            I => \N__24018\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__24018\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__4099\ : InMux
    port map (
            O => \N__24015\,
            I => \N__24011\
        );

    \I__4098\ : InMux
    port map (
            O => \N__24014\,
            I => \N__24008\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__24011\,
            I => \N__24005\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__24008\,
            I => \N__24002\
        );

    \I__4095\ : Span4Mux_s2_v
    port map (
            O => \N__24005\,
            I => \N__23999\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__24002\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__23999\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__4092\ : InMux
    port map (
            O => \N__23994\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__4091\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23988\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__23988\,
            I => \N__23985\
        );

    \I__4089\ : Odrv4
    port map (
            O => \N__23985\,
            I => \VPP_VDDQ.un1_count_2_1_axb_14\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__23982\,
            I => \N__23979\
        );

    \I__4087\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23975\
        );

    \I__4086\ : InMux
    port map (
            O => \N__23978\,
            I => \N__23972\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__23975\,
            I => \N__23968\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__23972\,
            I => \N__23965\
        );

    \I__4083\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23962\
        );

    \I__4082\ : Span4Mux_h
    port map (
            O => \N__23968\,
            I => \N__23959\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__23965\,
            I => \N__23956\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__23962\,
            I => \N__23953\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__23959\,
            I => \VPP_VDDQ.count_2_rst_10\
        );

    \I__4078\ : Odrv4
    port map (
            O => \N__23956\,
            I => \VPP_VDDQ.count_2_rst_10\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__23953\,
            I => \VPP_VDDQ.count_2_rst_10\
        );

    \I__4076\ : InMux
    port map (
            O => \N__23946\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__4075\ : InMux
    port map (
            O => \N__23943\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__4074\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23935\
        );

    \I__4073\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23932\
        );

    \I__4072\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23929\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__23935\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__23932\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__23929\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__4068\ : InMux
    port map (
            O => \N__23922\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__4067\ : InMux
    port map (
            O => \N__23919\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__4066\ : InMux
    port map (
            O => \N__23916\,
            I => \N__23913\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__23913\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__4064\ : InMux
    port map (
            O => \N__23910\,
            I => \N__23907\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__23907\,
            I => \N__23903\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__23906\,
            I => \N__23900\
        );

    \I__4061\ : Span4Mux_s1_v
    port map (
            O => \N__23903\,
            I => \N__23897\
        );

    \I__4060\ : InMux
    port map (
            O => \N__23900\,
            I => \N__23894\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__23897\,
            I => \VPP_VDDQ.count_2_rst_4\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__23894\,
            I => \VPP_VDDQ.count_2_rst_4\
        );

    \I__4057\ : InMux
    port map (
            O => \N__23889\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__4056\ : InMux
    port map (
            O => \N__23886\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__4055\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23879\
        );

    \I__4054\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23876\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__23879\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__23876\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__4051\ : InMux
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__23868\,
            I => \N__23865\
        );

    \I__4049\ : Span4Mux_s1_v
    port map (
            O => \N__23865\,
            I => \N__23861\
        );

    \I__4048\ : InMux
    port map (
            O => \N__23864\,
            I => \N__23858\
        );

    \I__4047\ : Odrv4
    port map (
            O => \N__23861\,
            I => \VPP_VDDQ.count_2_rst_2\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__23858\,
            I => \VPP_VDDQ.count_2_rst_2\
        );

    \I__4045\ : InMux
    port map (
            O => \N__23853\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__4044\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23847\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__23847\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__4042\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23839\
        );

    \I__4041\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23834\
        );

    \I__4040\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23834\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__23839\,
            I => \VPP_VDDQ.count_2_rst_1\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__23834\,
            I => \VPP_VDDQ.count_2_rst_1\
        );

    \I__4037\ : InMux
    port map (
            O => \N__23829\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__4036\ : InMux
    port map (
            O => \N__23826\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__4035\ : CascadeMux
    port map (
            O => \N__23823\,
            I => \N__23820\
        );

    \I__4034\ : InMux
    port map (
            O => \N__23820\,
            I => \N__23817\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__23817\,
            I => \N__23814\
        );

    \I__4032\ : Span4Mux_h
    port map (
            O => \N__23814\,
            I => \N__23811\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__23811\,
            I => \POWERLED.un1_dutycycle_53_axb_13_1\
        );

    \I__4030\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23803\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__23807\,
            I => \N__23800\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__23806\,
            I => \N__23787\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__23803\,
            I => \N__23784\
        );

    \I__4026\ : InMux
    port map (
            O => \N__23800\,
            I => \N__23779\
        );

    \I__4025\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23779\
        );

    \I__4024\ : InMux
    port map (
            O => \N__23798\,
            I => \N__23774\
        );

    \I__4023\ : InMux
    port map (
            O => \N__23797\,
            I => \N__23774\
        );

    \I__4022\ : InMux
    port map (
            O => \N__23796\,
            I => \N__23767\
        );

    \I__4021\ : InMux
    port map (
            O => \N__23795\,
            I => \N__23767\
        );

    \I__4020\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23767\
        );

    \I__4019\ : InMux
    port map (
            O => \N__23793\,
            I => \N__23756\
        );

    \I__4018\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23756\
        );

    \I__4017\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23756\
        );

    \I__4016\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23756\
        );

    \I__4015\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23756\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__23784\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_7\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__23779\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_7\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__23774\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_7\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__23767\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_7\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__23756\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_7\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__4008\ : InMux
    port map (
            O => \N__23742\,
            I => \N__23739\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__4006\ : Span4Mux_h
    port map (
            O => \N__23736\,
            I => \N__23733\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__23733\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__4004\ : InMux
    port map (
            O => \N__23730\,
            I => \N__23727\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__23727\,
            I => \N__23724\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__23724\,
            I => \VPP_VDDQ.count_2_0_4\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__23721\,
            I => \VPP_VDDQ.count_2Z0Z_4_cascade_\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__23718\,
            I => \VPP_VDDQ.count_2_rst_8_cascade_\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__23715\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__23712\,
            I => \VPP_VDDQ.count_2_rst_7_cascade_\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__23709\,
            I => \VPP_VDDQ.count_2Z0Z_1_cascade_\
        );

    \I__3996\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23703\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__23703\,
            I => \VPP_VDDQ.count_2_0_1\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__23700\,
            I => \N__23695\
        );

    \I__3993\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23687\
        );

    \I__3992\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23687\
        );

    \I__3991\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23680\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__23694\,
            I => \N__23675\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__23693\,
            I => \N__23671\
        );

    \I__3988\ : InMux
    port map (
            O => \N__23692\,
            I => \N__23664\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__23687\,
            I => \N__23661\
        );

    \I__3986\ : InMux
    port map (
            O => \N__23686\,
            I => \N__23654\
        );

    \I__3985\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23654\
        );

    \I__3984\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23654\
        );

    \I__3983\ : InMux
    port map (
            O => \N__23683\,
            I => \N__23651\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__23680\,
            I => \N__23648\
        );

    \I__3981\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23640\
        );

    \I__3980\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23640\
        );

    \I__3979\ : InMux
    port map (
            O => \N__23675\,
            I => \N__23637\
        );

    \I__3978\ : InMux
    port map (
            O => \N__23674\,
            I => \N__23634\
        );

    \I__3977\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23629\
        );

    \I__3976\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23629\
        );

    \I__3975\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23624\
        );

    \I__3974\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23624\
        );

    \I__3973\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23621\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__23664\,
            I => \N__23614\
        );

    \I__3971\ : Span4Mux_s3_v
    port map (
            O => \N__23661\,
            I => \N__23614\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__23654\,
            I => \N__23614\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__23651\,
            I => \N__23611\
        );

    \I__3968\ : Span4Mux_h
    port map (
            O => \N__23648\,
            I => \N__23608\
        );

    \I__3967\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23603\
        );

    \I__3966\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23603\
        );

    \I__3965\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23600\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23591\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__23637\,
            I => \N__23591\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__23634\,
            I => \N__23591\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__23629\,
            I => \N__23591\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23584\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23584\
        );

    \I__3958\ : Span4Mux_h
    port map (
            O => \N__23614\,
            I => \N__23584\
        );

    \I__3957\ : Span4Mux_v
    port map (
            O => \N__23611\,
            I => \N__23581\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__23608\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__23603\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__23600\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__3953\ : Odrv12
    port map (
            O => \N__23591\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__3952\ : Odrv4
    port map (
            O => \N__23584\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__23581\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__23568\,
            I => \POWERLED.N_161_N_cascade_\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__23565\,
            I => \N__23562\
        );

    \I__3948\ : InMux
    port map (
            O => \N__23562\,
            I => \N__23559\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__23559\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__3946\ : InMux
    port map (
            O => \N__23556\,
            I => \N__23550\
        );

    \I__3945\ : InMux
    port map (
            O => \N__23555\,
            I => \N__23550\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__23550\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__3943\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23530\
        );

    \I__3942\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23517\
        );

    \I__3941\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23514\
        );

    \I__3940\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23507\
        );

    \I__3939\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23507\
        );

    \I__3938\ : InMux
    port map (
            O => \N__23542\,
            I => \N__23507\
        );

    \I__3937\ : InMux
    port map (
            O => \N__23541\,
            I => \N__23500\
        );

    \I__3936\ : InMux
    port map (
            O => \N__23540\,
            I => \N__23500\
        );

    \I__3935\ : InMux
    port map (
            O => \N__23539\,
            I => \N__23500\
        );

    \I__3934\ : InMux
    port map (
            O => \N__23538\,
            I => \N__23491\
        );

    \I__3933\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23491\
        );

    \I__3932\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23491\
        );

    \I__3931\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23491\
        );

    \I__3930\ : InMux
    port map (
            O => \N__23534\,
            I => \N__23486\
        );

    \I__3929\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23486\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__23530\,
            I => \N__23483\
        );

    \I__3927\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23480\
        );

    \I__3926\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23475\
        );

    \I__3925\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23475\
        );

    \I__3924\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23466\
        );

    \I__3923\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23466\
        );

    \I__3922\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23466\
        );

    \I__3921\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23466\
        );

    \I__3920\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23463\
        );

    \I__3919\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23458\
        );

    \I__3918\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23458\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__23517\,
            I => \N__23444\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23441\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__23507\,
            I => \N__23436\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__23500\,
            I => \N__23436\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__23491\,
            I => \N__23423\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23423\
        );

    \I__3911\ : Span4Mux_s1_v
    port map (
            O => \N__23483\,
            I => \N__23423\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__23480\,
            I => \N__23423\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23423\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__23466\,
            I => \N__23423\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__23463\,
            I => \N__23417\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__23458\,
            I => \N__23417\
        );

    \I__3905\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23414\
        );

    \I__3904\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23405\
        );

    \I__3903\ : InMux
    port map (
            O => \N__23455\,
            I => \N__23405\
        );

    \I__3902\ : InMux
    port map (
            O => \N__23454\,
            I => \N__23405\
        );

    \I__3901\ : InMux
    port map (
            O => \N__23453\,
            I => \N__23405\
        );

    \I__3900\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23402\
        );

    \I__3899\ : InMux
    port map (
            O => \N__23451\,
            I => \N__23399\
        );

    \I__3898\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23390\
        );

    \I__3897\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23390\
        );

    \I__3896\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23390\
        );

    \I__3895\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23390\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__23444\,
            I => \N__23381\
        );

    \I__3893\ : Span4Mux_v
    port map (
            O => \N__23441\,
            I => \N__23381\
        );

    \I__3892\ : Span4Mux_v
    port map (
            O => \N__23436\,
            I => \N__23381\
        );

    \I__3891\ : Span4Mux_v
    port map (
            O => \N__23423\,
            I => \N__23381\
        );

    \I__3890\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23378\
        );

    \I__3889\ : Span4Mux_s3_v
    port map (
            O => \N__23417\,
            I => \N__23375\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23370\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__23405\,
            I => \N__23370\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__23402\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__23399\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__23390\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3883\ : Odrv4
    port map (
            O => \N__23381\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__23378\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__23375\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3880\ : Odrv12
    port map (
            O => \N__23370\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__23355\,
            I => \POWERLED.dutycycle_en_12_cascade_\
        );

    \I__3878\ : InMux
    port map (
            O => \N__23352\,
            I => \N__23346\
        );

    \I__3877\ : InMux
    port map (
            O => \N__23351\,
            I => \N__23346\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__23346\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__3875\ : SRMux
    port map (
            O => \N__23343\,
            I => \N__23338\
        );

    \I__3874\ : SRMux
    port map (
            O => \N__23342\,
            I => \N__23331\
        );

    \I__3873\ : SRMux
    port map (
            O => \N__23341\,
            I => \N__23327\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__23338\,
            I => \N__23324\
        );

    \I__3871\ : SRMux
    port map (
            O => \N__23337\,
            I => \N__23321\
        );

    \I__3870\ : SRMux
    port map (
            O => \N__23336\,
            I => \N__23318\
        );

    \I__3869\ : SRMux
    port map (
            O => \N__23335\,
            I => \N__23315\
        );

    \I__3868\ : SRMux
    port map (
            O => \N__23334\,
            I => \N__23312\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__23331\,
            I => \N__23308\
        );

    \I__3866\ : SRMux
    port map (
            O => \N__23330\,
            I => \N__23305\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23298\
        );

    \I__3864\ : Span4Mux_s3_v
    port map (
            O => \N__23324\,
            I => \N__23298\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__23321\,
            I => \N__23298\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23294\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23291\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23288\
        );

    \I__3859\ : SRMux
    port map (
            O => \N__23311\,
            I => \N__23285\
        );

    \I__3858\ : Span4Mux_v
    port map (
            O => \N__23308\,
            I => \N__23282\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23277\
        );

    \I__3856\ : Span4Mux_h
    port map (
            O => \N__23298\,
            I => \N__23277\
        );

    \I__3855\ : SRMux
    port map (
            O => \N__23297\,
            I => \N__23274\
        );

    \I__3854\ : Span4Mux_v
    port map (
            O => \N__23294\,
            I => \N__23269\
        );

    \I__3853\ : Span4Mux_v
    port map (
            O => \N__23291\,
            I => \N__23269\
        );

    \I__3852\ : Span4Mux_s2_h
    port map (
            O => \N__23288\,
            I => \N__23266\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__23285\,
            I => \N__23263\
        );

    \I__3850\ : Span4Mux_h
    port map (
            O => \N__23282\,
            I => \N__23260\
        );

    \I__3849\ : Span4Mux_s2_h
    port map (
            O => \N__23277\,
            I => \N__23257\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__23274\,
            I => \N__23252\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__23269\,
            I => \N__23252\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__23266\,
            I => \POWERLED.N_229_iZ0\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__23263\,
            I => \POWERLED.N_229_iZ0\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__23260\,
            I => \POWERLED.N_229_iZ0\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__23257\,
            I => \POWERLED.N_229_iZ0\
        );

    \I__3842\ : Odrv4
    port map (
            O => \N__23252\,
            I => \POWERLED.N_229_iZ0\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__23241\,
            I => \POWERLED.un1_dutycycle_53_49_0_1_cascade_\
        );

    \I__3840\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__23235\,
            I => \POWERLED.un1_dutycycle_53_49_0_0\
        );

    \I__3838\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23226\
        );

    \I__3837\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23226\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__23226\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_6\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__23223\,
            I => \POWERLED.un1_dutycycle_53_9_1_cascade_\
        );

    \I__3834\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23217\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__23217\,
            I => \POWERLED.un1_dutycycle_53_2_1_0_tz\
        );

    \I__3832\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23199\
        );

    \I__3831\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23192\
        );

    \I__3830\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23192\
        );

    \I__3829\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23192\
        );

    \I__3828\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23187\
        );

    \I__3827\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23187\
        );

    \I__3826\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23184\
        );

    \I__3825\ : InMux
    port map (
            O => \N__23207\,
            I => \N__23173\
        );

    \I__3824\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23173\
        );

    \I__3823\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23173\
        );

    \I__3822\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23173\
        );

    \I__3821\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23173\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__23202\,
            I => \N__23165\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23161\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__23192\,
            I => \N__23158\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__23187\,
            I => \N__23155\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__23184\,
            I => \N__23152\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__23173\,
            I => \N__23149\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__23172\,
            I => \N__23144\
        );

    \I__3813\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23141\
        );

    \I__3812\ : InMux
    port map (
            O => \N__23170\,
            I => \N__23130\
        );

    \I__3811\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23130\
        );

    \I__3810\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23130\
        );

    \I__3809\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23130\
        );

    \I__3808\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23130\
        );

    \I__3807\ : Span4Mux_s2_h
    port map (
            O => \N__23161\,
            I => \N__23119\
        );

    \I__3806\ : Span4Mux_s1_v
    port map (
            O => \N__23158\,
            I => \N__23119\
        );

    \I__3805\ : Span4Mux_s2_h
    port map (
            O => \N__23155\,
            I => \N__23119\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__23152\,
            I => \N__23119\
        );

    \I__3803\ : Span4Mux_s1_v
    port map (
            O => \N__23149\,
            I => \N__23119\
        );

    \I__3802\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23114\
        );

    \I__3801\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23114\
        );

    \I__3800\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23111\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__23141\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__23130\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__23119\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__23114\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__23111\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__23100\,
            I => \POWERLED.dutycycleZ0Z_11_cascade_\
        );

    \I__3793\ : InMux
    port map (
            O => \N__23097\,
            I => \N__23094\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__23094\,
            I => \POWERLED.un1_i1_mux\
        );

    \I__3791\ : InMux
    port map (
            O => \N__23091\,
            I => \N__23088\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__23088\,
            I => \N__23085\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__23085\,
            I => \N__23082\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__23082\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_7\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__23079\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_11_cascade_\
        );

    \I__3786\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23073\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__23073\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_7\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__23070\,
            I => \POWERLED.un1_dutycycle_53_axb_12_cascade_\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__23067\,
            I => \POWERLED.dutycycleZ0Z_10_cascade_\
        );

    \I__3782\ : CascadeMux
    port map (
            O => \N__23064\,
            I => \POWERLED.N_156_N_cascade_\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__3780\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__23055\,
            I => \POWERLED.dutycycle_en_10\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__23052\,
            I => \POWERLED.dutycycle_en_10_cascade_\
        );

    \I__3777\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23045\
        );

    \I__3776\ : InMux
    port map (
            O => \N__23048\,
            I => \N__23042\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__23045\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__23042\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__3773\ : InMux
    port map (
            O => \N__23037\,
            I => \N__23033\
        );

    \I__3772\ : InMux
    port map (
            O => \N__23036\,
            I => \N__23030\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__23033\,
            I => \POWERLED.dutycycleZ1Z_13\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__23030\,
            I => \POWERLED.dutycycleZ1Z_13\
        );

    \I__3769\ : CascadeMux
    port map (
            O => \N__23025\,
            I => \POWERLED.dutycycleZ0Z_13_cascade_\
        );

    \I__3768\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23016\
        );

    \I__3767\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23016\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__23016\,
            I => \N__23008\
        );

    \I__3765\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23005\
        );

    \I__3764\ : InMux
    port map (
            O => \N__23014\,
            I => \N__23000\
        );

    \I__3763\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23000\
        );

    \I__3762\ : InMux
    port map (
            O => \N__23012\,
            I => \N__22993\
        );

    \I__3761\ : InMux
    port map (
            O => \N__23011\,
            I => \N__22993\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__23008\,
            I => \N__22988\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__23005\,
            I => \N__22988\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__23000\,
            I => \N__22985\
        );

    \I__3757\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22980\
        );

    \I__3756\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22980\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__22993\,
            I => \N__22977\
        );

    \I__3754\ : Span4Mux_s3_v
    port map (
            O => \N__22988\,
            I => \N__22972\
        );

    \I__3753\ : Span4Mux_s3_v
    port map (
            O => \N__22985\,
            I => \N__22972\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__22980\,
            I => \POWERLED.N_143_N\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__22977\,
            I => \POWERLED.N_143_N\
        );

    \I__3750\ : Odrv4
    port map (
            O => \N__22972\,
            I => \POWERLED.N_143_N\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__22965\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__3748\ : CascadeMux
    port map (
            O => \N__22962\,
            I => \POWERLED.N_158_N_cascade_\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__22959\,
            I => \N__22956\
        );

    \I__3746\ : InMux
    port map (
            O => \N__22956\,
            I => \N__22953\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__22953\,
            I => \POWERLED.dutycycle_en_11\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__22950\,
            I => \POWERLED.dutycycle_en_11_cascade_\
        );

    \I__3743\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22943\
        );

    \I__3742\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22940\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__22943\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__22940\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__3739\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22932\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__22932\,
            I => \N__22929\
        );

    \I__3737\ : Span4Mux_h
    port map (
            O => \N__22929\,
            I => \N__22926\
        );

    \I__3736\ : Span4Mux_s3_h
    port map (
            O => \N__22926\,
            I => \N__22922\
        );

    \I__3735\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22919\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__22922\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__22919\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__22914\,
            I => \N__22911\
        );

    \I__3731\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22905\
        );

    \I__3730\ : InMux
    port map (
            O => \N__22910\,
            I => \N__22905\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__22905\,
            I => \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HHZ0Z1\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__22902\,
            I => \N__22898\
        );

    \I__3727\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22893\
        );

    \I__3726\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22893\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__22893\,
            I => \POWERLED.dutycycleZ1Z_11\
        );

    \I__3724\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22884\
        );

    \I__3723\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22884\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__22884\,
            I => \N__22881\
        );

    \I__3721\ : Odrv12
    port map (
            O => \N__22881\,
            I => \POWERLED.dutycycle_eena_7\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__22878\,
            I => \POWERLED.dutycycleZ0Z_8_cascade_\
        );

    \I__3719\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22869\
        );

    \I__3718\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22869\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__22869\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__3716\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22862\
        );

    \I__3715\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22859\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__22862\,
            I => \N__22854\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__22859\,
            I => \N__22854\
        );

    \I__3712\ : Odrv12
    port map (
            O => \N__22854\,
            I => \POWERLED.dutycycle_eena_9\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__22851\,
            I => \N__22848\
        );

    \I__3710\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22842\
        );

    \I__3709\ : InMux
    port map (
            O => \N__22847\,
            I => \N__22842\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__22842\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__22839\,
            I => \N__22834\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__22838\,
            I => \N__22831\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__22837\,
            I => \N__22828\
        );

    \I__3704\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22818\
        );

    \I__3703\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22818\
        );

    \I__3702\ : InMux
    port map (
            O => \N__22828\,
            I => \N__22818\
        );

    \I__3701\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22815\
        );

    \I__3700\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22812\
        );

    \I__3699\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22809\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22803\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22803\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22798\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22798\
        );

    \I__3694\ : CascadeMux
    port map (
            O => \N__22808\,
            I => \N__22795\
        );

    \I__3693\ : Span4Mux_v
    port map (
            O => \N__22803\,
            I => \N__22790\
        );

    \I__3692\ : Span4Mux_v
    port map (
            O => \N__22798\,
            I => \N__22790\
        );

    \I__3691\ : InMux
    port map (
            O => \N__22795\,
            I => \N__22787\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__22790\,
            I => \POWERLED.N_164\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__22787\,
            I => \POWERLED.N_164\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__22782\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\
        );

    \I__3687\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22776\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__22776\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_1_0\
        );

    \I__3685\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22769\
        );

    \I__3684\ : InMux
    port map (
            O => \N__22772\,
            I => \N__22766\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__22769\,
            I => \N__22763\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__22766\,
            I => \N__22760\
        );

    \I__3681\ : Odrv4
    port map (
            O => \N__22763\,
            I => \POWERLED.N_228\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__22760\,
            I => \POWERLED.N_228\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__22755\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\
        );

    \I__3678\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22737\
        );

    \I__3677\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22737\
        );

    \I__3676\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22730\
        );

    \I__3675\ : InMux
    port map (
            O => \N__22749\,
            I => \N__22727\
        );

    \I__3674\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22724\
        );

    \I__3673\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22720\
        );

    \I__3672\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22717\
        );

    \I__3671\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22712\
        );

    \I__3670\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22712\
        );

    \I__3669\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22709\
        );

    \I__3668\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22706\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__22737\,
            I => \N__22703\
        );

    \I__3666\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22694\
        );

    \I__3665\ : InMux
    port map (
            O => \N__22735\,
            I => \N__22694\
        );

    \I__3664\ : InMux
    port map (
            O => \N__22734\,
            I => \N__22694\
        );

    \I__3663\ : InMux
    port map (
            O => \N__22733\,
            I => \N__22694\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__22730\,
            I => \N__22680\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22680\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__22724\,
            I => \N__22680\
        );

    \I__3659\ : InMux
    port map (
            O => \N__22723\,
            I => \N__22677\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22672\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22672\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__22712\,
            I => \N__22665\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__22709\,
            I => \N__22665\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__22706\,
            I => \N__22665\
        );

    \I__3653\ : Span4Mux_v
    port map (
            O => \N__22703\,
            I => \N__22660\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__22694\,
            I => \N__22660\
        );

    \I__3651\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22657\
        );

    \I__3650\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22654\
        );

    \I__3649\ : InMux
    port map (
            O => \N__22691\,
            I => \N__22647\
        );

    \I__3648\ : InMux
    port map (
            O => \N__22690\,
            I => \N__22647\
        );

    \I__3647\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22647\
        );

    \I__3646\ : InMux
    port map (
            O => \N__22688\,
            I => \N__22642\
        );

    \I__3645\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22642\
        );

    \I__3644\ : Span4Mux_v
    port map (
            O => \N__22680\,
            I => \N__22639\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__22677\,
            I => \N__22628\
        );

    \I__3642\ : Span4Mux_v
    port map (
            O => \N__22672\,
            I => \N__22628\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__22665\,
            I => \N__22628\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__22660\,
            I => \N__22628\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__22657\,
            I => \N__22628\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__22654\,
            I => \POWERLED.func_state\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__22647\,
            I => \POWERLED.func_state\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__22642\,
            I => \POWERLED.func_state\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__22639\,
            I => \POWERLED.func_state\
        );

    \I__3634\ : Odrv4
    port map (
            O => \N__22628\,
            I => \POWERLED.func_state\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__22617\,
            I => \N__22608\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \N__22603\
        );

    \I__3631\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22596\
        );

    \I__3630\ : InMux
    port map (
            O => \N__22614\,
            I => \N__22596\
        );

    \I__3629\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22589\
        );

    \I__3628\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22589\
        );

    \I__3627\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22589\
        );

    \I__3626\ : InMux
    port map (
            O => \N__22608\,
            I => \N__22582\
        );

    \I__3625\ : InMux
    port map (
            O => \N__22607\,
            I => \N__22582\
        );

    \I__3624\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22582\
        );

    \I__3623\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22577\
        );

    \I__3622\ : InMux
    port map (
            O => \N__22602\,
            I => \N__22577\
        );

    \I__3621\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22574\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__22596\,
            I => \N__22569\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__22589\,
            I => \N__22569\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__22582\,
            I => \N__22564\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22564\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__22574\,
            I => \N__22561\
        );

    \I__3615\ : Span4Mux_v
    port map (
            O => \N__22569\,
            I => \N__22556\
        );

    \I__3614\ : Span4Mux_v
    port map (
            O => \N__22564\,
            I => \N__22556\
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__22561\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__22556\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3611\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22546\
        );

    \I__3610\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22543\
        );

    \I__3609\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22540\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__22546\,
            I => \N__22537\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22534\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__22540\,
            I => \N__22530\
        );

    \I__3605\ : Span4Mux_h
    port map (
            O => \N__22537\,
            I => \N__22527\
        );

    \I__3604\ : Span4Mux_h
    port map (
            O => \N__22534\,
            I => \N__22524\
        );

    \I__3603\ : InMux
    port map (
            O => \N__22533\,
            I => \N__22521\
        );

    \I__3602\ : Odrv12
    port map (
            O => \N__22530\,
            I => \POWERLED.func_state_RNI_0Z0Z_1\
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__22527\,
            I => \POWERLED.func_state_RNI_0Z0Z_1\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__22524\,
            I => \POWERLED.func_state_RNI_0Z0Z_1\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__22521\,
            I => \POWERLED.func_state_RNI_0Z0Z_1\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__22512\,
            I => \POWERLED.dutycycle_eena_5_d_cascade_\
        );

    \I__3597\ : InMux
    port map (
            O => \N__22509\,
            I => \N__22506\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22503\
        );

    \I__3595\ : Span4Mux_h
    port map (
            O => \N__22503\,
            I => \N__22500\
        );

    \I__3594\ : Odrv4
    port map (
            O => \N__22500\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0\
        );

    \I__3593\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22494\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__22494\,
            I => \POWERLED.dutycycle_RNIB8FGCZ0Z_7\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__22491\,
            I => \N__22488\
        );

    \I__3590\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22482\
        );

    \I__3589\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22482\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__22482\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__22479\,
            I => \POWERLED.dutycycle_RNIB8FGCZ0Z_7_cascade_\
        );

    \I__3586\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22470\
        );

    \I__3585\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22470\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__22470\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__22467\,
            I => \N__22464\
        );

    \I__3582\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22461\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__22461\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1\
        );

    \I__3580\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22454\
        );

    \I__3579\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22451\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__22454\,
            I => \N__22448\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__22451\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__22448\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__22443\,
            I => \POWERLED.count_clkZ0Z_8_cascade_\
        );

    \I__3574\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22433\
        );

    \I__3573\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22433\
        );

    \I__3572\ : InMux
    port map (
            O => \N__22438\,
            I => \N__22430\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__22433\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__22430\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__3569\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22419\
        );

    \I__3568\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22419\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__22419\,
            I => \N__22415\
        );

    \I__3566\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22412\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__22415\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__22412\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__22407\,
            I => \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\
        );

    \I__3562\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22398\
        );

    \I__3561\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22398\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__22398\,
            I => \N__22395\
        );

    \I__3559\ : Odrv4
    port map (
            O => \N__22395\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__3557\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22386\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__22386\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__3555\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22378\
        );

    \I__3554\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22373\
        );

    \I__3553\ : InMux
    port map (
            O => \N__22381\,
            I => \N__22373\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__22378\,
            I => \N__22370\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__22373\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__22370\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__3549\ : InMux
    port map (
            O => \N__22365\,
            I => \N__22359\
        );

    \I__3548\ : InMux
    port map (
            O => \N__22364\,
            I => \N__22359\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__22356\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__3544\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22347\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__22347\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__3542\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__3540\ : Span4Mux_s2_v
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__22335\,
            I => \POWERLED.un1_N_1_i\
        );

    \I__3538\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22326\
        );

    \I__3537\ : InMux
    port map (
            O => \N__22331\,
            I => \N__22326\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__3535\ : Span12Mux_s4_v
    port map (
            O => \N__22323\,
            I => \N__22320\
        );

    \I__3534\ : Odrv12
    port map (
            O => \N__22320\,
            I => \POWERLED.g3_0_3_0_0\
        );

    \I__3533\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22313\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22310\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22307\
        );

    \I__3530\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22304\
        );

    \I__3529\ : Odrv4
    port map (
            O => \N__22307\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__22304\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__3527\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22293\
        );

    \I__3526\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22293\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__22293\,
            I => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\
        );

    \I__3524\ : InMux
    port map (
            O => \N__22290\,
            I => \POWERLED.un1_count_clk_2_cry_9\
        );

    \I__3523\ : InMux
    port map (
            O => \N__22287\,
            I => \N__22283\
        );

    \I__3522\ : InMux
    port map (
            O => \N__22286\,
            I => \N__22280\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__22283\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__22280\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__3519\ : InMux
    port map (
            O => \N__22275\,
            I => \N__22269\
        );

    \I__3518\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22269\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__22269\,
            I => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\
        );

    \I__3516\ : InMux
    port map (
            O => \N__22266\,
            I => \POWERLED.un1_count_clk_2_cry_10\
        );

    \I__3515\ : InMux
    port map (
            O => \N__22263\,
            I => \N__22259\
        );

    \I__3514\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22256\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__22259\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__22256\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__3511\ : InMux
    port map (
            O => \N__22251\,
            I => \POWERLED.un1_count_clk_2_cry_11\
        );

    \I__3510\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22245\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__22245\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__3508\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22236\
        );

    \I__3507\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22236\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__22236\,
            I => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\
        );

    \I__3505\ : InMux
    port map (
            O => \N__22233\,
            I => \POWERLED.un1_count_clk_2_cry_12\
        );

    \I__3504\ : InMux
    port map (
            O => \N__22230\,
            I => \POWERLED.un1_count_clk_2_cry_13\
        );

    \I__3503\ : InMux
    port map (
            O => \N__22227\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__3502\ : InMux
    port map (
            O => \N__22224\,
            I => \N__22220\
        );

    \I__3501\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22217\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__22220\,
            I => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__22217\,
            I => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__22212\,
            I => \N__22209\
        );

    \I__3497\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22206\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__22206\,
            I => \N__22203\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__22203\,
            I => \POWERLED.count_clk_0_12\
        );

    \I__3494\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22194\
        );

    \I__3493\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22194\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__22194\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__3491\ : InMux
    port map (
            O => \N__22191\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__3490\ : InMux
    port map (
            O => \N__22188\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__3489\ : InMux
    port map (
            O => \N__22185\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__3488\ : InMux
    port map (
            O => \N__22182\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__3487\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22173\
        );

    \I__3486\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22173\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__22173\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__3484\ : InMux
    port map (
            O => \N__22170\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__3483\ : InMux
    port map (
            O => \N__22167\,
            I => \N__22161\
        );

    \I__3482\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22161\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__22161\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__3480\ : InMux
    port map (
            O => \N__22158\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__3479\ : InMux
    port map (
            O => \N__22155\,
            I => \POWERLED.un1_count_clk_2_cry_7\
        );

    \I__3478\ : InMux
    port map (
            O => \N__22152\,
            I => \bfn_6_10_0_\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__22149\,
            I => \N__22146\
        );

    \I__3476\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22140\
        );

    \I__3475\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22140\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__22140\,
            I => \POWERLED.count_off_1_13\
        );

    \I__3473\ : InMux
    port map (
            O => \N__22137\,
            I => \N__22134\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__22134\,
            I => \POWERLED.count_off_0_13\
        );

    \I__3471\ : CascadeMux
    port map (
            O => \N__22131\,
            I => \N__22128\
        );

    \I__3470\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22122\
        );

    \I__3469\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22122\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__22122\,
            I => \POWERLED.count_off_1_14\
        );

    \I__3467\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__22116\,
            I => \POWERLED.count_off_0_14\
        );

    \I__3465\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22107\
        );

    \I__3464\ : InMux
    port map (
            O => \N__22112\,
            I => \N__22107\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__22107\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIPVUTZ0Z2\
        );

    \I__3462\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22101\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__22101\,
            I => \POWERLED.count_off_0_15\
        );

    \I__3460\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22095\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__22095\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__3458\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22088\
        );

    \I__3457\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22085\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__22088\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__22085\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3454\ : InMux
    port map (
            O => \N__22080\,
            I => \N__22076\
        );

    \I__3453\ : InMux
    port map (
            O => \N__22079\,
            I => \N__22073\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__22076\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__22073\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__22068\,
            I => \POWERLED.count_offZ0Z_15_cascade_\
        );

    \I__3449\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22061\
        );

    \I__3448\ : InMux
    port map (
            O => \N__22064\,
            I => \N__22058\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__22061\,
            I => \N__22055\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__22058\,
            I => \N__22050\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__22055\,
            I => \N__22047\
        );

    \I__3444\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22042\
        );

    \I__3443\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22042\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__22050\,
            I => \N__22039\
        );

    \I__3441\ : Odrv4
    port map (
            O => \N__22047\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__22042\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3439\ : Odrv4
    port map (
            O => \N__22039\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3438\ : InMux
    port map (
            O => \N__22032\,
            I => \N__22029\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__22029\,
            I => \POWERLED.un34_clk_100khz_10\
        );

    \I__3436\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22023\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22020\
        );

    \I__3434\ : Span4Mux_h
    port map (
            O => \N__22020\,
            I => \N__22017\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__22017\,
            I => \POWERLED.count_off_0_6\
        );

    \I__3432\ : InMux
    port map (
            O => \N__22014\,
            I => \N__22010\
        );

    \I__3431\ : InMux
    port map (
            O => \N__22013\,
            I => \N__22007\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__22010\,
            I => \N__22004\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__22007\,
            I => \POWERLED.count_off_1_6\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__22004\,
            I => \POWERLED.count_off_1_6\
        );

    \I__3427\ : InMux
    port map (
            O => \N__21999\,
            I => \N__21995\
        );

    \I__3426\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21992\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__21995\,
            I => \N__21989\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__21992\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__21989\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__21984\,
            I => \N__21981\
        );

    \I__3421\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21975\
        );

    \I__3420\ : InMux
    port map (
            O => \N__21980\,
            I => \N__21975\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__21975\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__21972\,
            I => \N__21969\
        );

    \I__3417\ : InMux
    port map (
            O => \N__21969\,
            I => \N__21963\
        );

    \I__3416\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21963\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__21963\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__21960\,
            I => \N__21956\
        );

    \I__3413\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21951\
        );

    \I__3412\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21951\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__21951\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3410\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21944\
        );

    \I__3409\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21941\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__21944\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__21941\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__21936\,
            I => \N__21933\
        );

    \I__3405\ : InMux
    port map (
            O => \N__21933\,
            I => \N__21930\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__21930\,
            I => \N__21927\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__21927\,
            I => \N__21924\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__21924\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__3401\ : InMux
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__21918\,
            I => \POWERLED.count_off_0_9\
        );

    \I__3399\ : InMux
    port map (
            O => \N__21915\,
            I => \N__21909\
        );

    \I__3398\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21909\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__21909\,
            I => \POWERLED.count_off_1_9\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__21906\,
            I => \N__21903\
        );

    \I__3395\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21900\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__21900\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__21897\,
            I => \POWERLED.count_offZ0Z_9_cascade_\
        );

    \I__3392\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21891\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__21891\,
            I => \POWERLED.un34_clk_100khz_11\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__21888\,
            I => \N__21884\
        );

    \I__3389\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21881\
        );

    \I__3388\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21878\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__21881\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__21878\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3385\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21867\
        );

    \I__3384\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21867\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__21867\,
            I => \POWERLED.count_off_1_10\
        );

    \I__3382\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__21861\,
            I => \POWERLED.count_off_0_10\
        );

    \I__3380\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21854\
        );

    \I__3379\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21851\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__21854\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__21851\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3376\ : InMux
    port map (
            O => \N__21846\,
            I => \N__21840\
        );

    \I__3375\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21840\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__21840\,
            I => \POWERLED.count_off_1_11\
        );

    \I__3373\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21834\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__21834\,
            I => \POWERLED.count_off_0_11\
        );

    \I__3371\ : InMux
    port map (
            O => \N__21831\,
            I => \N__21828\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__21828\,
            I => \POWERLED.count_off_0_12\
        );

    \I__3369\ : InMux
    port map (
            O => \N__21825\,
            I => \N__21821\
        );

    \I__3368\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21818\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__21821\,
            I => \POWERLED.count_off_1_12\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__21818\,
            I => \POWERLED.count_off_1_12\
        );

    \I__3365\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21809\
        );

    \I__3364\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21806\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__21809\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__21806\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__21801\,
            I => \N__21797\
        );

    \I__3360\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21794\
        );

    \I__3359\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21791\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__21794\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__21791\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3356\ : InMux
    port map (
            O => \N__21786\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__3355\ : InMux
    port map (
            O => \N__21783\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__3354\ : InMux
    port map (
            O => \N__21780\,
            I => \bfn_6_6_0_\
        );

    \I__3353\ : InMux
    port map (
            O => \N__21777\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__3352\ : InMux
    port map (
            O => \N__21774\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__3351\ : InMux
    port map (
            O => \N__21771\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__3350\ : InMux
    port map (
            O => \N__21768\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__3349\ : InMux
    port map (
            O => \N__21765\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__3348\ : InMux
    port map (
            O => \N__21762\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__3347\ : InMux
    port map (
            O => \N__21759\,
            I => \N__21755\
        );

    \I__3346\ : InMux
    port map (
            O => \N__21758\,
            I => \N__21752\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__21755\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__21752\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3343\ : InMux
    port map (
            O => \N__21747\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__21744\,
            I => \N__21740\
        );

    \I__3341\ : InMux
    port map (
            O => \N__21743\,
            I => \N__21737\
        );

    \I__3340\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21734\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__21737\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__21734\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3337\ : InMux
    port map (
            O => \N__21729\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__3336\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21722\
        );

    \I__3335\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21719\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__21722\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__21719\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3332\ : InMux
    port map (
            O => \N__21714\,
            I => \bfn_6_5_0_\
        );

    \I__3331\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21707\
        );

    \I__3330\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21704\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__21707\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__21704\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3327\ : InMux
    port map (
            O => \N__21699\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__3326\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21692\
        );

    \I__3325\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21689\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__21692\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__21689\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3322\ : InMux
    port map (
            O => \N__21684\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__3321\ : InMux
    port map (
            O => \N__21681\,
            I => \N__21677\
        );

    \I__3320\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21674\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__21677\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__21674\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3317\ : InMux
    port map (
            O => \N__21669\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__3316\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21662\
        );

    \I__3315\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21659\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__21662\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__21659\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3312\ : InMux
    port map (
            O => \N__21654\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__3311\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21647\
        );

    \I__3310\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21644\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__21647\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__21644\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3307\ : InMux
    port map (
            O => \N__21639\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__3306\ : InMux
    port map (
            O => \N__21636\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__3305\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21629\
        );

    \I__3304\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21626\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__21629\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__21626\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3301\ : InMux
    port map (
            O => \N__21621\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__3300\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21614\
        );

    \I__3299\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21611\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__21614\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__21611\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3296\ : InMux
    port map (
            O => \N__21606\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__3295\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21599\
        );

    \I__3294\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21596\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__21599\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__21596\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3291\ : InMux
    port map (
            O => \N__21591\,
            I => \bfn_6_4_0_\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__21588\,
            I => \N__21584\
        );

    \I__3289\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21581\
        );

    \I__3288\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21578\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__21581\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__21578\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3285\ : InMux
    port map (
            O => \N__21573\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__3284\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21566\
        );

    \I__3283\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21563\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__21566\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__21563\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3280\ : InMux
    port map (
            O => \N__21558\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__3279\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21551\
        );

    \I__3278\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21548\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__21551\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__21548\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3275\ : InMux
    port map (
            O => \N__21543\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__21540\,
            I => \N__21536\
        );

    \I__3273\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21533\
        );

    \I__3272\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21530\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__21533\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__21530\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3269\ : InMux
    port map (
            O => \N__21525\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__3268\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21518\
        );

    \I__3267\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21515\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__21518\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__21515\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3264\ : InMux
    port map (
            O => \N__21510\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__21507\,
            I => \N__21504\
        );

    \I__3262\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21501\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__21501\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__3260\ : InMux
    port map (
            O => \N__21498\,
            I => \N__21494\
        );

    \I__3259\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21491\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__21494\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__21491\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__3256\ : CascadeMux
    port map (
            O => \N__21486\,
            I => \VPP_VDDQ.count_2Z0Z_11_cascade_\
        );

    \I__3255\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21480\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__21480\,
            I => \VPP_VDDQ.un29_clk_100khz_1\
        );

    \I__3253\ : CascadeMux
    port map (
            O => \N__21477\,
            I => \N__21473\
        );

    \I__3252\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21470\
        );

    \I__3251\ : InMux
    port map (
            O => \N__21473\,
            I => \N__21466\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__21470\,
            I => \N__21463\
        );

    \I__3249\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21460\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__21466\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__21463\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__21460\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__21453\,
            I => \N__21450\
        );

    \I__3244\ : InMux
    port map (
            O => \N__21450\,
            I => \N__21445\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__21449\,
            I => \N__21442\
        );

    \I__3242\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21438\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__21445\,
            I => \N__21435\
        );

    \I__3240\ : InMux
    port map (
            O => \N__21442\,
            I => \N__21430\
        );

    \I__3239\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21430\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__21438\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__21435\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__21430\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3235\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21418\
        );

    \I__3234\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21415\
        );

    \I__3233\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21412\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__21418\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__21415\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__21412\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__3229\ : InMux
    port map (
            O => \N__21405\,
            I => \N__21402\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__21402\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__3227\ : InMux
    port map (
            O => \N__21399\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__3226\ : InMux
    port map (
            O => \N__21396\,
            I => \N__21393\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__21393\,
            I => \N__21388\
        );

    \I__3224\ : InMux
    port map (
            O => \N__21392\,
            I => \N__21383\
        );

    \I__3223\ : InMux
    port map (
            O => \N__21391\,
            I => \N__21383\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__21388\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__21383\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__3220\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21375\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21372\
        );

    \I__3218\ : Span4Mux_v
    port map (
            O => \N__21372\,
            I => \N__21369\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__21369\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__3216\ : InMux
    port map (
            O => \N__21366\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__3215\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21358\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__21362\,
            I => \N__21355\
        );

    \I__3213\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21352\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__21358\,
            I => \N__21349\
        );

    \I__3211\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21346\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__21352\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__21349\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__21346\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__3206\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__21333\,
            I => \N__21330\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__21330\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__3203\ : InMux
    port map (
            O => \N__21327\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__3202\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21319\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__21323\,
            I => \N__21316\
        );

    \I__3200\ : InMux
    port map (
            O => \N__21322\,
            I => \N__21313\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__21319\,
            I => \N__21310\
        );

    \I__3198\ : InMux
    port map (
            O => \N__21316\,
            I => \N__21307\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__21313\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__21310\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__21307\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3194\ : InMux
    port map (
            O => \N__21300\,
            I => \N__21297\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21294\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__21294\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__3191\ : InMux
    port map (
            O => \N__21291\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__3190\ : InMux
    port map (
            O => \N__21288\,
            I => \N__21283\
        );

    \I__3189\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21278\
        );

    \I__3188\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21278\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__21283\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__21278\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3185\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21270\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__21270\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__3183\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__21264\,
            I => \VPP_VDDQ.count_2_0_6\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__21261\,
            I => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__21258\,
            I => \N__21254\
        );

    \I__3179\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21251\
        );

    \I__3178\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21248\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__21251\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__21248\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__3175\ : CascadeMux
    port map (
            O => \N__21243\,
            I => \N__21240\
        );

    \I__3174\ : InMux
    port map (
            O => \N__21240\,
            I => \N__21237\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__21237\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__21234\,
            I => \VPP_VDDQ.count_2Z0Z_9_cascade_\
        );

    \I__3171\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21225\
        );

    \I__3170\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21225\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__21225\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__3168\ : InMux
    port map (
            O => \N__21222\,
            I => \N__21219\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__21219\,
            I => \VPP_VDDQ.un29_clk_100khz_0\
        );

    \I__3166\ : InMux
    port map (
            O => \N__21216\,
            I => \N__21213\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__21213\,
            I => \N__21210\
        );

    \I__3164\ : Span4Mux_s1_v
    port map (
            O => \N__21210\,
            I => \N__21204\
        );

    \I__3163\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21199\
        );

    \I__3162\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21199\
        );

    \I__3161\ : InMux
    port map (
            O => \N__21207\,
            I => \N__21196\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__21204\,
            I => \POWERLED.un1_dutycycle_53_44_d_1_0_tz\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__21199\,
            I => \POWERLED.un1_dutycycle_53_44_d_1_0_tz\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__21196\,
            I => \POWERLED.un1_dutycycle_53_44_d_1_0_tz\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__21189\,
            I => \POWERLED.dutycycle_er_RNIZ0Z_9_cascade_\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__21186\,
            I => \N__21182\
        );

    \I__3155\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21179\
        );

    \I__3154\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21176\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21173\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__21176\,
            I => \N__21170\
        );

    \I__3151\ : Span4Mux_h
    port map (
            O => \N__21173\,
            I => \N__21167\
        );

    \I__3150\ : Odrv4
    port map (
            O => \N__21170\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_4\
        );

    \I__3149\ : Odrv4
    port map (
            O => \N__21167\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_4\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__21162\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_4_cascade_\
        );

    \I__3147\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__21156\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_10\
        );

    \I__3145\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__21150\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_10\
        );

    \I__3143\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__21144\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__21141\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_10_cascade_\
        );

    \I__3140\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21135\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__21135\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__3138\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21126\
        );

    \I__3137\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21126\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__21126\,
            I => \N__21123\
        );

    \I__3135\ : Span4Mux_s1_v
    port map (
            O => \N__21123\,
            I => \N__21120\
        );

    \I__3134\ : Span4Mux_v
    port map (
            O => \N__21120\,
            I => \N__21117\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__21117\,
            I => \N__21114\
        );

    \I__3132\ : Odrv4
    port map (
            O => \N__21114\,
            I => \VPP_VDDQ.N_297_0\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__21111\,
            I => \N__21107\
        );

    \I__3130\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21102\
        );

    \I__3129\ : InMux
    port map (
            O => \N__21107\,
            I => \N__21102\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__21102\,
            I => \N__21099\
        );

    \I__3127\ : Odrv4
    port map (
            O => \N__21099\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__21096\,
            I => \VPP_VDDQ_delayed_vddq_ok_cascade_\
        );

    \I__3125\ : IoInMux
    port map (
            O => \N__21093\,
            I => \N__21090\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__21090\,
            I => vccst_pwrgd
        );

    \I__3123\ : IoInMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__21084\,
            I => \N__21081\
        );

    \I__3121\ : Span4Mux_s2_h
    port map (
            O => \N__21081\,
            I => \N__21077\
        );

    \I__3120\ : IoInMux
    port map (
            O => \N__21080\,
            I => \N__21074\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__21077\,
            I => \N__21071\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__21074\,
            I => \N__21068\
        );

    \I__3117\ : Sp12to4
    port map (
            O => \N__21071\,
            I => \N__21065\
        );

    \I__3116\ : IoSpan4Mux
    port map (
            O => \N__21068\,
            I => \N__21062\
        );

    \I__3115\ : Span12Mux_v
    port map (
            O => \N__21065\,
            I => \N__21059\
        );

    \I__3114\ : IoSpan4Mux
    port map (
            O => \N__21062\,
            I => \N__21056\
        );

    \I__3113\ : Odrv12
    port map (
            O => \N__21059\,
            I => pch_pwrok
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__21056\,
            I => pch_pwrok
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__21051\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__21048\,
            I => \N__21045\
        );

    \I__3109\ : InMux
    port map (
            O => \N__21045\,
            I => \N__21042\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__21042\,
            I => \POWERLED.un1_dutycycle_53_axb_7_1\
        );

    \I__3107\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__21036\,
            I => \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_1\
        );

    \I__3105\ : InMux
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__21030\,
            I => \POWERLED.un1_dutycycle_53_44_d_c_1_s_1\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__21027\,
            I => \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_2_cascade_\
        );

    \I__3102\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21021\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__21021\,
            I => \N__21018\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__21018\,
            I => \N__21015\
        );

    \I__3099\ : Odrv4
    port map (
            O => \N__21015\,
            I => \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_0\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__21012\,
            I => \N__21009\
        );

    \I__3097\ : InMux
    port map (
            O => \N__21009\,
            I => \N__21003\
        );

    \I__3096\ : InMux
    port map (
            O => \N__21008\,
            I => \N__21003\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__20999\
        );

    \I__3094\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20996\
        );

    \I__3093\ : Span4Mux_v
    port map (
            O => \N__20999\,
            I => \N__20993\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__20996\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__20993\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31\
        );

    \I__3090\ : InMux
    port map (
            O => \N__20988\,
            I => \POWERLED.un1_dutycycle_94_cry_8_cZ0\
        );

    \I__3089\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20979\
        );

    \I__3088\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20979\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__20979\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\
        );

    \I__3086\ : InMux
    port map (
            O => \N__20976\,
            I => \POWERLED.un1_dutycycle_94_cry_9_cZ0\
        );

    \I__3085\ : InMux
    port map (
            O => \N__20973\,
            I => \POWERLED.un1_dutycycle_94_cry_10\
        );

    \I__3084\ : InMux
    port map (
            O => \N__20970\,
            I => \POWERLED.un1_dutycycle_94_cry_11_cZ0\
        );

    \I__3083\ : InMux
    port map (
            O => \N__20967\,
            I => \POWERLED.un1_dutycycle_94_cry_12\
        );

    \I__3082\ : InMux
    port map (
            O => \N__20964\,
            I => \POWERLED.un1_dutycycle_94_cry_13\
        );

    \I__3081\ : InMux
    port map (
            O => \N__20961\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__3080\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20954\
        );

    \I__3079\ : InMux
    port map (
            O => \N__20957\,
            I => \N__20951\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__20954\,
            I => \N__20948\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__20951\,
            I => \N__20945\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__20948\,
            I => \N__20940\
        );

    \I__3075\ : Span4Mux_h
    port map (
            O => \N__20945\,
            I => \N__20940\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__20940\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__20937\,
            I => \POWERLED.un1_dutycycle_53_axb_7_cascade_\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20931\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__20931\,
            I => \N__20928\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__20928\,
            I => \N__20925\
        );

    \I__3069\ : Span4Mux_h
    port map (
            O => \N__20925\,
            I => \N__20922\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__20922\,
            I => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\
        );

    \I__3067\ : InMux
    port map (
            O => \N__20919\,
            I => \POWERLED.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__3066\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20913\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__20913\,
            I => \N__20910\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__20910\,
            I => \N__20907\
        );

    \I__3063\ : Span4Mux_h
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__20904\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNIZ0\
        );

    \I__3061\ : InMux
    port map (
            O => \N__20901\,
            I => \POWERLED.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__3059\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20889\
        );

    \I__3058\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20889\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__20889\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__3056\ : InMux
    port map (
            O => \N__20886\,
            I => \POWERLED.un1_dutycycle_94_cry_2\
        );

    \I__3055\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20879\
        );

    \I__3054\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20876\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__20879\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__20876\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__3051\ : InMux
    port map (
            O => \N__20871\,
            I => \POWERLED.un1_dutycycle_94_cry_3_cZ0\
        );

    \I__3050\ : InMux
    port map (
            O => \N__20868\,
            I => \N__20865\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20862\
        );

    \I__3048\ : Odrv12
    port map (
            O => \N__20862\,
            I => \POWERLED.N_308\
        );

    \I__3047\ : InMux
    port map (
            O => \N__20859\,
            I => \POWERLED.un1_dutycycle_94_cry_4\
        );

    \I__3046\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20853\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__3044\ : Span4Mux_h
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__20847\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\
        );

    \I__3042\ : InMux
    port map (
            O => \N__20844\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3041\ : InMux
    port map (
            O => \N__20841\,
            I => \POWERLED.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__20838\,
            I => \N__20834\
        );

    \I__3039\ : InMux
    port map (
            O => \N__20837\,
            I => \N__20829\
        );

    \I__3038\ : InMux
    port map (
            O => \N__20834\,
            I => \N__20829\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__20829\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\
        );

    \I__3036\ : InMux
    port map (
            O => \N__20826\,
            I => \bfn_5_14_0_\
        );

    \I__3035\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20817\
        );

    \I__3034\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20817\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__20817\,
            I => \POWERLED.func_state_RNI_1Z0Z_0\
        );

    \I__3032\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__20811\,
            I => \POWERLED.N_321\
        );

    \I__3030\ : InMux
    port map (
            O => \N__20808\,
            I => \N__20805\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__20805\,
            I => \POWERLED.un1_clk_100khz_43_and_i_0_d_0\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \POWERLED.un1_clk_100khz_40_and_i_0_0_0_cascade_\
        );

    \I__3027\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__20796\,
            I => \POWERLED.dutycycle_en_8\
        );

    \I__3025\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20787\
        );

    \I__3024\ : InMux
    port map (
            O => \N__20792\,
            I => \N__20787\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__20787\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__20784\,
            I => \POWERLED.dutycycle_en_8_cascade_\
        );

    \I__3021\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__20778\,
            I => \POWERLED.un1_clk_100khz_40_and_i_0_0_0\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__20775\,
            I => \POWERLED.un1_clk_100khz_40_and_i_0_d_0_cascade_\
        );

    \I__3018\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20769\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__20769\,
            I => \N__20766\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__20766\,
            I => \POWERLED.dutycycle_en_6\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__20763\,
            I => \POWERLED.dutycycle_en_6_cascade_\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__20760\,
            I => \N__20757\
        );

    \I__3013\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20754\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__20754\,
            I => \N__20750\
        );

    \I__3011\ : InMux
    port map (
            O => \N__20753\,
            I => \N__20747\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__20750\,
            I => \N__20744\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__20747\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__20744\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__20739\,
            I => \N__20736\
        );

    \I__3006\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20733\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__20733\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__3004\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__20727\,
            I => \POWERLED.N_388_N\
        );

    \I__3002\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20721\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__20721\,
            I => \N__20718\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__20715\,
            I => \POWERLED.un1_func_state25_6_0_1\
        );

    \I__2998\ : InMux
    port map (
            O => \N__20712\,
            I => \N__20709\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__20709\,
            I => \POWERLED.un1_func_state25_4_i_a2_1\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__20706\,
            I => \N__20703\
        );

    \I__2995\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20700\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__20700\,
            I => \POWERLED.un1_func_state25_6_0_1_1\
        );

    \I__2993\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__20694\,
            I => \POWERLED.N_425\
        );

    \I__2991\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__20685\,
            I => \POWERLED.count_clk_RNI0TA81Z0Z_7\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__20682\,
            I => \POWERLED.count_clk_RNI0TA81Z0Z_7_cascade_\
        );

    \I__2987\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20651\
        );

    \I__2986\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20651\
        );

    \I__2985\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20651\
        );

    \I__2984\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20651\
        );

    \I__2983\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20644\
        );

    \I__2982\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20644\
        );

    \I__2981\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20644\
        );

    \I__2980\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20639\
        );

    \I__2979\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20639\
        );

    \I__2978\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20632\
        );

    \I__2977\ : InMux
    port map (
            O => \N__20669\,
            I => \N__20632\
        );

    \I__2976\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20632\
        );

    \I__2975\ : InMux
    port map (
            O => \N__20667\,
            I => \N__20627\
        );

    \I__2974\ : InMux
    port map (
            O => \N__20666\,
            I => \N__20627\
        );

    \I__2973\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20614\
        );

    \I__2972\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20614\
        );

    \I__2971\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20614\
        );

    \I__2970\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20614\
        );

    \I__2969\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20614\
        );

    \I__2968\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20614\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__20651\,
            I => \N__20605\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20605\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__20639\,
            I => \N__20605\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__20632\,
            I => \N__20605\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20600\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__20614\,
            I => \N__20600\
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__20605\,
            I => \POWERLED.N_128\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__20600\,
            I => \POWERLED.N_128\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__20595\,
            I => \POWERLED.N_431_cascade_\
        );

    \I__2958\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20581\
        );

    \I__2957\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20576\
        );

    \I__2956\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20576\
        );

    \I__2955\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20569\
        );

    \I__2954\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20569\
        );

    \I__2953\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20569\
        );

    \I__2952\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20566\
        );

    \I__2951\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20562\
        );

    \I__2950\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20559\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20552\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__20576\,
            I => \N__20552\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__20569\,
            I => \N__20552\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20549\
        );

    \I__2945\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20546\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20541\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__20559\,
            I => \N__20541\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__20552\,
            I => \N__20538\
        );

    \I__2941\ : Odrv12
    port map (
            O => \N__20549\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__20546\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2939\ : Odrv4
    port map (
            O => \N__20541\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__20538\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__2937\ : InMux
    port map (
            O => \N__20529\,
            I => \N__20526\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__20526\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__2935\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__20520\,
            I => \N__20512\
        );

    \I__2933\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20505\
        );

    \I__2932\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20496\
        );

    \I__2931\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20496\
        );

    \I__2930\ : InMux
    port map (
            O => \N__20516\,
            I => \N__20496\
        );

    \I__2929\ : InMux
    port map (
            O => \N__20515\,
            I => \N__20496\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__20512\,
            I => \N__20490\
        );

    \I__2927\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20480\
        );

    \I__2926\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20480\
        );

    \I__2925\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20480\
        );

    \I__2924\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20480\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20475\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__20496\,
            I => \N__20475\
        );

    \I__2921\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20468\
        );

    \I__2920\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20468\
        );

    \I__2919\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20468\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__20490\,
            I => \N__20463\
        );

    \I__2917\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20460\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__20480\,
            I => \N__20457\
        );

    \I__2915\ : Span4Mux_s1_h
    port map (
            O => \N__20475\,
            I => \N__20452\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__20468\,
            I => \N__20452\
        );

    \I__2913\ : InMux
    port map (
            O => \N__20467\,
            I => \N__20447\
        );

    \I__2912\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20447\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__20463\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__20460\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__20457\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__20452\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__20447\,
            I => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\
        );

    \I__2906\ : SRMux
    port map (
            O => \N__20436\,
            I => \N__20427\
        );

    \I__2905\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20422\
        );

    \I__2904\ : SRMux
    port map (
            O => \N__20434\,
            I => \N__20422\
        );

    \I__2903\ : InMux
    port map (
            O => \N__20433\,
            I => \N__20417\
        );

    \I__2902\ : SRMux
    port map (
            O => \N__20432\,
            I => \N__20417\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__20431\,
            I => \N__20414\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__20430\,
            I => \N__20411\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__20427\,
            I => \N__20401\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__20422\,
            I => \N__20396\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__20417\,
            I => \N__20396\
        );

    \I__2896\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20385\
        );

    \I__2895\ : InMux
    port map (
            O => \N__20411\,
            I => \N__20385\
        );

    \I__2894\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20385\
        );

    \I__2893\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20385\
        );

    \I__2892\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20385\
        );

    \I__2891\ : SRMux
    port map (
            O => \N__20407\,
            I => \N__20370\
        );

    \I__2890\ : SRMux
    port map (
            O => \N__20406\,
            I => \N__20367\
        );

    \I__2889\ : SRMux
    port map (
            O => \N__20405\,
            I => \N__20364\
        );

    \I__2888\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20361\
        );

    \I__2887\ : Span4Mux_v
    port map (
            O => \N__20401\,
            I => \N__20349\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__20396\,
            I => \N__20349\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__20385\,
            I => \N__20349\
        );

    \I__2884\ : InMux
    port map (
            O => \N__20384\,
            I => \N__20344\
        );

    \I__2883\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20344\
        );

    \I__2882\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20339\
        );

    \I__2881\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20339\
        );

    \I__2880\ : InMux
    port map (
            O => \N__20380\,
            I => \N__20332\
        );

    \I__2879\ : InMux
    port map (
            O => \N__20379\,
            I => \N__20332\
        );

    \I__2878\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20332\
        );

    \I__2877\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20327\
        );

    \I__2876\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20327\
        );

    \I__2875\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20324\
        );

    \I__2874\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20321\
        );

    \I__2873\ : SRMux
    port map (
            O => \N__20373\,
            I => \N__20318\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__20370\,
            I => \N__20315\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__20367\,
            I => \N__20312\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__20364\,
            I => \N__20307\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__20361\,
            I => \N__20307\
        );

    \I__2868\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20300\
        );

    \I__2867\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20300\
        );

    \I__2866\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20300\
        );

    \I__2865\ : InMux
    port map (
            O => \N__20357\,
            I => \N__20295\
        );

    \I__2864\ : InMux
    port map (
            O => \N__20356\,
            I => \N__20295\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__20349\,
            I => \N__20288\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__20344\,
            I => \N__20288\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__20339\,
            I => \N__20288\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__20332\,
            I => \N__20281\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__20327\,
            I => \N__20281\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__20324\,
            I => \N__20281\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__20321\,
            I => \N__20278\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__20318\,
            I => \N__20275\
        );

    \I__2855\ : Span4Mux_h
    port map (
            O => \N__20315\,
            I => \N__20270\
        );

    \I__2854\ : Span4Mux_h
    port map (
            O => \N__20312\,
            I => \N__20270\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__20307\,
            I => \N__20263\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__20300\,
            I => \N__20263\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20263\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__20288\,
            I => \N__20256\
        );

    \I__2849\ : Span4Mux_v
    port map (
            O => \N__20281\,
            I => \N__20256\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__20278\,
            I => \N__20256\
        );

    \I__2847\ : Odrv12
    port map (
            O => \N__20275\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__20270\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__20263\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__20256\,
            I => \RSMRST_PWRGD.count_0_sqmuxa\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__20247\,
            I => \N__20243\
        );

    \I__2842\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20240\
        );

    \I__2841\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20237\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__20240\,
            I => \N__20234\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__20237\,
            I => \N__20228\
        );

    \I__2838\ : Span12Mux_s8_v
    port map (
            O => \N__20234\,
            I => \N__20225\
        );

    \I__2837\ : InMux
    port map (
            O => \N__20233\,
            I => \N__20218\
        );

    \I__2836\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20218\
        );

    \I__2835\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20218\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__20228\,
            I => \N__20215\
        );

    \I__2833\ : Odrv12
    port map (
            O => \N__20225\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__20218\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__20215\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__2830\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20205\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__20205\,
            I => \N__20202\
        );

    \I__2828\ : Span4Mux_v
    port map (
            O => \N__20202\,
            I => \N__20199\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__20199\,
            I => \RSMRST_PWRGD.count_rst_5\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__2825\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__20190\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \POWERLED.count_clkZ0Z_13_cascade_\
        );

    \I__2822\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__20181\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__20178\,
            I => \POWERLED.un34_clk_100khz_9_cascade_\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__20175\,
            I => \N__20171\
        );

    \I__2818\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20168\
        );

    \I__2817\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20165\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__20168\,
            I => \N__20162\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__20165\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__20162\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__2813\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20154\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__20154\,
            I => \POWERLED.un34_clk_100khz_8\
        );

    \I__2811\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20148\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__20148\,
            I => \POWERLED.count_off_0_5\
        );

    \I__2809\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20141\
        );

    \I__2808\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20138\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__20141\,
            I => \N__20135\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__20138\,
            I => \POWERLED.count_off_1_5\
        );

    \I__2805\ : Odrv4
    port map (
            O => \N__20135\,
            I => \POWERLED.count_off_1_5\
        );

    \I__2804\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20126\
        );

    \I__2803\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20123\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__20126\,
            I => \N__20120\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__20123\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__20120\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__20115\,
            I => \N__20111\
        );

    \I__2798\ : InMux
    port map (
            O => \N__20114\,
            I => \N__20106\
        );

    \I__2797\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20106\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__20106\,
            I => \N__20103\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__20103\,
            I => \POWERLED.count_off_1_2\
        );

    \I__2794\ : InMux
    port map (
            O => \N__20100\,
            I => \N__20097\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__20097\,
            I => \POWERLED.count_off_0_2\
        );

    \I__2792\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20091\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__20091\,
            I => \POWERLED.count_off_0_4\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__20088\,
            I => \N__20085\
        );

    \I__2789\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20079\
        );

    \I__2788\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20079\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__20079\,
            I => \N__20076\
        );

    \I__2786\ : Odrv12
    port map (
            O => \N__20076\,
            I => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__20073\,
            I => \N__20070\
        );

    \I__2784\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20066\
        );

    \I__2783\ : InMux
    port map (
            O => \N__20069\,
            I => \N__20063\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__20066\,
            I => \N__20060\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__20063\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__20060\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__2779\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__20052\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__20049\,
            I => \N__20046\
        );

    \I__2776\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20043\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__20043\,
            I => \POWERLED.count_clk_0_10\
        );

    \I__2774\ : InMux
    port map (
            O => \N__20040\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__2773\ : InMux
    port map (
            O => \N__20037\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__2772\ : InMux
    port map (
            O => \N__20034\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__2771\ : InMux
    port map (
            O => \N__20031\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__2770\ : InMux
    port map (
            O => \N__20028\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__2769\ : InMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__20019\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__20016\,
            I => \N__20013\
        );

    \I__2765\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__20010\,
            I => \N__20005\
        );

    \I__2763\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20002\
        );

    \I__2762\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19999\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__20005\,
            I => \N__19996\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__20002\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__19999\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__19996\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__19989\,
            I => \POWERLED.count_offZ0Z_2_cascade_\
        );

    \I__2756\ : InMux
    port map (
            O => \N__19986\,
            I => \POWERLED.un3_count_off_1_cry_1\
        );

    \I__2755\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19977\
        );

    \I__2754\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19977\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__19977\,
            I => \N__19974\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__19974\,
            I => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\
        );

    \I__2751\ : InMux
    port map (
            O => \N__19971\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__2750\ : InMux
    port map (
            O => \N__19968\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__2749\ : InMux
    port map (
            O => \N__19965\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__2748\ : InMux
    port map (
            O => \N__19962\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__2747\ : InMux
    port map (
            O => \N__19959\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__2746\ : InMux
    port map (
            O => \N__19956\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__2745\ : InMux
    port map (
            O => \N__19953\,
            I => \bfn_5_7_0_\
        );

    \I__2744\ : InMux
    port map (
            O => \N__19950\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__19947\,
            I => \N__19944\
        );

    \I__2742\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19941\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__19941\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__2739\ : InMux
    port map (
            O => \N__19935\,
            I => \N__19932\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__19932\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__19929\,
            I => \N__19926\
        );

    \I__2736\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__19923\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__2734\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19915\
        );

    \I__2733\ : InMux
    port map (
            O => \N__19919\,
            I => \N__19912\
        );

    \I__2732\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19909\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19899\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__19912\,
            I => \N__19899\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__19909\,
            I => \N__19899\
        );

    \I__2728\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19896\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__19907\,
            I => \N__19893\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19889\
        );

    \I__2725\ : Span4Mux_v
    port map (
            O => \N__19899\,
            I => \N__19878\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__19896\,
            I => \N__19878\
        );

    \I__2723\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19873\
        );

    \I__2722\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19873\
        );

    \I__2721\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19868\
        );

    \I__2720\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19868\
        );

    \I__2719\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19857\
        );

    \I__2718\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19857\
        );

    \I__2717\ : InMux
    port map (
            O => \N__19885\,
            I => \N__19857\
        );

    \I__2716\ : InMux
    port map (
            O => \N__19884\,
            I => \N__19857\
        );

    \I__2715\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19857\
        );

    \I__2714\ : Span4Mux_v
    port map (
            O => \N__19878\,
            I => \N__19854\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__19873\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__19868\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__19857\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__19854\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__2709\ : IoInMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__2707\ : Span4Mux_s0_h
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__2706\ : Span4Mux_h
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__19833\,
            I => \N__19830\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__19830\,
            I => hda_sdo_atp
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__19827\,
            I => \HDA_STRAP.curr_stateZ0Z_1_cascade_\
        );

    \I__2702\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__19821\,
            I => \HDA_STRAP.curr_state_3_1\
        );

    \I__2700\ : InMux
    port map (
            O => \N__19818\,
            I => \N__19806\
        );

    \I__2699\ : InMux
    port map (
            O => \N__19817\,
            I => \N__19806\
        );

    \I__2698\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19806\
        );

    \I__2697\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19806\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__19806\,
            I => \HDA_STRAP.N_208\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__19803\,
            I => \N__19799\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__19802\,
            I => \N__19796\
        );

    \I__2693\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19792\
        );

    \I__2692\ : InMux
    port map (
            O => \N__19796\,
            I => \N__19787\
        );

    \I__2691\ : InMux
    port map (
            O => \N__19795\,
            I => \N__19787\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__19792\,
            I => \HDA_STRAP.curr_state_i_2\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__19787\,
            I => \HDA_STRAP.curr_state_i_2\
        );

    \I__2688\ : InMux
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__19779\,
            I => \HDA_STRAP.HDA_SDO_ATP_0\
        );

    \I__2686\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19773\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__19773\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__2683\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19764\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__19764\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__2680\ : InMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__19755\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__2678\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19748\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__19751\,
            I => \N__19745\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__19748\,
            I => \N__19736\
        );

    \I__2675\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19733\
        );

    \I__2674\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19730\
        );

    \I__2673\ : InMux
    port map (
            O => \N__19743\,
            I => \N__19719\
        );

    \I__2672\ : InMux
    port map (
            O => \N__19742\,
            I => \N__19719\
        );

    \I__2671\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19719\
        );

    \I__2670\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19719\
        );

    \I__2669\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19719\
        );

    \I__2668\ : Span4Mux_s3_v
    port map (
            O => \N__19736\,
            I => \N__19716\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__19733\,
            I => \N__19713\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19710\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__19719\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__19716\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__19713\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__19710\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__19701\,
            I => \N_392_cascade_\
        );

    \I__2660\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19693\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__19697\,
            I => \N__19686\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__19696\,
            I => \N__19683\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__19693\,
            I => \N__19679\
        );

    \I__2656\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19676\
        );

    \I__2655\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19673\
        );

    \I__2654\ : InMux
    port map (
            O => \N__19690\,
            I => \N__19662\
        );

    \I__2653\ : InMux
    port map (
            O => \N__19689\,
            I => \N__19662\
        );

    \I__2652\ : InMux
    port map (
            O => \N__19686\,
            I => \N__19662\
        );

    \I__2651\ : InMux
    port map (
            O => \N__19683\,
            I => \N__19662\
        );

    \I__2650\ : InMux
    port map (
            O => \N__19682\,
            I => \N__19662\
        );

    \I__2649\ : Span4Mux_s3_v
    port map (
            O => \N__19679\,
            I => \N__19659\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__19676\,
            I => \N__19656\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__19673\,
            I => \N__19653\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__19662\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2645\ : Odrv4
    port map (
            O => \N__19659\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2644\ : Odrv12
    port map (
            O => \N__19656\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__19653\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__2642\ : CascadeMux
    port map (
            O => \N__19644\,
            I => \N__19640\
        );

    \I__2641\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19634\
        );

    \I__2640\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19625\
        );

    \I__2639\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19625\
        );

    \I__2638\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19625\
        );

    \I__2637\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19625\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19622\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19619\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__19622\,
            I => \N__19616\
        );

    \I__2633\ : Span4Mux_s2_h
    port map (
            O => \N__19619\,
            I => \N__19613\
        );

    \I__2632\ : Sp12to4
    port map (
            O => \N__19616\,
            I => \N__19610\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__19613\,
            I => \N__19607\
        );

    \I__2630\ : Span12Mux_v
    port map (
            O => \N__19610\,
            I => \N__19604\
        );

    \I__2629\ : Span4Mux_v
    port map (
            O => \N__19607\,
            I => \N__19601\
        );

    \I__2628\ : Odrv12
    port map (
            O => \N__19604\,
            I => \RSMRSTn_0\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__19601\,
            I => \RSMRSTn_0\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__19596\,
            I => \VPP_VDDQ.count_2Z0Z_13_cascade_\
        );

    \I__2625\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__19590\,
            I => \VPP_VDDQ.un29_clk_100khz_2\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__19587\,
            I => \VPP_VDDQ.un29_clk_100khz_3_cascade_\
        );

    \I__2622\ : InMux
    port map (
            O => \N__19584\,
            I => \N__19578\
        );

    \I__2621\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19578\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__19578\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__19575\,
            I => \HDA_STRAP.i4_mux_cascade_\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__19572\,
            I => \HDA_STRAP.curr_state_i_2_cascade_\
        );

    \I__2617\ : InMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__19566\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__2615\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__19560\,
            I => \POWERLED.un1_dutycycle_53_39_c_1\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__19557\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_\
        );

    \I__2612\ : CascadeMux
    port map (
            O => \N__19554\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_10_cascade_\
        );

    \I__2611\ : IoInMux
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__19548\,
            I => \N__19544\
        );

    \I__2609\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19541\
        );

    \I__2608\ : Span4Mux_s2_h
    port map (
            O => \N__19544\,
            I => \N__19538\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__19541\,
            I => \N__19535\
        );

    \I__2606\ : Sp12to4
    port map (
            O => \N__19538\,
            I => \N__19532\
        );

    \I__2605\ : Sp12to4
    port map (
            O => \N__19535\,
            I => \N__19529\
        );

    \I__2604\ : Span12Mux_s11_v
    port map (
            O => \N__19532\,
            I => \N__19526\
        );

    \I__2603\ : Span12Mux_s11_v
    port map (
            O => \N__19529\,
            I => \N__19523\
        );

    \I__2602\ : Odrv12
    port map (
            O => \N__19526\,
            I => v1p8a_ok
        );

    \I__2601\ : Odrv12
    port map (
            O => \N__19523\,
            I => v1p8a_ok
        );

    \I__2600\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19515\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__2597\ : Span4Mux_h
    port map (
            O => \N__19509\,
            I => \N__19506\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__19506\,
            I => v5a_ok
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \POWERLED.dutycycleZ0Z_2_cascade_\
        );

    \I__2594\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19497\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__19497\,
            I => \POWERLED.dutycycle_RNIANIR7Z0Z_10\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__19494\,
            I => \N__19491\
        );

    \I__2591\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19485\
        );

    \I__2590\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19485\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__19485\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__2588\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19476\
        );

    \I__2587\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19476\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19473\
        );

    \I__2585\ : Span4Mux_s3_v
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__19470\,
            I => \POWERLED.dutycycle_eena_3_d_0\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__19467\,
            I => \N__19463\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__19466\,
            I => \N__19460\
        );

    \I__2581\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19455\
        );

    \I__2580\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19455\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__19455\,
            I => \N__19452\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__19452\,
            I => \N__19449\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__19446\,
            I => \POWERLED.dutycycle_eena_3_0_0\
        );

    \I__2575\ : InMux
    port map (
            O => \N__19443\,
            I => \N__19440\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__19440\,
            I => \POWERLED.dutycycle_RNIANIR7Z0Z_8\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \POWERLED.dutycycle_RNIANIR7Z0Z_8_cascade_\
        );

    \I__2572\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19430\
        );

    \I__2571\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19427\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__19430\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__19427\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__2568\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19419\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__19419\,
            I => \N__19416\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__19413\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_3\
        );

    \I__2564\ : InMux
    port map (
            O => \N__19410\,
            I => \N__19406\
        );

    \I__2563\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19403\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__19406\,
            I => \N__19400\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19397\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__19400\,
            I => \POWERLED.func_state_RNI8H551_0Z0Z_0\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__19397\,
            I => \POWERLED.func_state_RNI8H551_0Z0Z_0\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__19392\,
            I => \N__19387\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__19391\,
            I => \N__19384\
        );

    \I__2556\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19380\
        );

    \I__2555\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19375\
        );

    \I__2554\ : InMux
    port map (
            O => \N__19384\,
            I => \N__19375\
        );

    \I__2553\ : InMux
    port map (
            O => \N__19383\,
            I => \N__19372\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__19380\,
            I => \N__19369\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__19375\,
            I => \N__19363\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__19372\,
            I => \N__19363\
        );

    \I__2549\ : Span4Mux_s2_v
    port map (
            O => \N__19369\,
            I => \N__19360\
        );

    \I__2548\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19357\
        );

    \I__2547\ : Span4Mux_v
    port map (
            O => \N__19363\,
            I => \N__19354\
        );

    \I__2546\ : Odrv4
    port map (
            O => \N__19360\,
            I => \POWERLED.N_372\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__19357\,
            I => \POWERLED.N_372\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__19354\,
            I => \POWERLED.N_372\
        );

    \I__2543\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__19344\,
            I => \N__19339\
        );

    \I__2541\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19334\
        );

    \I__2540\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19334\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__19339\,
            I => \N__19331\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__19334\,
            I => \POWERLED.func_state_RNIZ0Z_0\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__19331\,
            I => \POWERLED.func_state_RNIZ0Z_0\
        );

    \I__2536\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19323\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__19317\,
            I => \POWERLED.un1_clk_100khz_36_and_i_a2_6_0_0_0\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__19314\,
            I => \POWERLED.un1_dutycycle_53_7_a0_1_a1_0_cascade_\
        );

    \I__2531\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19308\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__19308\,
            I => \N__19305\
        );

    \I__2529\ : Span4Mux_h
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__19302\,
            I => \POWERLED.un1_dutycycle_53_7_a0_2\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__19299\,
            I => \POWERLED.un1_dutycycle_53_axb_13_1_0_cascade_\
        );

    \I__2526\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19293\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__19293\,
            I => \POWERLED.un1_dutycycle_53_7_a0_3\
        );

    \I__2524\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19287\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__19287\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_12\
        );

    \I__2522\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__19281\,
            I => \POWERLED.func_state_RNI8H551Z0Z_0\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__19278\,
            I => \POWERLED.dutycycle_RNIANIR7Z0Z_10_cascade_\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__19275\,
            I => \POWERLED.dutycycleZ0Z_6_cascade_\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__19272\,
            I => \N__19269\
        );

    \I__2517\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19257\
        );

    \I__2516\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19257\
        );

    \I__2515\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19257\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__19266\,
            I => \N__19254\
        );

    \I__2513\ : InMux
    port map (
            O => \N__19265\,
            I => \N__19250\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__19264\,
            I => \N__19247\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19240\
        );

    \I__2510\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19237\
        );

    \I__2509\ : InMux
    port map (
            O => \N__19253\,
            I => \N__19234\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__19250\,
            I => \N__19229\
        );

    \I__2507\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19222\
        );

    \I__2506\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19222\
        );

    \I__2505\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19222\
        );

    \I__2504\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19217\
        );

    \I__2503\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19217\
        );

    \I__2502\ : Span4Mux_s3_h
    port map (
            O => \N__19240\,
            I => \N__19209\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__19237\,
            I => \N__19209\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__19234\,
            I => \N__19209\
        );

    \I__2499\ : InMux
    port map (
            O => \N__19233\,
            I => \N__19204\
        );

    \I__2498\ : InMux
    port map (
            O => \N__19232\,
            I => \N__19204\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__19229\,
            I => \N__19199\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__19222\,
            I => \N__19199\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__19217\,
            I => \N__19196\
        );

    \I__2494\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19193\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__19209\,
            I => \N__19180\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__19204\,
            I => \N__19180\
        );

    \I__2491\ : Span4Mux_v
    port map (
            O => \N__19199\,
            I => \N__19173\
        );

    \I__2490\ : Span4Mux_v
    port map (
            O => \N__19196\,
            I => \N__19173\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__19193\,
            I => \N__19173\
        );

    \I__2488\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19160\
        );

    \I__2487\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19160\
        );

    \I__2486\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19160\
        );

    \I__2485\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19160\
        );

    \I__2484\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19160\
        );

    \I__2483\ : InMux
    port map (
            O => \N__19187\,
            I => \N__19160\
        );

    \I__2482\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19155\
        );

    \I__2481\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19155\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__19180\,
            I => \N__19152\
        );

    \I__2479\ : IoSpan4Mux
    port map (
            O => \N__19173\,
            I => \N__19149\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__19160\,
            I => \N__19144\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19144\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__19152\,
            I => slp_s4n
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__19149\,
            I => slp_s4n
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__19144\,
            I => slp_s4n
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__19137\,
            I => \N__19134\
        );

    \I__2472\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19121\
        );

    \I__2471\ : InMux
    port map (
            O => \N__19133\,
            I => \N__19121\
        );

    \I__2470\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19121\
        );

    \I__2469\ : InMux
    port map (
            O => \N__19131\,
            I => \N__19114\
        );

    \I__2468\ : InMux
    port map (
            O => \N__19130\,
            I => \N__19114\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__19129\,
            I => \N__19110\
        );

    \I__2466\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19106\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19103\
        );

    \I__2464\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19098\
        );

    \I__2463\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19098\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19094\
        );

    \I__2461\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19089\
        );

    \I__2460\ : InMux
    port map (
            O => \N__19110\,
            I => \N__19089\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__19109\,
            I => \N__19086\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__19106\,
            I => \N__19078\
        );

    \I__2457\ : Span4Mux_v
    port map (
            O => \N__19103\,
            I => \N__19073\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__19098\,
            I => \N__19073\
        );

    \I__2455\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19070\
        );

    \I__2454\ : Span4Mux_v
    port map (
            O => \N__19094\,
            I => \N__19065\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__19089\,
            I => \N__19065\
        );

    \I__2452\ : InMux
    port map (
            O => \N__19086\,
            I => \N__19062\
        );

    \I__2451\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19051\
        );

    \I__2450\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19051\
        );

    \I__2449\ : InMux
    port map (
            O => \N__19083\,
            I => \N__19051\
        );

    \I__2448\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19051\
        );

    \I__2447\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19051\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__19078\,
            I => \N__19045\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__19073\,
            I => \N__19045\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__19070\,
            I => \N__19042\
        );

    \I__2443\ : Span4Mux_s2_h
    port map (
            O => \N__19065\,
            I => \N__19035\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__19062\,
            I => \N__19035\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__19051\,
            I => \N__19035\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__19050\,
            I => \N__19031\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__19045\,
            I => \N__19026\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__19042\,
            I => \N__19026\
        );

    \I__2437\ : Span4Mux_h
    port map (
            O => \N__19035\,
            I => \N__19023\
        );

    \I__2436\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19018\
        );

    \I__2435\ : InMux
    port map (
            O => \N__19031\,
            I => \N__19018\
        );

    \I__2434\ : Span4Mux_h
    port map (
            O => \N__19026\,
            I => \N__19015\
        );

    \I__2433\ : Span4Mux_h
    port map (
            O => \N__19023\,
            I => \N__19012\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__19018\,
            I => \N__19009\
        );

    \I__2431\ : IoSpan4Mux
    port map (
            O => \N__19015\,
            I => \N__19006\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__19012\,
            I => \N__19003\
        );

    \I__2429\ : Span12Mux_s10_h
    port map (
            O => \N__19009\,
            I => \N__19000\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__19006\,
            I => slp_s3n
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__19003\,
            I => slp_s3n
        );

    \I__2426\ : Odrv12
    port map (
            O => \N__19000\,
            I => slp_s3n
        );

    \I__2425\ : InMux
    port map (
            O => \N__18993\,
            I => \N__18989\
        );

    \I__2424\ : InMux
    port map (
            O => \N__18992\,
            I => \N__18986\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__18989\,
            I => \POWERLED.un1_clk_100khz_42_and_i_o2_1_1\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__18986\,
            I => \POWERLED.un1_clk_100khz_42_and_i_o2_1_1\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__18981\,
            I => \POWERLED.func_state_RNI8H551Z0Z_0_cascade_\
        );

    \I__2420\ : IoInMux
    port map (
            O => \N__18978\,
            I => \N__18975\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__18975\,
            I => \N__18972\
        );

    \I__2418\ : IoSpan4Mux
    port map (
            O => \N__18972\,
            I => \N__18961\
        );

    \I__2417\ : InMux
    port map (
            O => \N__18971\,
            I => \N__18958\
        );

    \I__2416\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18955\
        );

    \I__2415\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18948\
        );

    \I__2414\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18948\
        );

    \I__2413\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18948\
        );

    \I__2412\ : InMux
    port map (
            O => \N__18966\,
            I => \N__18943\
        );

    \I__2411\ : InMux
    port map (
            O => \N__18965\,
            I => \N__18938\
        );

    \I__2410\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18938\
        );

    \I__2409\ : Span4Mux_s2_v
    port map (
            O => \N__18961\,
            I => \N__18933\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__18958\,
            I => \N__18933\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__18955\,
            I => \N__18928\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__18948\,
            I => \N__18928\
        );

    \I__2405\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18923\
        );

    \I__2404\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18923\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__18943\,
            I => rsmrstn
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__18938\,
            I => rsmrstn
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__18933\,
            I => rsmrstn
        );

    \I__2400\ : Odrv4
    port map (
            O => \N__18928\,
            I => rsmrstn
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__18923\,
            I => rsmrstn
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__18912\,
            I => \POWERLED.N_143_N_cascade_\
        );

    \I__2397\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18906\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__18903\,
            I => \POWERLED.N_116_f0\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__18900\,
            I => \POWERLED.N_116_f0_cascade_\
        );

    \I__2393\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18891\
        );

    \I__2392\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18891\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__18891\,
            I => \N__18888\
        );

    \I__2390\ : Odrv4
    port map (
            O => \N__18888\,
            I => \POWERLED.dutycycle_erZ0Z_9\
        );

    \I__2389\ : CEMux
    port map (
            O => \N__18885\,
            I => \N__18882\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__18882\,
            I => \N__18879\
        );

    \I__2387\ : Odrv4
    port map (
            O => \N__18879\,
            I => \POWERLED.dutycycle_en_2\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__18876\,
            I => \N__18868\
        );

    \I__2385\ : CascadeMux
    port map (
            O => \N__18875\,
            I => \N__18862\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__18874\,
            I => \N__18859\
        );

    \I__2383\ : InMux
    port map (
            O => \N__18873\,
            I => \N__18854\
        );

    \I__2382\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18854\
        );

    \I__2381\ : CascadeMux
    port map (
            O => \N__18871\,
            I => \N__18851\
        );

    \I__2380\ : InMux
    port map (
            O => \N__18868\,
            I => \N__18843\
        );

    \I__2379\ : InMux
    port map (
            O => \N__18867\,
            I => \N__18838\
        );

    \I__2378\ : InMux
    port map (
            O => \N__18866\,
            I => \N__18838\
        );

    \I__2377\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18835\
        );

    \I__2376\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18830\
        );

    \I__2375\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18830\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__18854\,
            I => \N__18827\
        );

    \I__2373\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18820\
        );

    \I__2372\ : InMux
    port map (
            O => \N__18850\,
            I => \N__18820\
        );

    \I__2371\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18820\
        );

    \I__2370\ : InMux
    port map (
            O => \N__18848\,
            I => \N__18817\
        );

    \I__2369\ : InMux
    port map (
            O => \N__18847\,
            I => \N__18812\
        );

    \I__2368\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18812\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__18843\,
            I => \N__18804\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__18838\,
            I => \N__18804\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18801\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__18830\,
            I => \N__18796\
        );

    \I__2363\ : Span4Mux_s2_h
    port map (
            O => \N__18827\,
            I => \N__18796\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__18820\,
            I => \N__18793\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__18817\,
            I => \N__18788\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__18812\,
            I => \N__18788\
        );

    \I__2359\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18781\
        );

    \I__2358\ : InMux
    port map (
            O => \N__18810\,
            I => \N__18781\
        );

    \I__2357\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18781\
        );

    \I__2356\ : Span4Mux_s3_v
    port map (
            O => \N__18804\,
            I => \N__18778\
        );

    \I__2355\ : Span4Mux_s2_h
    port map (
            O => \N__18801\,
            I => \N__18773\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__18796\,
            I => \N__18773\
        );

    \I__2353\ : Span4Mux_s3_h
    port map (
            O => \N__18793\,
            I => \N__18768\
        );

    \I__2352\ : Span4Mux_s3_h
    port map (
            O => \N__18788\,
            I => \N__18768\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__18781\,
            I => \N__18765\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__18778\,
            I => \POWERLED.N_3168_i\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__18773\,
            I => \POWERLED.N_3168_i\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__18768\,
            I => \POWERLED.N_3168_i\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__18765\,
            I => \POWERLED.N_3168_i\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__18756\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__18753\,
            I => \POWERLED.un1_clk_100khz_42_and_i_o2_1_1_cascade_\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__2343\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18743\
        );

    \I__2342\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18740\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__18743\,
            I => \N__18735\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18735\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__18735\,
            I => \POWERLED.N_171\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__18732\,
            I => \POWERLED.N_171_cascade_\
        );

    \I__2337\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18726\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__18726\,
            I => \POWERLED.N_387\
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__18723\,
            I => \POWERLED.dutycycle_m1_0_a2_0_cascade_\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__18720\,
            I => \N__18717\
        );

    \I__2333\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18714\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__18714\,
            I => \POWERLED.N_145_N\
        );

    \I__2331\ : InMux
    port map (
            O => \N__18711\,
            I => \N__18708\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__18708\,
            I => \N__18705\
        );

    \I__2329\ : Span4Mux_v
    port map (
            O => \N__18705\,
            I => \N__18702\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__18702\,
            I => \POWERLED.g1Z0Z_3\
        );

    \I__2327\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18696\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__18696\,
            I => \N__18693\
        );

    \I__2325\ : Span4Mux_v
    port map (
            O => \N__18693\,
            I => \N__18690\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__18690\,
            I => \POWERLED.g2_2\
        );

    \I__2323\ : InMux
    port map (
            O => \N__18687\,
            I => \N__18684\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__18684\,
            I => \N__18681\
        );

    \I__2321\ : Span4Mux_s3_h
    port map (
            O => \N__18681\,
            I => \N__18678\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__18678\,
            I => \POWERLED.func_state_1_m2_am_1_0\
        );

    \I__2319\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18672\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__18672\,
            I => \N__18669\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__18669\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3_out\
        );

    \I__2316\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18663\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__18663\,
            I => \N__18660\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__18660\,
            I => \POWERLED.un1_clk_100khz_2_i_o3_0\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__18657\,
            I => \POWERLED.func_state_RNI3IN21_1Z0Z_1_cascade_\
        );

    \I__2312\ : InMux
    port map (
            O => \N__18654\,
            I => \N__18651\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__18651\,
            I => \N__18644\
        );

    \I__2310\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18641\
        );

    \I__2309\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18638\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__18648\,
            I => \N__18631\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__18647\,
            I => \N__18626\
        );

    \I__2306\ : Span4Mux_h
    port map (
            O => \N__18644\,
            I => \N__18623\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18618\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__18638\,
            I => \N__18618\
        );

    \I__2303\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18613\
        );

    \I__2302\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18613\
        );

    \I__2301\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18610\
        );

    \I__2300\ : InMux
    port map (
            O => \N__18634\,
            I => \N__18599\
        );

    \I__2299\ : InMux
    port map (
            O => \N__18631\,
            I => \N__18599\
        );

    \I__2298\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18599\
        );

    \I__2297\ : InMux
    port map (
            O => \N__18629\,
            I => \N__18599\
        );

    \I__2296\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18599\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__18623\,
            I => \clk_100Khz_signalkeep_4_rep1\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__18618\,
            I => \clk_100Khz_signalkeep_4_rep1\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__18613\,
            I => \clk_100Khz_signalkeep_4_rep1\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__18610\,
            I => \clk_100Khz_signalkeep_4_rep1\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__18599\,
            I => \clk_100Khz_signalkeep_4_rep1\
        );

    \I__2290\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18585\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__18585\,
            I => \POWERLED.func_state_0_sqmuxa_0_o2_xZ0\
        );

    \I__2288\ : InMux
    port map (
            O => \N__18582\,
            I => \N__18579\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__18579\,
            I => \N__18576\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__18576\,
            I => \POWERLED.N_233_N\
        );

    \I__2285\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18565\
        );

    \I__2284\ : InMux
    port map (
            O => \N__18572\,
            I => \N__18553\
        );

    \I__2283\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18553\
        );

    \I__2282\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18553\
        );

    \I__2281\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18553\
        );

    \I__2280\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18553\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__18565\,
            I => \N__18550\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__18564\,
            I => \N__18545\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18541\
        );

    \I__2276\ : Span4Mux_s3_h
    port map (
            O => \N__18550\,
            I => \N__18538\
        );

    \I__2275\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18531\
        );

    \I__2274\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18531\
        );

    \I__2273\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18531\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__18544\,
            I => \N__18528\
        );

    \I__2271\ : Span4Mux_s3_h
    port map (
            O => \N__18541\,
            I => \N__18525\
        );

    \I__2270\ : Sp12to4
    port map (
            O => \N__18538\,
            I => \N__18520\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__18531\,
            I => \N__18520\
        );

    \I__2268\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18517\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__18525\,
            I => \curr_state_RNIR5QD1_0_0\
        );

    \I__2266\ : Odrv12
    port map (
            O => \N__18520\,
            I => \curr_state_RNIR5QD1_0_0\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__18517\,
            I => \curr_state_RNIR5QD1_0_0\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__18510\,
            I => \N__18507\
        );

    \I__2263\ : InMux
    port map (
            O => \N__18507\,
            I => \N__18504\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__18504\,
            I => \N__18501\
        );

    \I__2261\ : Span4Mux_s3_h
    port map (
            O => \N__18501\,
            I => \N__18497\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__18500\,
            I => \N__18492\
        );

    \I__2259\ : Span4Mux_v
    port map (
            O => \N__18497\,
            I => \N__18489\
        );

    \I__2258\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18485\
        );

    \I__2257\ : InMux
    port map (
            O => \N__18495\,
            I => \N__18480\
        );

    \I__2256\ : InMux
    port map (
            O => \N__18492\,
            I => \N__18480\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__18489\,
            I => \N__18477\
        );

    \I__2254\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18474\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__18485\,
            I => \N__18469\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__18480\,
            I => \N__18469\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__18477\,
            I => \clk_100Khz_signalkeep_4_fast\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__18474\,
            I => \clk_100Khz_signalkeep_4_fast\
        );

    \I__2249\ : Odrv12
    port map (
            O => \N__18469\,
            I => \clk_100Khz_signalkeep_4_fast\
        );

    \I__2248\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18453\
        );

    \I__2247\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18453\
        );

    \I__2246\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18453\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__18453\,
            I => \N__18450\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__18450\,
            I => \RSMRST_PWRGD_RSMRSTn_fast\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__18447\,
            I => \rsmrstn_cascade_\
        );

    \I__2242\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18441\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__18441\,
            I => \POWERLED.count_off_0_3\
        );

    \I__2240\ : InMux
    port map (
            O => \N__18438\,
            I => \N__18435\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__18435\,
            I => \POWERLED.count_off_0_0\
        );

    \I__2238\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18429\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__18429\,
            I => \N__18426\
        );

    \I__2236\ : Span4Mux_s3_h
    port map (
            O => \N__18426\,
            I => \N__18423\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__18423\,
            I => \POWERLED.func_state_RNI3IN21_2Z0Z_1\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__18420\,
            I => \N__18415\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__18419\,
            I => \N__18412\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__18418\,
            I => \N__18409\
        );

    \I__2231\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18405\
        );

    \I__2230\ : InMux
    port map (
            O => \N__18412\,
            I => \N__18398\
        );

    \I__2229\ : InMux
    port map (
            O => \N__18409\,
            I => \N__18398\
        );

    \I__2228\ : InMux
    port map (
            O => \N__18408\,
            I => \N__18395\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__18405\,
            I => \N__18392\
        );

    \I__2226\ : InMux
    port map (
            O => \N__18404\,
            I => \N__18387\
        );

    \I__2225\ : InMux
    port map (
            O => \N__18403\,
            I => \N__18387\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__18398\,
            I => \N__18384\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__18395\,
            I => \N__18381\
        );

    \I__2222\ : Odrv12
    port map (
            O => \N__18392\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__18387\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__18384\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__18381\,
            I => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__18372\,
            I => \POWERLED.N_425_cascade_\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__18369\,
            I => \POWERLED.N_175_cascade_\
        );

    \I__2216\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18363\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__18363\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_bm_1\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__18360\,
            I => \POWERLED.count_clk_en_0_cascade_\
        );

    \I__2213\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18354\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__18354\,
            I => \POWERLED.count_clk_en_2\
        );

    \I__2211\ : InMux
    port map (
            O => \N__18351\,
            I => \N__18348\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__18348\,
            I => \RSMRST_PWRGD.curr_state_2_0\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__18345\,
            I => \RSMRST_PWRGD.m4_0_0_cascade_\
        );

    \I__2208\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18336\
        );

    \I__2207\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18336\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__18336\,
            I => \N__18333\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__18333\,
            I => \RSMRST_PWRGD.N_423\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__18330\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__2203\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18324\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__18324\,
            I => \RSMRST_PWRGD.curr_state_7_1\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__18321\,
            I => \POWERLED.count_off_1_0_cascade_\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__18318\,
            I => \POWERLED.count_offZ0Z_0_cascade_\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__18315\,
            I => \POWERLED.count_off_RNIZ0Z_1_cascade_\
        );

    \I__2198\ : InMux
    port map (
            O => \N__18312\,
            I => \N__18309\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__18309\,
            I => \POWERLED.count_off_RNIZ0Z_1\
        );

    \I__2196\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18303\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__18303\,
            I => \POWERLED.count_off_0_1\
        );

    \I__2194\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18296\
        );

    \I__2193\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18293\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__18296\,
            I => \N__18290\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__18293\,
            I => \N__18287\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__18290\,
            I => \N__18284\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__18287\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__18284\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__2187\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18276\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__18276\,
            I => \N__18273\
        );

    \I__2185\ : Span4Mux_s3_h
    port map (
            O => \N__18273\,
            I => \N__18270\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__18270\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__18267\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__18264\,
            I => \curr_state_RNIR5QD1_0_0_cascade_\
        );

    \I__2181\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18258\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__18258\,
            I => \RSMRST_PWRGD.curr_state_1_1\
        );

    \I__2179\ : InMux
    port map (
            O => \N__18255\,
            I => \bfn_4_5_0_\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__18252\,
            I => \RSMRST_PWRGD.N_423_cascade_\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__18249\,
            I => \N__18246\
        );

    \I__2176\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18237\
        );

    \I__2175\ : InMux
    port map (
            O => \N__18245\,
            I => \N__18237\
        );

    \I__2174\ : InMux
    port map (
            O => \N__18244\,
            I => \N__18237\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__18237\,
            I => \N__18234\
        );

    \I__2172\ : Span4Mux_h
    port map (
            O => \N__18234\,
            I => \N__18231\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__18231\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__2170\ : InMux
    port map (
            O => \N__18228\,
            I => \N__18222\
        );

    \I__2169\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18222\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__18222\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__2167\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18213\
        );

    \I__2166\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18213\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__18213\,
            I => \N__18210\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__18210\,
            I => \N__18207\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__18207\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__2162\ : InMux
    port map (
            O => \N__18204\,
            I => \N__18201\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__18201\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__2160\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18195\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__18195\,
            I => \N__18191\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18188\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__18191\,
            I => \N__18185\
        );

    \I__2156\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18182\
        );

    \I__2155\ : Span4Mux_s1_h
    port map (
            O => \N__18185\,
            I => \N__18179\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__18182\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__18179\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__18174\,
            I => \N__18170\
        );

    \I__2151\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18166\
        );

    \I__2150\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18163\
        );

    \I__2149\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18160\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__18166\,
            I => \N__18157\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__18163\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__18160\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__18157\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__18150\,
            I => \N__18147\
        );

    \I__2143\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18144\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18141\
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__18141\,
            I => \PCH_PWRGD.N_278_0\
        );

    \I__2140\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18132\
        );

    \I__2139\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18132\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__18132\,
            I => \N__18129\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__18129\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__18126\,
            I => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0_cascade_\
        );

    \I__2135\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__18120\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__2133\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18113\
        );

    \I__2132\ : InMux
    port map (
            O => \N__18116\,
            I => \N__18110\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__18113\,
            I => \N__18107\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__18110\,
            I => \N__18104\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__18107\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__18104\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__18099\,
            I => \N__18095\
        );

    \I__2126\ : InMux
    port map (
            O => \N__18098\,
            I => \N__18087\
        );

    \I__2125\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18087\
        );

    \I__2124\ : InMux
    port map (
            O => \N__18094\,
            I => \N__18087\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__18087\,
            I => \PCH_PWRGD.N_3122_i\
        );

    \I__2122\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18076\
        );

    \I__2121\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18076\
        );

    \I__2120\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18073\
        );

    \I__2119\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18070\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__18076\,
            I => \PCH_PWRGD.N_3120_i\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__18073\,
            I => \PCH_PWRGD.N_3120_i\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__18070\,
            I => \PCH_PWRGD.N_3120_i\
        );

    \I__2115\ : InMux
    port map (
            O => \N__18063\,
            I => \N__18060\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__18060\,
            I => \PCH_PWRGD.N_413\
        );

    \I__2113\ : InMux
    port map (
            O => \N__18057\,
            I => \N__18045\
        );

    \I__2112\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18045\
        );

    \I__2111\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18045\
        );

    \I__2110\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18045\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__18045\,
            I => \N__18042\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__18042\,
            I => \N__18039\
        );

    \I__2107\ : Span4Mux_v
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__2106\ : Odrv4
    port map (
            O => \N__18036\,
            I => vr_ready_vccin
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__18033\,
            I => \PCH_PWRGD.N_413_cascade_\
        );

    \I__2104\ : InMux
    port map (
            O => \N__18030\,
            I => \N__18027\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__18027\,
            I => \PCH_PWRGD.N_277_0\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__18021\
        );

    \I__2101\ : InMux
    port map (
            O => \N__18021\,
            I => \N__18015\
        );

    \I__2100\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18015\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__18015\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__18012\,
            I => \N__18007\
        );

    \I__2097\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18001\
        );

    \I__2096\ : InMux
    port map (
            O => \N__18010\,
            I => \N__18001\
        );

    \I__2095\ : InMux
    port map (
            O => \N__18007\,
            I => \N__17996\
        );

    \I__2094\ : InMux
    port map (
            O => \N__18006\,
            I => \N__17996\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__18001\,
            I => \PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__17996\,
            I => \PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__17991\,
            I => \PCH_PWRGD.N_277_0_cascade_\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__17988\,
            I => \PCH_PWRGD.delayed_vccin_okZ0_cascade_\
        );

    \I__2089\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17982\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__2087\ : Span4Mux_s2_v
    port map (
            O => \N__17979\,
            I => \N__17976\
        );

    \I__2086\ : Span4Mux_s1_h
    port map (
            O => \N__17976\,
            I => \N__17973\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__17973\,
            I => \PCH_PWRGD.un12_clk_100khz_1\
        );

    \I__2084\ : InMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__2082\ : Span4Mux_s3_h
    port map (
            O => \N__17964\,
            I => \N__17961\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__17961\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__17958\,
            I => \PCH_PWRGD.N_3120_i_cascade_\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \PCH_PWRGD.curr_state_7_0_cascade_\
        );

    \I__2078\ : InMux
    port map (
            O => \N__17952\,
            I => \N__17949\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__17949\,
            I => \PCH_PWRGD.curr_state_1_0\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__17946\,
            I => \N__17942\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__17945\,
            I => \N__17936\
        );

    \I__2074\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17926\
        );

    \I__2073\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17926\
        );

    \I__2072\ : InMux
    port map (
            O => \N__17940\,
            I => \N__17926\
        );

    \I__2071\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17926\
        );

    \I__2070\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17922\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__17935\,
            I => \N__17915\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__17926\,
            I => \N__17904\
        );

    \I__2067\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17901\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__17922\,
            I => \N__17898\
        );

    \I__2065\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17889\
        );

    \I__2064\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17889\
        );

    \I__2063\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17889\
        );

    \I__2062\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17889\
        );

    \I__2061\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17880\
        );

    \I__2060\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17880\
        );

    \I__2059\ : InMux
    port map (
            O => \N__17913\,
            I => \N__17880\
        );

    \I__2058\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17880\
        );

    \I__2057\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17877\
        );

    \I__2056\ : InMux
    port map (
            O => \N__17910\,
            I => \N__17870\
        );

    \I__2055\ : InMux
    port map (
            O => \N__17909\,
            I => \N__17870\
        );

    \I__2054\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17870\
        );

    \I__2053\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17867\
        );

    \I__2052\ : Span4Mux_s1_v
    port map (
            O => \N__17904\,
            I => \N__17864\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__17901\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__17898\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__17889\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__17880\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__17877\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__17870\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__17867\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__17864\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__17847\,
            I => \PCH_PWRGD.curr_state_7_1_cascade_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__17844\,
            I => \N__17841\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__17841\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__2040\ : InMux
    port map (
            O => \N__17838\,
            I => \N__17826\
        );

    \I__2039\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17826\
        );

    \I__2038\ : InMux
    port map (
            O => \N__17836\,
            I => \N__17826\
        );

    \I__2037\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17826\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__17826\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__17823\,
            I => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__17820\,
            I => \POWERLED.un1_dutycycle_53_7_a0_2_0_cascade_\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__17817\,
            I => \N__17814\
        );

    \I__2032\ : InMux
    port map (
            O => \N__17814\,
            I => \N__17811\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__17811\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_3\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__17808\,
            I => \POWERLED.un1_dutycycle_53_34_1_cascade_\
        );

    \I__2029\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__17802\,
            I => \POWERLED.un1_dutycycle_53_34_0\
        );

    \I__2027\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__17796\,
            I => \POWERLED.un1_dutycycle_53_36_0\
        );

    \I__2025\ : CascadeMux
    port map (
            O => \N__17793\,
            I => \POWERLED.un1_m2_0_a0_0_cascade_\
        );

    \I__2024\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17787\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__17787\,
            I => \POWERLED.un1_m2_0_a0_1\
        );

    \I__2022\ : InMux
    port map (
            O => \N__17784\,
            I => \N__17775\
        );

    \I__2021\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17775\
        );

    \I__2020\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17775\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__17775\,
            I => \N__17772\
        );

    \I__2018\ : Span12Mux_s2_v
    port map (
            O => \N__17772\,
            I => \N__17767\
        );

    \I__2017\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17762\
        );

    \I__2016\ : InMux
    port map (
            O => \N__17770\,
            I => \N__17762\
        );

    \I__2015\ : Odrv12
    port map (
            O => \N__17767\,
            I => \POWERLED.N_371\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__17762\,
            I => \POWERLED.N_371\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__17757\,
            I => \POWERLED.N_371_cascade_\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__17754\,
            I => \POWERLED.N_372_cascade_\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__17751\,
            I => \POWERLED.un1_m5_2_cascade_\
        );

    \I__2010\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17745\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__17745\,
            I => \POWERLED.un1_dutycycle_53_30_0_0\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__17742\,
            I => \POWERLED.un1_dutycycle_53_30_1_cascade_\
        );

    \I__2007\ : InMux
    port map (
            O => \N__17739\,
            I => \N__17733\
        );

    \I__2006\ : InMux
    port map (
            O => \N__17738\,
            I => \N__17733\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__17733\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__17730\,
            I => \POWERLED.dutycycle_er_RNIT8CS1Z0Z_9_cascade_\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__17727\,
            I => \POWERLED.dutycycleZ1Z_9_cascade_\
        );

    \I__2002\ : InMux
    port map (
            O => \N__17724\,
            I => \N__17721\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__17721\,
            I => \POWERLED.dutycycle_i3_mux\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__17718\,
            I => \POWERLED.N_235_N_cascade_\
        );

    \I__1999\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17712\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__17712\,
            I => \POWERLED.N_434_N\
        );

    \I__1997\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17706\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__17706\,
            I => \POWERLED.N_235_N\
        );

    \I__1995\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17700\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__17700\,
            I => \POWERLED.un1_clk_100khz_42_and_i_a2_3_0\
        );

    \I__1993\ : InMux
    port map (
            O => \N__17697\,
            I => \N__17694\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__17694\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_2\
        );

    \I__1991\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17685\
        );

    \I__1990\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17685\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__17685\,
            I => \POWERLED.dutycycle_RNIHGUM6Z0Z_2\
        );

    \I__1988\ : InMux
    port map (
            O => \N__17682\,
            I => \N__17676\
        );

    \I__1987\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17676\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__17676\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__17673\,
            I => \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\
        );

    \I__1984\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17667\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__17667\,
            I => \POWERLED.N_301\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__17664\,
            I => \POWERLED.un1_func_state25_6_0_a2_0_cascade_\
        );

    \I__1981\ : InMux
    port map (
            O => \N__17661\,
            I => \N__17658\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__17658\,
            I => \POWERLED.un1_func_state25_6_0_2\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__17655\,
            I => \POWERLED.dutycycle_set_1_cascade_\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__17652\,
            I => \POWERLED.dutycycleZ1Z_5_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__17649\,
            I => \N__17646\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__17646\,
            I => \POWERLED.dutycycle_set_1\
        );

    \I__1975\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17637\
        );

    \I__1974\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17637\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__17637\,
            I => \N__17634\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__17634\,
            I => \POWERLED.dutycycle_eena_14_0_0_1\
        );

    \I__1971\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17628\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__17628\,
            I => \POWERLED.N_118_f0\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__17625\,
            I => \POWERLED.dutycycle_eena_3_0_0_sx_cascade_\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__17622\,
            I => \N__17619\
        );

    \I__1967\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17613\
        );

    \I__1966\ : InMux
    port map (
            O => \N__17618\,
            I => \N__17613\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__17613\,
            I => \N__17610\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__17610\,
            I => \POWERLED.N_393\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__17607\,
            I => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2_cascade_\
        );

    \I__1962\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17601\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__17601\,
            I => \N__17597\
        );

    \I__1960\ : InMux
    port map (
            O => \N__17600\,
            I => \N__17594\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__17597\,
            I => \POWERLED.dutycycle_RNI0DTG7Z0Z_6\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__17594\,
            I => \POWERLED.dutycycle_RNI0DTG7Z0Z_6\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__17589\,
            I => \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__17586\,
            I => \POWERLED.dutycycle_cascade_\
        );

    \I__1955\ : InMux
    port map (
            O => \N__17583\,
            I => \N__17580\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__17580\,
            I => \POWERLED.dutycycle_set_0_0\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__17577\,
            I => \POWERLED.dutycycle_set_0_0_cascade_\
        );

    \I__1952\ : InMux
    port map (
            O => \N__17574\,
            I => \N__17568\
        );

    \I__1951\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17568\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__17568\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__17565\,
            I => \POWERLED.N_346_cascade_\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__17562\,
            I => \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_\
        );

    \I__1947\ : InMux
    port map (
            O => \N__17559\,
            I => \N__17556\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__17556\,
            I => \POWERLED.func_state_RNIQBTF3_0Z0Z_1\
        );

    \I__1945\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17550\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__17550\,
            I => \N__17547\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__17547\,
            I => \POWERLED.func_state_1_ss0_i_0_o2_1\
        );

    \I__1942\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17541\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__17541\,
            I => \POWERLED.func_state_RNIQBTF3_1Z0Z_1\
        );

    \I__1940\ : InMux
    port map (
            O => \N__17538\,
            I => \N__17535\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__17535\,
            I => \POWERLED.N_343\
        );

    \I__1938\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17526\
        );

    \I__1937\ : InMux
    port map (
            O => \N__17531\,
            I => \N__17526\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__17526\,
            I => \RSMRST_PWRGD.count_5_1\
        );

    \I__1935\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17515\
        );

    \I__1934\ : CEMux
    port map (
            O => \N__17522\,
            I => \N__17515\
        );

    \I__1933\ : CEMux
    port map (
            O => \N__17521\,
            I => \N__17511\
        );

    \I__1932\ : CEMux
    port map (
            O => \N__17520\,
            I => \N__17504\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__17515\,
            I => \N__17500\
        );

    \I__1930\ : CEMux
    port map (
            O => \N__17514\,
            I => \N__17497\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__17511\,
            I => \N__17490\
        );

    \I__1928\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17482\
        );

    \I__1927\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17475\
        );

    \I__1926\ : InMux
    port map (
            O => \N__17508\,
            I => \N__17475\
        );

    \I__1925\ : CEMux
    port map (
            O => \N__17507\,
            I => \N__17475\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__17504\,
            I => \N__17472\
        );

    \I__1923\ : CEMux
    port map (
            O => \N__17503\,
            I => \N__17469\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__17500\,
            I => \N__17466\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__17497\,
            I => \N__17463\
        );

    \I__1920\ : CEMux
    port map (
            O => \N__17496\,
            I => \N__17460\
        );

    \I__1919\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17453\
        );

    \I__1918\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17453\
        );

    \I__1917\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17453\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__17490\,
            I => \N__17450\
        );

    \I__1915\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17447\
        );

    \I__1914\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17438\
        );

    \I__1913\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17438\
        );

    \I__1912\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17438\
        );

    \I__1911\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17438\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__17482\,
            I => \N__17423\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17423\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__17472\,
            I => \N__17420\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17415\
        );

    \I__1906\ : Sp12to4
    port map (
            O => \N__17466\,
            I => \N__17415\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__17463\,
            I => \N__17412\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__17460\,
            I => \N__17407\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__17453\,
            I => \N__17407\
        );

    \I__1902\ : Span4Mux_s1_h
    port map (
            O => \N__17450\,
            I => \N__17400\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17400\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__17438\,
            I => \N__17400\
        );

    \I__1899\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17391\
        );

    \I__1898\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17391\
        );

    \I__1897\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17391\
        );

    \I__1896\ : InMux
    port map (
            O => \N__17434\,
            I => \N__17391\
        );

    \I__1895\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17384\
        );

    \I__1894\ : InMux
    port map (
            O => \N__17432\,
            I => \N__17384\
        );

    \I__1893\ : InMux
    port map (
            O => \N__17431\,
            I => \N__17384\
        );

    \I__1892\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17377\
        );

    \I__1891\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17377\
        );

    \I__1890\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17377\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__17423\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__17420\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1887\ : Odrv12
    port map (
            O => \N__17415\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__17412\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1885\ : Odrv12
    port map (
            O => \N__17407\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__17400\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__17391\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__17384\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__17377\,
            I => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__17358\,
            I => \RSMRST_PWRGD.count_rst_6_cascade_\
        );

    \I__1879\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17350\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__17354\,
            I => \N__17347\
        );

    \I__1877\ : InMux
    port map (
            O => \N__17353\,
            I => \N__17344\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__17350\,
            I => \N__17340\
        );

    \I__1875\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17337\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__17344\,
            I => \N__17334\
        );

    \I__1873\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17331\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__17340\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__17337\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__17334\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__17331\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1868\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__17319\,
            I => \RSMRST_PWRGD.un12_clk_100khz_2\
        );

    \I__1866\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__17313\,
            I => \POWERLED.func_state_RNIAE974Z0Z_0\
        );

    \I__1864\ : CascadeMux
    port map (
            O => \N__17310\,
            I => \POWERLED.func_state_1_m2_am_1_1_cascade_\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__17307\,
            I => \POWERLED.func_state_1_m2s2_i_1_cascade_\
        );

    \I__1862\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17301\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__17301\,
            I => \POWERLED.N_79\
        );

    \I__1860\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17295\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__17295\,
            I => \POWERLED.func_state_RNIQTLM2Z0Z_1\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__17292\,
            I => \POWERLED.N_79_cascade_\
        );

    \I__1857\ : InMux
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__17286\,
            I => \POWERLED.func_state_1_m2_1\
        );

    \I__1855\ : InMux
    port map (
            O => \N__17283\,
            I => \N__17277\
        );

    \I__1854\ : InMux
    port map (
            O => \N__17282\,
            I => \N__17277\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__17277\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__1852\ : InMux
    port map (
            O => \N__17274\,
            I => \N__17267\
        );

    \I__1851\ : InMux
    port map (
            O => \N__17273\,
            I => \N__17267\
        );

    \I__1850\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17264\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__17267\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__17264\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__17259\,
            I => \POWERLED.func_state_1_m2_1_cascade_\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__17256\,
            I => \N__17252\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__17255\,
            I => \N__17249\
        );

    \I__1844\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17246\
        );

    \I__1843\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17243\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__17246\,
            I => \N__17240\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__17243\,
            I => \RSMRST_PWRGD.un2_count_1_axb_4\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__17240\,
            I => \RSMRST_PWRGD.un2_count_1_axb_4\
        );

    \I__1839\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17229\
        );

    \I__1838\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17229\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17226\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__17226\,
            I => \N__17223\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__17223\,
            I => \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1834\ : InMux
    port map (
            O => \N__17220\,
            I => \N__17214\
        );

    \I__1833\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17214\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__17214\,
            I => \RSMRST_PWRGD.count_5_4\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__17211\,
            I => \RSMRST_PWRGD.un2_count_1_axb_1_cascade_\
        );

    \I__1830\ : InMux
    port map (
            O => \N__17208\,
            I => \N__17205\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__17205\,
            I => \N__17202\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__17202\,
            I => \N__17198\
        );

    \I__1827\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17195\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__17198\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__17195\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__17190\,
            I => \N__17187\
        );

    \I__1823\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17183\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__17186\,
            I => \N__17180\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__17183\,
            I => \N__17177\
        );

    \I__1820\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17174\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__17177\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__17174\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1817\ : InMux
    port map (
            O => \N__17169\,
            I => \N__17165\
        );

    \I__1816\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17162\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__17165\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__17162\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1813\ : InMux
    port map (
            O => \N__17157\,
            I => \N__17154\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__17154\,
            I => \RSMRST_PWRGD.un12_clk_100khz_4\
        );

    \I__1811\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17148\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__17148\,
            I => \RSMRST_PWRGD.un12_clk_100khz_5\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__17145\,
            I => \RSMRST_PWRGD.un12_clk_100khz_11_cascade_\
        );

    \I__1808\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17139\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__17139\,
            I => \RSMRST_PWRGD.un12_clk_100khz_12\
        );

    \I__1806\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17133\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__17133\,
            I => \RSMRST_PWRGD.count_5_0\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__17130\,
            I => \RSMRST_PWRGD.countZ0Z_0_cascade_\
        );

    \I__1803\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17123\
        );

    \I__1802\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17120\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17117\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__17120\,
            I => \RSMRST_PWRGD.un2_count_1_axb_1\
        );

    \I__1799\ : Odrv4
    port map (
            O => \N__17117\,
            I => \RSMRST_PWRGD.un2_count_1_axb_1\
        );

    \I__1798\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17109\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__17109\,
            I => \RSMRST_PWRGD.count_rst_6\
        );

    \I__1796\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__1795\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17100\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__17100\,
            I => \RSMRST_PWRGD.count_rst_11\
        );

    \I__1793\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17094\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__17094\,
            I => \RSMRST_PWRGD.count_5_6\
        );

    \I__1791\ : InMux
    port map (
            O => \N__17091\,
            I => \N__17088\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__17088\,
            I => \RSMRST_PWRGD.count_5_7\
        );

    \I__1789\ : InMux
    port map (
            O => \N__17085\,
            I => \N__17081\
        );

    \I__1788\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17078\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__17081\,
            I => \RSMRST_PWRGD.count_rst_12\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__17078\,
            I => \RSMRST_PWRGD.count_rst_12\
        );

    \I__1785\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17070\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__17070\,
            I => \N__17067\
        );

    \I__1783\ : Odrv4
    port map (
            O => \N__17067\,
            I => \RSMRST_PWRGD.un2_count_1_axb_2\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__17064\,
            I => \RSMRST_PWRGD.un2_count_1_axb_4_cascade_\
        );

    \I__1781\ : InMux
    port map (
            O => \N__17061\,
            I => \N__17058\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__17058\,
            I => \RSMRST_PWRGD.count_rst_9\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__17055\,
            I => \RSMRST_PWRGD.count_rst_9_cascade_\
        );

    \I__1778\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17048\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__17051\,
            I => \N__17045\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__17048\,
            I => \N__17041\
        );

    \I__1775\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17038\
        );

    \I__1774\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17035\
        );

    \I__1773\ : Odrv12
    port map (
            O => \N__17041\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__17038\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__17035\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1770\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17025\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__17025\,
            I => \N__17022\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__17022\,
            I => \N__17019\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__17019\,
            I => \RSMRST_PWRGD.un12_clk_100khz_1\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__17016\,
            I => \RSMRST_PWRGD.un12_clk_100khz_0_cascade_\
        );

    \I__1765\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17007\
        );

    \I__1764\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17007\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__17007\,
            I => \RSMRST_PWRGD.count_5_2\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__17004\,
            I => \N__17000\
        );

    \I__1761\ : InMux
    port map (
            O => \N__17003\,
            I => \N__16992\
        );

    \I__1760\ : InMux
    port map (
            O => \N__17000\,
            I => \N__16992\
        );

    \I__1759\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16992\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__16992\,
            I => \N__16989\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__16989\,
            I => \RSMRST_PWRGD.count_rst_7\
        );

    \I__1756\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16983\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16979\
        );

    \I__1754\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16976\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__16979\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__16976\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1751\ : InMux
    port map (
            O => \N__16971\,
            I => \N__16968\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__16968\,
            I => \RSMRST_PWRGD.un12_clk_100khz_3\
        );

    \I__1749\ : InMux
    port map (
            O => \N__16965\,
            I => \N__16962\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__16962\,
            I => \N__16958\
        );

    \I__1747\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16955\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__16958\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__16955\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1744\ : InMux
    port map (
            O => \N__16950\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__1743\ : InMux
    port map (
            O => \N__16947\,
            I => \N__16941\
        );

    \I__1742\ : InMux
    port map (
            O => \N__16946\,
            I => \N__16941\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__16941\,
            I => \N__16938\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__16938\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__1739\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16931\
        );

    \I__1738\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16928\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__16931\,
            I => \N__16925\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__16928\,
            I => \RSMRST_PWRGD.count_rst_8\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__16925\,
            I => \RSMRST_PWRGD.count_rst_8\
        );

    \I__1734\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16917\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16914\
        );

    \I__1732\ : Span4Mux_s1_h
    port map (
            O => \N__16914\,
            I => \N__16911\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__16911\,
            I => \RSMRST_PWRGD.count_5_3\
        );

    \I__1730\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16905\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__16905\,
            I => \N__16901\
        );

    \I__1728\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16898\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__16901\,
            I => \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__16898\,
            I => \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\
        );

    \I__1725\ : InMux
    port map (
            O => \N__16893\,
            I => \N__16890\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__16890\,
            I => \N__16887\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__16887\,
            I => \RSMRST_PWRGD.count_5_13\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__16884\,
            I => \RSMRST_PWRGD.count_rst_2_cascade_\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__16881\,
            I => \RSMRST_PWRGD.count_rst_13_cascade_\
        );

    \I__1720\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16872\
        );

    \I__1719\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16872\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__16872\,
            I => \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__16869\,
            I => \RSMRST_PWRGD.countZ0Z_8_cascade_\
        );

    \I__1716\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16863\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__16863\,
            I => \RSMRST_PWRGD.count_5_8\
        );

    \I__1714\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16857\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__16857\,
            I => \N__16851\
        );

    \I__1712\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16844\
        );

    \I__1711\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16844\
        );

    \I__1710\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16844\
        );

    \I__1709\ : Odrv12
    port map (
            O => \N__16851\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__16844\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1707\ : InMux
    port map (
            O => \N__16839\,
            I => \N__16833\
        );

    \I__1706\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16833\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__16833\,
            I => \N__16830\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__16830\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__1703\ : InMux
    port map (
            O => \N__16827\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__1702\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16821\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__16821\,
            I => \N__16816\
        );

    \I__1700\ : InMux
    port map (
            O => \N__16820\,
            I => \N__16811\
        );

    \I__1699\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16811\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__16816\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__16811\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__16806\,
            I => \N__16802\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__16805\,
            I => \N__16799\
        );

    \I__1694\ : InMux
    port map (
            O => \N__16802\,
            I => \N__16794\
        );

    \I__1693\ : InMux
    port map (
            O => \N__16799\,
            I => \N__16794\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__16794\,
            I => \N__16791\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__16791\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1690\ : InMux
    port map (
            O => \N__16788\,
            I => \bfn_2_4_0_\
        );

    \I__1689\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16782\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__16782\,
            I => \N__16779\
        );

    \I__1687\ : Span4Mux_v
    port map (
            O => \N__16779\,
            I => \N__16774\
        );

    \I__1686\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16769\
        );

    \I__1685\ : InMux
    port map (
            O => \N__16777\,
            I => \N__16769\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__16774\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__16769\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1682\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16758\
        );

    \I__1681\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16758\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__16758\,
            I => \N__16755\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__16755\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1678\ : InMux
    port map (
            O => \N__16752\,
            I => \PCH_PWRGD.un2_count_1_cry_8\
        );

    \I__1677\ : InMux
    port map (
            O => \N__16749\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__1676\ : InMux
    port map (
            O => \N__16746\,
            I => \N__16742\
        );

    \I__1675\ : InMux
    port map (
            O => \N__16745\,
            I => \N__16739\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__16742\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__16739\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__16734\,
            I => \N__16730\
        );

    \I__1671\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16725\
        );

    \I__1670\ : InMux
    port map (
            O => \N__16730\,
            I => \N__16725\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__16725\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1668\ : InMux
    port map (
            O => \N__16722\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__1667\ : InMux
    port map (
            O => \N__16719\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__1666\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16712\
        );

    \I__1665\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16709\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__16712\,
            I => \N__16706\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__16709\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__16706\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1661\ : InMux
    port map (
            O => \N__16701\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__1660\ : InMux
    port map (
            O => \N__16698\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__1659\ : InMux
    port map (
            O => \N__16695\,
            I => \N__16692\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__16692\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__16689\,
            I => \N__16686\
        );

    \I__1656\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16683\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__16683\,
            I => \PCH_PWRGD.un2_count_1_axb_0\
        );

    \I__1654\ : InMux
    port map (
            O => \N__16680\,
            I => \PCH_PWRGD.un2_count_1_cry_0\
        );

    \I__1653\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16674\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__16674\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__1651\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16666\
        );

    \I__1650\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16661\
        );

    \I__1649\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16661\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__16666\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__16661\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1646\ : InMux
    port map (
            O => \N__16656\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__1645\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16649\
        );

    \I__1644\ : InMux
    port map (
            O => \N__16652\,
            I => \N__16645\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__16649\,
            I => \N__16642\
        );

    \I__1642\ : InMux
    port map (
            O => \N__16648\,
            I => \N__16639\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__16645\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__16642\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__16639\,
            I => \PCH_PWRGD.un2_count_1_axb_3\
        );

    \I__1638\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16628\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__16631\,
            I => \N__16625\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__16628\,
            I => \N__16622\
        );

    \I__1635\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16619\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__16622\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__16619\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__1632\ : InMux
    port map (
            O => \N__16614\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__1631\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16606\
        );

    \I__1630\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16601\
        );

    \I__1629\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16601\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__16606\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__16601\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__16596\,
            I => \N__16592\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__16595\,
            I => \N__16589\
        );

    \I__1624\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16584\
        );

    \I__1623\ : InMux
    port map (
            O => \N__16589\,
            I => \N__16584\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__16584\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1621\ : InMux
    port map (
            O => \N__16581\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__1620\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16575\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__16575\,
            I => \N__16571\
        );

    \I__1618\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16568\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__16571\,
            I => \PCH_PWRGD.un2_count_1_axb_5\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__16568\,
            I => \PCH_PWRGD.un2_count_1_axb_5\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__16563\,
            I => \N__16559\
        );

    \I__1614\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16554\
        );

    \I__1613\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16554\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__16551\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1610\ : InMux
    port map (
            O => \N__16548\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__16545\,
            I => \N__16541\
        );

    \I__1608\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16538\
        );

    \I__1607\ : InMux
    port map (
            O => \N__16541\,
            I => \N__16535\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__16538\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__16535\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1604\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16524\
        );

    \I__1603\ : InMux
    port map (
            O => \N__16529\,
            I => \N__16524\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__16524\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__1601\ : InMux
    port map (
            O => \N__16521\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__1600\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16512\
        );

    \I__1599\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16512\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__16512\,
            I => \PCH_PWRGD.count_rst_9\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__16509\,
            I => \PCH_PWRGD.un2_count_1_axb_5_cascade_\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__16506\,
            I => \N__16503\
        );

    \I__1595\ : InMux
    port map (
            O => \N__16503\,
            I => \N__16497\
        );

    \I__1594\ : InMux
    port map (
            O => \N__16502\,
            I => \N__16497\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__16497\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__1592\ : InMux
    port map (
            O => \N__16494\,
            I => \N__16491\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__16491\,
            I => \PCH_PWRGD.count_rst_11\
        );

    \I__1590\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16485\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__16485\,
            I => \N__16482\
        );

    \I__1588\ : Span4Mux_s2_h
    port map (
            O => \N__16482\,
            I => \N__16478\
        );

    \I__1587\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16475\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__16478\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__16475\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__16470\,
            I => \PCH_PWRGD.count_rst_11_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16463\
        );

    \I__1582\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16460\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__16463\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__16460\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1579\ : InMux
    port map (
            O => \N__16455\,
            I => \N__16452\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__16452\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__16449\,
            I => \POWERLED.g2_0_cascade_\
        );

    \I__1576\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16443\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__16443\,
            I => \N__16440\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__16440\,
            I => \POWERLED.g0_10_0_0_0\
        );

    \I__1573\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16434\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__16434\,
            I => \POWERLED.g0_8_1\
        );

    \I__1571\ : InMux
    port map (
            O => \N__16431\,
            I => \N__16428\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__16428\,
            I => \N__16425\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__16425\,
            I => \N__16422\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__16422\,
            I => \POWERLED.g1_1_0_1_0\
        );

    \I__1567\ : InMux
    port map (
            O => \N__16419\,
            I => \N__16413\
        );

    \I__1566\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16413\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__16413\,
            I => \POWERLED.un1_dutycycle_inv_4_0\
        );

    \I__1564\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16407\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__16407\,
            I => \PCH_PWRGD.un12_clk_100khz_5\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__16404\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__1561\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16398\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__16398\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__1559\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16392\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__16392\,
            I => \N__16389\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__16389\,
            I => \POWERLED.un1_dutycycle_164_0\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__16386\,
            I => \POWERLED.un1_dutycycle_172_m1_0_cascade_\
        );

    \I__1555\ : InMux
    port map (
            O => \N__16383\,
            I => \N__16380\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__16380\,
            I => \POWERLED.g0_0_m2_1\
        );

    \I__1553\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16374\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__16374\,
            I => \POWERLED.un1_dutycycle_172_m1_1_0\
        );

    \I__1551\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16368\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__16368\,
            I => \POWERLED.N_134\
        );

    \I__1549\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16362\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__16362\,
            I => \POWERLED.un1_dutycycle_168_0_0_1\
        );

    \I__1547\ : InMux
    port map (
            O => \N__16359\,
            I => \N__16356\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__16356\,
            I => \POWERLED.g1_1_0\
        );

    \I__1545\ : CascadeMux
    port map (
            O => \N__16353\,
            I => \POWERLED.g2_0_1_cascade_\
        );

    \I__1544\ : InMux
    port map (
            O => \N__16350\,
            I => \N__16347\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__16347\,
            I => \N__16344\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__16344\,
            I => \POWERLED.g0_10_0_0_1\
        );

    \I__1541\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16338\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__16338\,
            I => \POWERLED.g2_1\
        );

    \I__1539\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16332\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__16332\,
            I => \POWERLED.un1_dutycycle_172_m0_0\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__16329\,
            I => \POWERLED.g2_0_0_1_0_cascade_\
        );

    \I__1536\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16323\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__16323\,
            I => \N__16320\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__16320\,
            I => \POWERLED.N_237\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__16317\,
            I => \POWERLED.N_3297_0_0_0_cascade_\
        );

    \I__1532\ : InMux
    port map (
            O => \N__16314\,
            I => \N__16311\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__16311\,
            I => \POWERLED.g1_0_1_0_1\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__16308\,
            I => \N__16305\
        );

    \I__1529\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16302\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__16302\,
            I => \N__16299\
        );

    \I__1527\ : Odrv12
    port map (
            O => \N__16299\,
            I => \POWERLED.N_3297_0_0_2\
        );

    \I__1526\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16293\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__16293\,
            I => \POWERLED.un1_dutycycle_172_m3_0_0_0\
        );

    \I__1524\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16287\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__16287\,
            I => \N__16284\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__16284\,
            I => \POWERLED.un1_clk_100khz_52_and_i_0\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__16281\,
            I => \POWERLED.un1_clk_100khz_52_and_i_o2_0_0_1_cascade_\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__16278\,
            I => \POWERLED.dutycycle_eena_0_cascade_\
        );

    \I__1519\ : InMux
    port map (
            O => \N__16275\,
            I => \N__16272\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__16272\,
            I => \POWERLED.dutycycle_1_0_1\
        );

    \I__1517\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16263\
        );

    \I__1516\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16263\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__16263\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__16260\,
            I => \POWERLED.g0_18_1_cascade_\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__16257\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16251\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__16251\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_5\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__16248\,
            I => \N__16243\
        );

    \I__1509\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16238\
        );

    \I__1508\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16238\
        );

    \I__1507\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16235\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__16238\,
            I => \N__16232\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__16235\,
            I => \N__16229\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__16232\,
            I => \N__16225\
        );

    \I__1503\ : Span4Mux_s1_h
    port map (
            O => \N__16229\,
            I => \N__16222\
        );

    \I__1502\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16219\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__16225\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__1500\ : Odrv4
    port map (
            O => \N__16222\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__16219\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_0\
        );

    \I__1498\ : InMux
    port map (
            O => \N__16212\,
            I => \N__16209\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__16209\,
            I => vpp_ok
        );

    \I__1496\ : IoInMux
    port map (
            O => \N__16206\,
            I => \N__16203\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__16203\,
            I => \N__16200\
        );

    \I__1494\ : Span4Mux_s0_v
    port map (
            O => \N__16200\,
            I => \N__16197\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__16197\,
            I => vddq_en
        );

    \I__1492\ : InMux
    port map (
            O => \N__16194\,
            I => \N__16191\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__16191\,
            I => \POWERLED.N_189_i\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__16188\,
            I => \POWERLED.dutycycleZ0Z_1_cascade_\
        );

    \I__1489\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16182\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__16182\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__16179\,
            I => \POWERLED.dutycycle_eena_cascade_\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__16176\,
            I => \N__16172\
        );

    \I__1485\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16169\
        );

    \I__1484\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16166\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__16169\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__16166\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__16161\,
            I => \POWERLED.dutycycle_1_0_1_cascade_\
        );

    \I__1480\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16152\
        );

    \I__1479\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16152\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__16152\,
            I => \POWERLED.dutycycle_1_0_0\
        );

    \I__1477\ : InMux
    port map (
            O => \N__16149\,
            I => \N__16143\
        );

    \I__1476\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16143\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__16143\,
            I => \POWERLED.N_120_f0_1\
        );

    \I__1474\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16137\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__16137\,
            I => \POWERLED.dutycycle_eena_0\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__16134\,
            I => \POWERLED.un1_func_state25_6_0_a3_1_cascade_\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__16131\,
            I => \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__16128\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__16125\,
            I => \POWERLED.N_189_i_cascade_\
        );

    \I__1468\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16119\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__16119\,
            I => \N__16116\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__16116\,
            I => \POWERLED.N_238\
        );

    \I__1465\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16110\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__16110\,
            I => \POWERLED.func_state_1_m2_0\
        );

    \I__1463\ : InMux
    port map (
            O => \N__16107\,
            I => \N__16101\
        );

    \I__1462\ : InMux
    port map (
            O => \N__16106\,
            I => \N__16101\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__16101\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__16098\,
            I => \POWERLED.func_state_1_m2_0_cascade_\
        );

    \I__1459\ : IoInMux
    port map (
            O => \N__16095\,
            I => \N__16092\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__16092\,
            I => vccst_en
        );

    \I__1457\ : InMux
    port map (
            O => \N__16089\,
            I => \N__16086\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__16086\,
            I => \RSMRST_PWRGD.N_240_0\
        );

    \I__1455\ : InMux
    port map (
            O => \N__16083\,
            I => \N__16080\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16077\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__16077\,
            I => \N__16074\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__16074\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1451\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16065\
        );

    \I__1450\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16065\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__16065\,
            I => \N__16061\
        );

    \I__1448\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16058\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__16061\,
            I => \RSMRST_PWRGD.count_rst_1\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__16058\,
            I => \RSMRST_PWRGD.count_rst_1\
        );

    \I__1445\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16049\
        );

    \I__1444\ : InMux
    port map (
            O => \N__16052\,
            I => \N__16046\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__16049\,
            I => \N__16043\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__16046\,
            I => \RSMRST_PWRGD.count_5_12\
        );

    \I__1441\ : Odrv12
    port map (
            O => \N__16043\,
            I => \RSMRST_PWRGD.count_5_12\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__16038\,
            I => \RSMRST_PWRGD.countZ0Z_15_cascade_\
        );

    \I__1439\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16029\
        );

    \I__1438\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16029\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__16029\,
            I => \N__16026\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__16026\,
            I => \RSMRST_PWRGD.count_rst_4\
        );

    \I__1435\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16020\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__16020\,
            I => \RSMRST_PWRGD.count_5_15\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__16017\,
            I => \POWERLED.func_state_enZ0_cascade_\
        );

    \I__1432\ : InMux
    port map (
            O => \N__16014\,
            I => \RSMRST_PWRGD.un2_count_1_cry_14\
        );

    \I__1431\ : InMux
    port map (
            O => \N__16011\,
            I => \N__16008\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__16008\,
            I => \RSMRST_PWRGD.un2_count_1_axb_12\
        );

    \I__1429\ : InMux
    port map (
            O => \N__16005\,
            I => \N__16002\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__16002\,
            I => \N__15999\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__15999\,
            I => \RSMRST_PWRGD.un2_count_1_axb_5\
        );

    \I__1426\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15993\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__15993\,
            I => \RSMRST_PWRGD.count_5_14\
        );

    \I__1424\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15984\
        );

    \I__1423\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15984\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__15984\,
            I => \RSMRST_PWRGD.count_rst_3\
        );

    \I__1421\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15978\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__15978\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1419\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15966\
        );

    \I__1418\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15966\
        );

    \I__1417\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15966\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__15966\,
            I => \N__15963\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__15963\,
            I => \RSMRST_PWRGD.count_rst_10\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__15960\,
            I => \RSMRST_PWRGD.countZ0Z_14_cascade_\
        );

    \I__1413\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15951\
        );

    \I__1412\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15951\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__15951\,
            I => \RSMRST_PWRGD.count_5_5\
        );

    \I__1410\ : InMux
    port map (
            O => \N__15948\,
            I => \N__15942\
        );

    \I__1409\ : InMux
    port map (
            O => \N__15947\,
            I => \N__15942\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__15942\,
            I => \RSMRST_PWRGD.count_rst_0\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15939\,
            I => \N__15936\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__15936\,
            I => \RSMRST_PWRGD.count_5_11\
        );

    \I__1405\ : InMux
    port map (
            O => \N__15933\,
            I => \RSMRST_PWRGD.un2_count_1_cry_5\
        );

    \I__1404\ : InMux
    port map (
            O => \N__15930\,
            I => \RSMRST_PWRGD.un2_count_1_cry_6\
        );

    \I__1403\ : InMux
    port map (
            O => \N__15927\,
            I => \RSMRST_PWRGD.un2_count_1_cry_7\
        );

    \I__1402\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15920\
        );

    \I__1401\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15917\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__15920\,
            I => \N__15914\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__15917\,
            I => \RSMRST_PWRGD.un2_count_1_axb_9\
        );

    \I__1398\ : Odrv12
    port map (
            O => \N__15914\,
            I => \RSMRST_PWRGD.un2_count_1_axb_9\
        );

    \I__1397\ : InMux
    port map (
            O => \N__15909\,
            I => \N__15903\
        );

    \I__1396\ : InMux
    port map (
            O => \N__15908\,
            I => \N__15903\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__15903\,
            I => \N__15900\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__15900\,
            I => \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1393\ : InMux
    port map (
            O => \N__15897\,
            I => \bfn_1_6_0_\
        );

    \I__1392\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15889\
        );

    \I__1391\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15884\
        );

    \I__1390\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15884\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__15889\,
            I => \N__15881\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__15884\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1387\ : Odrv4
    port map (
            O => \N__15881\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__15876\,
            I => \N__15872\
        );

    \I__1385\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15869\
        );

    \I__1384\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15866\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__15869\,
            I => \N__15861\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__15866\,
            I => \N__15861\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__15861\,
            I => \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO\
        );

    \I__1380\ : InMux
    port map (
            O => \N__15858\,
            I => \RSMRST_PWRGD.un2_count_1_cry_9\
        );

    \I__1379\ : InMux
    port map (
            O => \N__15855\,
            I => \RSMRST_PWRGD.un2_count_1_cry_10\
        );

    \I__1378\ : InMux
    port map (
            O => \N__15852\,
            I => \RSMRST_PWRGD.un2_count_1_cry_11\
        );

    \I__1377\ : InMux
    port map (
            O => \N__15849\,
            I => \RSMRST_PWRGD.un2_count_1_cry_12\
        );

    \I__1376\ : InMux
    port map (
            O => \N__15846\,
            I => \RSMRST_PWRGD.un2_count_1_cry_13\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__15843\,
            I => \RSMRST_PWRGD.count_rst_cascade_\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__15840\,
            I => \RSMRST_PWRGD.countZ0Z_10_cascade_\
        );

    \I__1373\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15834\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__15834\,
            I => \RSMRST_PWRGD.count_5_10\
        );

    \I__1371\ : InMux
    port map (
            O => \N__15831\,
            I => \RSMRST_PWRGD.un2_count_1_cry_1\
        );

    \I__1370\ : InMux
    port map (
            O => \N__15828\,
            I => \RSMRST_PWRGD.un2_count_1_cry_2\
        );

    \I__1369\ : InMux
    port map (
            O => \N__15825\,
            I => \RSMRST_PWRGD.un2_count_1_cry_3\
        );

    \I__1368\ : InMux
    port map (
            O => \N__15822\,
            I => \RSMRST_PWRGD.un2_count_1_cry_4\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__15819\,
            I => \PCH_PWRGD.count_rst_3_cascade_\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \PCH_PWRGD.un2_count_1_axb_11_cascade_\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__15813\,
            I => \N__15810\
        );

    \I__1364\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15804\
        );

    \I__1363\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15804\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__15804\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__1361\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15798\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__15798\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__15795\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__15792\,
            I => \PCH_PWRGD.countZ0Z_4_cascade_\
        );

    \I__1357\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15786\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__15783\,
            I => \PCH_PWRGD.un12_clk_100khz_4\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__15780\,
            I => \RSMRST_PWRGD.un2_count_1_axb_9_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15774\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__15774\,
            I => \RSMRST_PWRGD.count_rst_14\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__15771\,
            I => \RSMRST_PWRGD.count_rst_14_cascade_\
        );

    \I__1350\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15762\
        );

    \I__1349\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15762\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__15762\,
            I => \RSMRST_PWRGD.count_5_9\
        );

    \I__1347\ : InMux
    port map (
            O => \N__15759\,
            I => \N__15756\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__15756\,
            I => \PCH_PWRGD.count_rst_14\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__15753\,
            I => \PCH_PWRGD.count_i_0_cascade_\
        );

    \I__1344\ : InMux
    port map (
            O => \N__15750\,
            I => \N__15747\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__15747\,
            I => \PCH_PWRGD.un12_clk_100khz_0\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__15744\,
            I => \PCH_PWRGD.un12_clk_100khz_9_cascade_\
        );

    \I__1341\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15738\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__15738\,
            I => \PCH_PWRGD.un12_clk_100khz_13\
        );

    \I__1339\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15729\
        );

    \I__1338\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15729\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__15729\,
            I => \PCH_PWRGD.count_i_0\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__15726\,
            I => \PCH_PWRGD.N_1_i_cascade_\
        );

    \I__1335\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15717\
        );

    \I__1334\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15717\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__15717\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__1332\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15711\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15708\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__15708\,
            I => \PCH_PWRGD.un12_clk_100khz_7\
        );

    \I__1329\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15702\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__15702\,
            I => \PCH_PWRGD.count_rst_3\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__15699\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__15696\,
            I => \PCH_PWRGD.countZ0Z_9_cascade_\
        );

    \I__1325\ : InMux
    port map (
            O => \N__15693\,
            I => \N__15690\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__15690\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__1323\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__15684\,
            I => \PCH_PWRGD.count_rst_6\
        );

    \I__1321\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15677\
        );

    \I__1320\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15674\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__15677\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__15674\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__15669\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__15666\,
            I => \PCH_PWRGD.un12_clk_100khz_6_cascade_\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__15663\,
            I => \PCH_PWRGD.count_rst_14_cascade_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un4_count_1_cry_8\,
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_16_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_9_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un2_count_1_cry_8\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un2_count_1_cry_16\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un2_count_1_cry_7\,
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \HDA_STRAP.count_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27147\,
            GLOBALBUFFEROUTPUT => \HDA_STRAP.count_en_g\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32559\,
            GLOBALBUFFEROUTPUT => \VPP_VDDQ_delayed_vddq_pwrgd_en_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNIPPJS1_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__17919\,
            in1 => \N__16763\,
            in2 => \N__24378\,
            in3 => \N__16778\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI64K95_9_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29876\,
            in1 => \_gnd_net_\,
            in2 => \N__15699\,
            in3 => \N__15693\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => \PCH_PWRGD.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_9_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__24346\,
            in2 => \N__15696\,
            in3 => \N__16764\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38412\,
            ce => \N__29879\,
            sr => \N__24389\
        );

    \PCH_PWRGD.count_8_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16820\,
            in1 => \N__24345\,
            in2 => \N__16806\,
            in3 => \N__17921\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38412\,
            ce => \N__29879\,
            sr => \N__24389\
        );

    \PCH_PWRGD.count_RNI41J95_8_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15687\,
            in1 => \N__29875\,
            in2 => \_gnd_net_\,
            in3 => \N__15680\,
            lcout => \PCH_PWRGD.un2_count_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNIONIS1_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16819\,
            in1 => \N__24344\,
            in2 => \N__16805\,
            in3 => \N__17918\,
            lcout => \PCH_PWRGD.count_rst_6\,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI41J95_0_8_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__15681\,
            in1 => \N__29877\,
            in2 => \N__15669\,
            in3 => \N__16777\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIK379L_3_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15714\,
            in1 => \N__16410\,
            in2 => \N__15666\,
            in3 => \N__15789\,
            lcout => \PCH_PWRGD.un12_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIUVFS4_0_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__15734\,
            in1 => \N__24335\,
            in2 => \_gnd_net_\,
            in3 => \N__17907\,
            lcout => \PCH_PWRGD.count_rst_14\,
            ltout => \PCH_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15723\,
            in2 => \N__15663\,
            in3 => \N__29866\,
            lcout => \PCH_PWRGD.un2_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOEC95_0_2_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__29867\,
            in1 => \N__16467\,
            in2 => \N__16545\,
            in3 => \N__16669\,
            lcout => \PCH_PWRGD.un12_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI410D3_0_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__15759\,
            in1 => \N__15722\,
            in2 => \_gnd_net_\,
            in3 => \N__29865\,
            lcout => \PCH_PWRGD.count_i_0\,
            ltout => \PCH_PWRGD.count_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI410D3_0_0_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__16715\,
            in1 => \N__29733\,
            in2 => \N__15753\,
            in3 => \N__16961\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un12_clk_100khz_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIV3OH31_2_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17985\,
            in1 => \N__15750\,
            in2 => \N__15744\,
            in3 => \N__15741\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => \PCH_PWRGD.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__15735\,
            in1 => \_gnd_net_\,
            in2 => \N__15726\,
            in3 => \N__24336\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38611\,
            ce => \N__29894\,
            sr => \N__24379\
        );

    \PCH_PWRGD.count_2_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16670\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38611\,
            ce => \N__29894\,
            sr => \N__24379\
        );

    \PCH_PWRGD.count_RNIOOMC5_0_11_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__15705\,
            in1 => \N__29832\,
            in2 => \N__15813\,
            in3 => \N__18117\,
            lcout => \PCH_PWRGD.un12_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__24339\,
            in1 => \N__16610\,
            in2 => \N__16596\,
            in3 => \N__17910\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38514\,
            ce => \N__29878\,
            sr => \N__24371\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNI237N1_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__17908\,
            in1 => \N__16745\,
            in2 => \N__16734\,
            in3 => \N__24337\,
            lcout => \PCH_PWRGD.count_rst_3\,
            ltout => \PCH_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOOMC5_11_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__29830\,
            in1 => \_gnd_net_\,
            in2 => \N__15819\,
            in3 => \N__15809\,
            lcout => \PCH_PWRGD.un2_count_1_axb_11\,
            ltout => \PCH_PWRGD.un2_count_1_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_11_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16733\,
            in1 => \N__17925\,
            in2 => \N__15816\,
            in3 => \N__24340\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38514\,
            ce => \N__29878\,
            sr => \N__24371\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNIKFES1_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__24338\,
            in1 => \N__16609\,
            in2 => \N__16595\,
            in3 => \N__17909\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISKE95_4_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__15801\,
            in1 => \N__29831\,
            in2 => \N__15795\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => \PCH_PWRGD.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQHD95_0_3_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__29833\,
            in1 => \N__16494\,
            in2 => \N__15792\,
            in3 => \N__16488\,
            lcout => \PCH_PWRGD.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIMCS06_9_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15767\,
            in1 => \N__15777\,
            in2 => \_gnd_net_\,
            in3 => \N__17493\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_9\,
            ltout => \RSMRST_PWRGD.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20408\,
            in1 => \N__15908\,
            in2 => \N__15780\,
            in3 => \N__20515\,
            lcout => \RSMRST_PWRGD.count_rst_14\,
            ltout => \RSMRST_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__15768\,
            in1 => \N__15892\,
            in2 => \N__15771\,
            in3 => \N__17495\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_9_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__15923\,
            in1 => \N__15909\,
            in2 => \N__20431\,
            in3 => \N__20518\,
            lcout => \RSMRST_PWRGD.count_5_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38622\,
            ce => \N__17514\,
            sr => \N__20407\
        );

    \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__20516\,
            in1 => \N__20409\,
            in2 => \N__15876\,
            in3 => \N__15893\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.count_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIV86M5_10_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17494\,
            in1 => \_gnd_net_\,
            in2 => \N__15843\,
            in3 => \N__15837\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => \RSMRST_PWRGD.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_10_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__20517\,
            in1 => \N__20410\,
            in2 => \N__15840\,
            in3 => \N__15875\,
            lcout => \RSMRST_PWRGD.count_5_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38622\,
            ce => \N__17514\,
            sr => \N__20407\
        );

    \RSMRST_PWRGD.count_13_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__20519\,
            in1 => \N__16908\,
            in2 => \N__20430\,
            in3 => \N__17353\,
            lcout => \RSMRST_PWRGD.count_5_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38622\,
            ce => \N__17514\,
            sr => \N__20407\
        );

    \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17127\,
            in2 => \N__20247\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20356\,
            in1 => \N__17073\,
            in2 => \_gnd_net_\,
            in3 => \N__15831\,
            lcout => \RSMRST_PWRGD.count_rst_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20358\,
            in1 => \N__16986\,
            in2 => \_gnd_net_\,
            in3 => \N__15828\,
            lcout => \RSMRST_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17256\,
            in3 => \N__15825\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20359\,
            in1 => \N__16005\,
            in2 => \_gnd_net_\,
            in3 => \N__15822\,
            lcout => \RSMRST_PWRGD.count_rst_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20357\,
            in1 => \N__17201\,
            in2 => \_gnd_net_\,
            in3 => \N__15933\,
            lcout => \RSMRST_PWRGD.count_rst_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__20360\,
            in1 => \_gnd_net_\,
            in2 => \N__17186\,
            in3 => \N__15930\,
            lcout => \RSMRST_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17044\,
            in2 => \_gnd_net_\,
            in3 => \N__15927\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_7\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15924\,
            in2 => \_gnd_net_\,
            in3 => \N__15897\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15894\,
            in2 => \_gnd_net_\,
            in3 => \N__15858\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20404\,
            in1 => \N__17168\,
            in2 => \_gnd_net_\,
            in3 => \N__15855\,
            lcout => \RSMRST_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20378\,
            in1 => \N__16011\,
            in2 => \_gnd_net_\,
            in3 => \N__15852\,
            lcout => \RSMRST_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17343\,
            in2 => \_gnd_net_\,
            in3 => \N__15849\,
            lcout => \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20379\,
            in1 => \N__15981\,
            in2 => \_gnd_net_\,
            in3 => \N__15846\,
            lcout => \RSMRST_PWRGD.count_rst_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un2_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16083\,
            in1 => \N__20380\,
            in2 => \_gnd_net_\,
            in3 => \N__16014\,
            lcout => \RSMRST_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIA43M5_12_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16053\,
            in1 => \N__16064\,
            in2 => \_gnd_net_\,
            in3 => \N__17489\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_14_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_5_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => \N__17496\,
            sr => \N__20405\
        );

    \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15956\,
            in1 => \N__17435\,
            in2 => \_gnd_net_\,
            in3 => \N__15973\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_5_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15974\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => \N__17496\,
            sr => \N__20405\
        );

    \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15996\,
            in1 => \N__17437\,
            in2 => \_gnd_net_\,
            in3 => \N__15989\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => \RSMRST_PWRGD.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000111"
        )
    port map (
            in0 => \N__15975\,
            in1 => \N__17510\,
            in2 => \N__15960\,
            in3 => \N__15957\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI812M5_11_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15939\,
            in1 => \N__17436\,
            in2 => \_gnd_net_\,
            in3 => \N__15947\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_11_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_5_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38589\,
            ce => \N__17496\,
            sr => \N__20405\
        );

    \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16920\,
            in1 => \N__17434\,
            in2 => \_gnd_net_\,
            in3 => \N__16935\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__16089\,
            in1 => \N__20375\,
            in2 => \N__19751\,
            in3 => \N__36046\,
            lcout => \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_12_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16070\,
            lcout => \RSMRST_PWRGD.count_5_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38581\,
            ce => \N__17507\,
            sr => \N__20406\
        );

    \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__32220\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19692\,
            lcout => \RSMRST_PWRGD.N_240_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIGD6M5_15_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17509\,
            in1 => \N__16023\,
            in2 => \_gnd_net_\,
            in3 => \N__16035\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => \RSMRST_PWRGD.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__16071\,
            in1 => \N__16052\,
            in2 => \N__16038\,
            in3 => \N__17508\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_15_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16034\,
            lcout => \RSMRST_PWRGD.count_5_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38581\,
            ce => \N__17507\,
            sr => \N__20406\
        );

    \POWERLED.func_state_en_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__32287\,
            in1 => \N__19265\,
            in2 => \_gnd_net_\,
            in3 => \N__36041\,
            lcout => \POWERLED.func_state_enZ0\,
            ltout => \POWERLED.func_state_enZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__36172\,
            in1 => \N__16113\,
            in2 => \N__16017\,
            in3 => \N__16107\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38576\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.G_146_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18635\,
            in2 => \_gnd_net_\,
            in3 => \N__19908\,
            lcout => \VPP_VDDQ_delayed_vddq_pwrgd_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI4Q6N7_1_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17316\,
            in1 => \N__17304\,
            in2 => \_gnd_net_\,
            in3 => \N__17544\,
            lcout => \POWERLED.func_state_1_m2_0\,
            ltout => \POWERLED.func_state_1_m2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8V1IA_0_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__16106\,
            in1 => \N__36171\,
            in2 => \N__16098\,
            in3 => \N__17272\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__29316\,
            in1 => \N__29270\,
            in2 => \_gnd_net_\,
            in3 => \N__29456\,
            lcout => \VPP_VDDQ.N_297_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29271\,
            in1 => \N__29315\,
            in2 => \N__29460\,
            in3 => \N__33367\,
            lcout => \VPP_VDDQ.count_2_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_0_i_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__19267\,
            in1 => \N__18568\,
            in2 => \N__19644\,
            in3 => \N__33390\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_0_o3_0_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101111111"
        )
    port map (
            in0 => \N__18569\,
            in1 => \N__19268\,
            in2 => \N__18647\,
            in3 => \N__19637\,
            lcout => \VCCST_EN_i_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.slp_s3n_signal_i_0_o3_2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101011111"
        )
    port map (
            in0 => \N__19638\,
            in1 => \N__18572\,
            in2 => \N__19137\,
            in3 => \N__18629\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_rep1_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18634\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19920\,
            lcout => \clk_100Khz_signalkeep_4_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__19132\,
            in1 => \N__18571\,
            in2 => \N__19272\,
            in3 => \N__18630\,
            lcout => \POWERLED.N_188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__18570\,
            in1 => \N__18675\,
            in2 => \N__18648\,
            in3 => \N__19639\,
            lcout => \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_0_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19133\,
            in1 => \N__20565\,
            in2 => \N__16248\,
            in3 => \N__19383\,
            lcout => \POWERLED.func_state_RNI2MQDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__36439\,
            in1 => \N__22692\,
            in2 => \_gnd_net_\,
            in3 => \N__18848\,
            lcout => \POWERLED.N_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__18404\,
            in1 => \_gnd_net_\,
            in2 => \N__19392\,
            in3 => \N__25109\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBADV5_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__16247\,
            in1 => \N__17661\,
            in2 => \N__16134\,
            in3 => \N__32569\,
            lcout => \POWERLED.dutycycle_RNIBADV5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI0TA81_0_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110111011"
        )
    port map (
            in0 => \N__18403\,
            in1 => \N__25160\,
            in2 => \N__19391\,
            in3 => \N__16246\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3F2B2_1_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__25108\,
            in1 => \_gnd_net_\,
            in2 => \N__16131\,
            in3 => \N__18432\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3P2F3_1_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33023\,
            in2 => \N__16128\,
            in3 => \N__32280\,
            lcout => \POWERLED.N_189_i\,
            ltout => \POWERLED.N_189_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3MDN4_2_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__32281\,
            in1 => \N__19246\,
            in2 => \N__16125\,
            in3 => \N__16122\,
            lcout => \POWERLED.N_118_f0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3MDN4_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101011"
        )
    port map (
            in0 => \N__16194\,
            in1 => \N__32282\,
            in2 => \N__19264\,
            in3 => \N__35497\,
            lcout => \POWERLED.N_120_f0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31RH1_5_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__32283\,
            in1 => \N__19245\,
            in2 => \N__33024\,
            in3 => \N__16326\,
            lcout => \POWERLED.un1_clk_100khz_52_and_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNISCB09_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__16157\,
            in1 => \N__32570\,
            in2 => \N__16176\,
            in3 => \N__16185\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => \POWERLED.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNICTP07_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111101"
        )
    port map (
            in0 => \N__23646\,
            in1 => \N__32301\,
            in2 => \N__16188\,
            in3 => \N__16148\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => \POWERLED.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__16158\,
            in1 => \N__32572\,
            in2 => \N__16179\,
            in3 => \N__16175\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => 'H',
            sr => \N__23334\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110011"
        )
    port map (
            in0 => \N__20584\,
            in1 => \N__20934\,
            in2 => \N__18418\,
            in3 => \N__22743\,
            lcout => \POWERLED.dutycycle_1_0_1\,
            ltout => \POWERLED.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI0O919_1_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__16140\,
            in1 => \N__32571\,
            in2 => \N__16161\,
            in3 => \N__16268\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0TA81_0_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__22746\,
            in1 => \N__31355\,
            in2 => \N__18419\,
            in3 => \N__20585\,
            lcout => \POWERLED.dutycycle_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNICTP07_1_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110011"
        )
    port map (
            in0 => \N__16149\,
            in1 => \N__23647\,
            in2 => \N__32316\,
            in3 => \N__36815\,
            lcout => \POWERLED.dutycycle_eena_0\,
            ltout => \POWERLED.dutycycle_eena_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__16269\,
            in1 => \N__32602\,
            in2 => \N__16278\,
            in3 => \N__16275\,
            lcout => \POWERLED.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38621\,
            ce => 'H',
            sr => \N__23334\
        );

    \POWERLED.dutycycle_RNI_7_5_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__36761\,
            in1 => \N__25633\,
            in2 => \_gnd_net_\,
            in3 => \N__17771\,
            lcout => OPEN,
            ltout => \POWERLED.g0_18_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_0_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__36817\,
            in1 => \N__31360\,
            in2 => \N__16260\,
            in3 => \N__29048\,
            lcout => \POWERLED.un1_dutycycle_164_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__29047\,
            in1 => \N__17770\,
            in2 => \N__31375\,
            in3 => \N__36816\,
            lcout => \POWERLED.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_5_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__28928\,
            in1 => \N__31361\,
            in2 => \N__36854\,
            in3 => \N__29046\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_5\,
            ltout => \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__18865\,
            in1 => \N__20586\,
            in2 => \N__16257\,
            in3 => \N__16228\,
            lcout => \POWERLED.func_state_RNIZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_5_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19368\,
            in2 => \_gnd_net_\,
            in3 => \N__16254\,
            lcout => \POWERLED.dutycycle_RNI_8Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_0_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__31359\,
            in1 => \N__29101\,
            in2 => \N__36855\,
            in3 => \N__25632\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16212\,
            in2 => \_gnd_net_\,
            in3 => \N__36189\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI64F52_5_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011011100"
        )
    port map (
            in0 => \N__36749\,
            in1 => \N__18699\,
            in2 => \N__25121\,
            in3 => \N__16371\,
            lcout => \POWERLED.un1_dutycycle_172_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_0_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000101"
        )
    port map (
            in0 => \N__16341\,
            in1 => \N__36750\,
            in2 => \N__25122\,
            in3 => \N__25176\,
            lcout => OPEN,
            ltout => \POWERLED.g2_0_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVB8J4_5_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__28929\,
            in1 => \N__16335\,
            in2 => \N__16329\,
            in3 => \N__16314\,
            lcout => \POWERLED.un1_dutycycle_172_m3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_0_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__25114\,
            in1 => \N__16350\,
            in2 => \N__36760\,
            in3 => \N__22332\,
            lcout => \POWERLED.N_3297_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_5_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000101"
        )
    port map (
            in0 => \N__28930\,
            in1 => \_gnd_net_\,
            in2 => \N__18871\,
            in3 => \N__22747\,
            lcout => \POWERLED.N_237\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_1_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__25113\,
            in1 => \N__16446\,
            in2 => \N__36759\,
            in3 => \N__22331\,
            lcout => OPEN,
            ltout => \POWERLED.N_3297_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIP7PD2_1_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__18850\,
            in1 => \N__16431\,
            in2 => \N__16317\,
            in3 => \N__23546\,
            lcout => \POWERLED.g1_0_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_1_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22742\,
            in2 => \_gnd_net_\,
            in3 => \N__18849\,
            lcout => \POWERLED.func_state_RNI_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5D218_0_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110111"
        )
    port map (
            in0 => \N__16383\,
            in1 => \N__16365\,
            in2 => \N__16308\,
            in3 => \N__16296\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_52_and_i_o2_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHL9SB_0_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111111111"
        )
    port map (
            in0 => \N__16290\,
            in1 => \N__32300\,
            in2 => \N__16281\,
            in3 => \N__23683\,
            lcout => \POWERLED.dutycycle_eena_14_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3F2B2_2_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010001000"
        )
    port map (
            in0 => \N__23542\,
            in1 => \N__16418\,
            in2 => \N__18420\,
            in3 => \N__16377\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI61QD3_0_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__18867\,
            in1 => \N__16395\,
            in2 => \N__16386\,
            in3 => \N__23544\,
            lcout => \POWERLED.g0_0_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_2_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111011101"
        )
    port map (
            in0 => \N__25646\,
            in1 => \N__16419\,
            in2 => \N__18876\,
            in3 => \N__36459\,
            lcout => \POWERLED.un1_dutycycle_172_m1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3IN21_0_5_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__18866\,
            in1 => \N__23543\,
            in2 => \_gnd_net_\,
            in3 => \N__25645\,
            lcout => \POWERLED.N_134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5DLR_2_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__19097\,
            in1 => \N__19216\,
            in2 => \_gnd_net_\,
            in3 => \N__36458\,
            lcout => \POWERLED.g0_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_0_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__29119\,
            in1 => \N__16359\,
            in2 => \N__31421\,
            in3 => \N__25177\,
            lcout => \POWERLED.un1_dutycycle_168_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_1_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__36869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17784\,
            lcout => \POWERLED.g1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_1_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__17783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36867\,
            lcout => OPEN,
            ltout => \POWERLED.g2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_0_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010001"
        )
    port map (
            in0 => \N__25178\,
            in1 => \N__31415\,
            in2 => \N__16353\,
            in3 => \N__29120\,
            lcout => \POWERLED.g0_10_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_0_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__17782\,
            in1 => \_gnd_net_\,
            in2 => \N__31422\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_1_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__36868\,
            in1 => \N__25179\,
            in2 => \N__16449\,
            in3 => \N__29121\,
            lcout => \POWERLED.g0_10_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIML1B1_2_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__16437\,
            in1 => \N__18573\,
            in2 => \N__18510\,
            in3 => \N__19643\,
            lcout => \POWERLED.g1_1_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_0_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25881\,
            in1 => \N__31416\,
            in2 => \N__36878\,
            in3 => \N__36762\,
            lcout => \POWERLED.un1_dutycycle_inv_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__16855\,
            in1 => \N__24363\,
            in2 => \N__17945\,
            in3 => \N__16838\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38320\,
            ce => \N__29904\,
            sr => \N__24387\
        );

    \PCH_PWRGD.count_RNIUNF95_0_5_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__29887\,
            in1 => \N__16517\,
            in2 => \N__16506\,
            in3 => \N__16854\,
            lcout => \PCH_PWRGD.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNILHFS1_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16574\,
            in1 => \N__24362\,
            in2 => \N__16563\,
            in3 => \N__17912\,
            lcout => \PCH_PWRGD.count_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNINLHS1_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__16839\,
            in1 => \N__16856\,
            in2 => \N__17935\,
            in3 => \N__24388\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI2UH95_7_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29886\,
            in2 => \N__16404\,
            in3 => \N__16401\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIUNF95_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__16502\,
            in1 => \N__16518\,
            in2 => \N__29896\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.un2_count_1_axb_5\,
            ltout => \PCH_PWRGD.un2_count_1_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_5_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16562\,
            in1 => \N__24364\,
            in2 => \N__16509\,
            in3 => \N__17914\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38320\,
            ce => \N__29904\,
            sr => \N__24387\
        );

    \PCH_PWRGD.count_3_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__17913\,
            in1 => \N__16632\,
            in2 => \N__24386\,
            in3 => \N__16653\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38320\,
            ce => \N__29904\,
            sr => \N__24387\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNIJDDS1_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__16648\,
            in1 => \N__24361\,
            in2 => \N__16631\,
            in3 => \N__17911\,
            lcout => \PCH_PWRGD.count_rst_11\,
            ltout => \PCH_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQHD95_3_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16481\,
            in2 => \N__16470\,
            in3 => \N__29868\,
            lcout => \PCH_PWRGD.un2_count_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOEC95_2_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29870\,
            in1 => \N__16466\,
            in2 => \_gnd_net_\,
            in3 => \N__16671\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI05RC5_15_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__16946\,
            in1 => \N__29873\,
            in2 => \_gnd_net_\,
            in3 => \N__16455\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16947\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__29872\,
            sr => \N__24390\
        );

    \PCH_PWRGD.count_RNI0RG95_6_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16530\,
            in1 => \N__16695\,
            in2 => \_gnd_net_\,
            in3 => \N__29871\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16529\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38610\,
            ce => \N__29872\,
            sr => \N__24390\
        );

    \PCH_PWRGD.count_RNISUOC5_13_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18279\,
            in1 => \N__18299\,
            in2 => \_gnd_net_\,
            in3 => \N__29869\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_0_c_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16689\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_0_c_RNIH9BS1_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24368\,
            in1 => \N__18116\,
            in2 => \_gnd_net_\,
            in3 => \N__16680\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_0\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNIIBCS1_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24369\,
            in1 => \N__16677\,
            in2 => \_gnd_net_\,
            in3 => \N__16656\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16652\,
            in2 => \_gnd_net_\,
            in3 => \N__16614\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16611\,
            in2 => \_gnd_net_\,
            in3 => \N__16581\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16578\,
            in2 => \_gnd_net_\,
            in3 => \N__16548\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNIMJGS1_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24370\,
            in1 => \N__16544\,
            in2 => \_gnd_net_\,
            in3 => \N__16521\,
            lcout => \PCH_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16860\,
            in2 => \_gnd_net_\,
            in3 => \N__16827\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16824\,
            in2 => \_gnd_net_\,
            in3 => \N__16788\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16785\,
            in2 => \_gnd_net_\,
            in3 => \N__16752\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIQRKS1_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24357\,
            in1 => \N__17970\,
            in2 => \_gnd_net_\,
            in3 => \N__16749\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16746\,
            in2 => \_gnd_net_\,
            in3 => \N__16722\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNI358N1_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24358\,
            in1 => \N__18198\,
            in2 => \_gnd_net_\,
            in3 => \N__16719\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNI479N1_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24372\,
            in1 => \N__16716\,
            in2 => \_gnd_net_\,
            in3 => \N__16701\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNI59AN1_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24359\,
            in1 => \N__29729\,
            in2 => \_gnd_net_\,
            in3 => \N__16698\,
            lcout => \PCH_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNI6BBN1_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16965\,
            in1 => \N__24360\,
            in2 => \_gnd_net_\,
            in3 => \N__16950\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_3_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16934\,
            lcout => \RSMRST_PWRGD.count_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38473\,
            ce => \N__17521\,
            sr => \N__20373\
        );

    \RSMRST_PWRGD.count_7_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17085\,
            lcout => \RSMRST_PWRGD.count_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38473\,
            ce => \N__17521\,
            sr => \N__20373\
        );

    \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20384\,
            in1 => \N__16904\,
            in2 => \N__17354\,
            in3 => \N__20494\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.count_rst_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIC74M5_13_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16893\,
            in2 => \N__16884\,
            in3 => \N__17488\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20383\,
            in1 => \N__16877\,
            in2 => \N__17051\,
            in3 => \N__20493\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIK9R06_8_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16866\,
            in2 => \N__16881\,
            in3 => \N__17487\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => \RSMRST_PWRGD.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_8_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20433\,
            in1 => \N__16878\,
            in2 => \N__16869\,
            in3 => \N__20495\,
            lcout => \RSMRST_PWRGD.count_5_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38422\,
            ce => \N__17520\,
            sr => \N__20432\
        );

    \RSMRST_PWRGD.count_RNIG3P06_6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17097\,
            in1 => \N__17105\,
            in2 => \_gnd_net_\,
            in3 => \N__17485\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_6_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17106\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38422\,
            ce => \N__17520\,
            sr => \N__20432\
        );

    \RSMRST_PWRGD.count_RNII6Q06_7_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17091\,
            in1 => \N__17084\,
            in2 => \_gnd_net_\,
            in3 => \N__17486\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_2_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.count_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38557\,
            ce => \N__17522\,
            sr => \N__20436\
        );

    \RSMRST_PWRGD.count_RNI8NK06_2_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17012\,
            in1 => \N__16999\,
            in2 => \_gnd_net_\,
            in3 => \N__17431\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNICTM06_4_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17433\,
            in1 => \N__17219\,
            in2 => \_gnd_net_\,
            in3 => \N__17061\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_4\,
            ltout => \RSMRST_PWRGD.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20376\,
            in1 => \N__17234\,
            in2 => \N__17064\,
            in3 => \N__20466\,
            lcout => \RSMRST_PWRGD.count_rst_9\,
            ltout => \RSMRST_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNICTM06_0_4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__17523\,
            in1 => \N__17220\,
            in2 => \N__17055\,
            in3 => \N__17052\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un12_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI91BKN_1_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17028\,
            in1 => \N__17322\,
            in2 => \N__17016\,
            in3 => \N__16971\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__17432\,
            in1 => \N__17013\,
            in2 => \N__17004\,
            in3 => \N__16982\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_4_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__20377\,
            in1 => \N__20467\,
            in2 => \N__17255\,
            in3 => \N__17235\,
            lcout => \RSMRST_PWRGD.count_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38557\,
            ce => \N__17522\,
            sr => \N__20436\
        );

    \RSMRST_PWRGD.count_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20435\,
            in1 => \N__20232\,
            in2 => \_gnd_net_\,
            in3 => \N__20489\,
            lcout => \RSMRST_PWRGD.count_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38529\,
            ce => \N__17503\,
            sr => \N__20434\
        );

    \RSMRST_PWRGD.count_RNIVV2I5_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17531\,
            in1 => \N__17429\,
            in2 => \_gnd_net_\,
            in3 => \N__17112\,
            lcout => \RSMRST_PWRGD.un2_count_1_axb_1\,
            ltout => \RSMRST_PWRGD.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20231\,
            in2 => \N__17211\,
            in3 => \N__20382\,
            lcout => \RSMRST_PWRGD.count_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38529\,
            ce => \N__17503\,
            sr => \N__20434\
        );

    \RSMRST_PWRGD.count_RNI_11_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20233\,
            in1 => \N__17208\,
            in2 => \N__17190\,
            in3 => \N__17169\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un12_clk_100khz_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI166B31_12_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17157\,
            in1 => \N__17151\,
            in2 => \N__17145\,
            in3 => \N__17142\,
            lcout => \RSMRST_PWRGD.count_RNI166B31Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIUU2I5_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17136\,
            in1 => \N__17428\,
            in2 => \_gnd_net_\,
            in3 => \N__20208\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => \RSMRST_PWRGD.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIAB7J1_1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20381\,
            in2 => \N__17130\,
            in3 => \N__17126\,
            lcout => \RSMRST_PWRGD.count_rst_6\,
            ltout => \RSMRST_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__17532\,
            in1 => \N__17430\,
            in2 => \N__17358\,
            in3 => \N__17355\,
            lcout => \RSMRST_PWRGD.un12_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__17274\,
            in1 => \N__17289\,
            in2 => \N__36188\,
            in3 => \N__17283\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38574\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIAE974_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100110011"
        )
    port map (
            in0 => \N__35466\,
            in1 => \N__18687\,
            in2 => \N__32832\,
            in3 => \N__22615\,
            lcout => \POWERLED.func_state_RNIAE974Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIC1SE1_1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__22689\,
            in1 => \N__23678\,
            in2 => \_gnd_net_\,
            in3 => \N__35465\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m2_am_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQTLM2_1_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001111"
        )
    port map (
            in0 => \N__18872\,
            in1 => \N__32828\,
            in2 => \N__17310\,
            in3 => \N__22614\,
            lcout => \POWERLED.func_state_RNIQTLM2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010001"
        )
    port map (
            in0 => \N__22690\,
            in1 => \N__18873\,
            in2 => \N__35433\,
            in3 => \N__17538\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m2s2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQBTF3_1_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110111"
        )
    port map (
            in0 => \N__23679\,
            in1 => \N__32890\,
            in2 => \N__17307\,
            in3 => \N__22691\,
            lcout => \POWERLED.N_79\,
            ltout => \POWERLED.N_79_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIK9J66_1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17298\,
            in2 => \N__17292\,
            in3 => \N__17559\,
            lcout => \POWERLED.func_state_1_m2_1\,
            ltout => \POWERLED.func_state_1_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIPFE19_1_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__17282\,
            in1 => \N__17273\,
            in2 => \N__17259\,
            in3 => \N__36173\,
            lcout => \POWERLED.func_state\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001001110"
        )
    port map (
            in0 => \N__17600\,
            in1 => \N__17574\,
            in2 => \N__23693\,
            in3 => \N__17583\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38533\,
            ce => 'H',
            sr => \N__23311\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIMU422_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__25120\,
            in1 => \N__23545\,
            in2 => \N__32867\,
            in3 => \N__20856\,
            lcout => \POWERLED.dutycycle_set_0_0\,
            ltout => \POWERLED.dutycycle_set_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMCG8B_6_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111000100"
        )
    port map (
            in0 => \N__23670\,
            in1 => \N__17604\,
            in2 => \N__17577\,
            in3 => \N__17573\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_0_0_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17618\,
            in1 => \N__22611\,
            in2 => \_gnd_net_\,
            in3 => \N__18846\,
            lcout => OPEN,
            ltout => \POWERLED.N_346_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIFJJH2_1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110111"
        )
    port map (
            in0 => \N__22612\,
            in1 => \N__23667\,
            in2 => \N__17565\,
            in3 => \N__25074\,
            lcout => \POWERLED.func_state_1_ss0_i_0_o2_1\,
            ltout => \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQBTF3_0_1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101011"
        )
    port map (
            in0 => \N__35468\,
            in1 => \N__32868\,
            in2 => \N__17562\,
            in3 => \N__22723\,
            lcout => \POWERLED.func_state_RNIQBTF3_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQBTF3_1_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__17553\,
            in1 => \N__32855\,
            in2 => \N__35467\,
            in3 => \N__22688\,
            lcout => \POWERLED.func_state_RNIQBTF3_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_0_1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22687\,
            in1 => \N__18847\,
            in2 => \N__17622\,
            in3 => \N__22613\,
            lcout => \POWERLED.N_343\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_229_i_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32972\,
            in1 => \N__33368\,
            in2 => \N__22837\,
            in3 => \N__18969\,
            lcout => \POWERLED.N_229_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHGUM6_2_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__32594\,
            in1 => \N__23645\,
            in2 => \_gnd_net_\,
            in3 => \N__17631\,
            lcout => \POWERLED.dutycycle_RNIHGUM6Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIESP71_0_0_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110111"
        )
    port map (
            in0 => \N__32974\,
            in1 => \N__18637\,
            in2 => \N__22839\,
            in3 => \N__24887\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_3_0_0_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8FSS1_0_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__24888\,
            in1 => \N__18970\,
            in2 => \N__17625\,
            in3 => \N__19919\,
            lcout => \POWERLED.dutycycle_eena_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_ss0_i_0_a2_3_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__19130\,
            in1 => \N__19243\,
            in2 => \_gnd_net_\,
            in3 => \N__18968\,
            lcout => \POWERLED.N_393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__19244\,
            in1 => \N__19131\,
            in2 => \_gnd_net_\,
            in3 => \N__22693\,
            lcout => \POWERLED.un1_clk_100khz_2_i_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__32973\,
            in1 => \N__18967\,
            in2 => \N__22838\,
            in3 => \N__18636\,
            lcout => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2\,
            ltout => \POWERLED.func_state_0_sqmuxa_0_oZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI0DTG7_6_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001010"
        )
    port map (
            in0 => \N__32595\,
            in1 => \N__18582\,
            in2 => \N__17607\,
            in3 => \N__35391\,
            lcout => \POWERLED.dutycycle_RNI0DTG7Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIGIKL1_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__22745\,
            in1 => \N__17670\,
            in2 => \N__19129\,
            in3 => \N__20916\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_0_2\,
            ltout => \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKGSL9_2_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__17681\,
            in1 => \N__18746\,
            in2 => \N__17589\,
            in3 => \N__17690\,
            lcout => \POWERLED.dutycycle\,
            ltout => \POWERLED.dutycycle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17586\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__17682\,
            in1 => \N__17697\,
            in2 => \N__18750\,
            in3 => \N__17691\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38550\,
            ce => 'H',
            sr => \N__23297\
        );

    \POWERLED.func_state_RNI34G9_0_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__32975\,
            in1 => \_gnd_net_\,
            in2 => \N__18874\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIESP71_1_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18650\,
            in1 => \N__22827\,
            in2 => \N__17673\,
            in3 => \N__22744\,
            lcout => \POWERLED.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_1_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__19113\,
            in1 => \_gnd_net_\,
            in2 => \N__18875\,
            in3 => \N__33011\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__22549\,
            in1 => \N__36180\,
            in2 => \N__17664\,
            in3 => \N__20724\,
            lcout => \POWERLED.un1_func_state25_6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI1UVG3_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011111"
        )
    port map (
            in0 => \N__23669\,
            in1 => \N__20868\,
            in2 => \N__32891\,
            in3 => \N__25119\,
            lcout => \POWERLED.dutycycle_set_1\,
            ltout => \POWERLED.dutycycle_set_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI7BG4G_5_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__32603\,
            in1 => \N__17738\,
            in2 => \N__17655\,
            in3 => \N__17642\,
            lcout => \POWERLED.dutycycleZ1Z_5\,
            ltout => \POWERLED.dutycycleZ1Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_5_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17652\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__17649\,
            in1 => \N__17643\,
            in2 => \N__32637\,
            in3 => \N__17739\,
            lcout => \POWERLED.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38618\,
            ce => 'H',
            sr => \N__23330\
        );

    \POWERLED.dutycycle_er_RNIT8CS1_9_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__18649\,
            in1 => \N__18896\,
            in2 => \N__21012\,
            in3 => \N__19918\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_er_RNIT8CS1Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_er_RNISPEN9_9_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18909\,
            in2 => \N__17730\,
            in3 => \N__17724\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => \POWERLED.dutycycleZ1Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_5_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__28927\,
            in1 => \N__29082\,
            in2 => \N__17727\,
            in3 => \N__20958\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_er_RNI9A8B3_9_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__18897\,
            in1 => \N__23668\,
            in2 => \N__32636\,
            in3 => \N__21008\,
            lcout => \POWERLED.dutycycle_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM6QF4_12_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110011"
        )
    port map (
            in0 => \N__17715\,
            in1 => \N__23015\,
            in2 => \N__26561\,
            in3 => \N__26448\,
            lcout => \POWERLED.N_235_N\,
            ltout => \POWERLED.N_235_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFJJH2_11_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100111111"
        )
    port map (
            in0 => \N__23540\,
            in1 => \N__23674\,
            in2 => \N__17718\,
            in3 => \N__26476\,
            lcout => \POWERLED.dutycycle_eena_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3IN21_2_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__17703\,
            in1 => \N__23539\,
            in2 => \N__25175\,
            in3 => \N__36419\,
            lcout => \POWERLED.N_434_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFJJH2_12_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111011111"
        )
    port map (
            in0 => \N__23541\,
            in1 => \N__26543\,
            in2 => \N__23694\,
            in3 => \N__17709\,
            lcout => \POWERLED.dutycycle_eena_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_14_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19343\,
            in1 => \_gnd_net_\,
            in2 => \N__25782\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_clk_100khz_42_and_i_a2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__26449\,
            in1 => \N__26544\,
            in2 => \_gnd_net_\,
            in3 => \N__25778\,
            lcout => \POWERLED.N_371\,
            ltout => \POWERLED.N_371_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17757\,
            in3 => \N__36418\,
            lcout => \POWERLED.N_372\,
            ltout => \POWERLED.N_372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_0_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17754\,
            in3 => \N__19342\,
            lcout => \POWERLED.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26148\,
            in1 => \N__23214\,
            in2 => \N__25555\,
            in3 => \N__26369\,
            lcout => OPEN,
            ltout => \POWERLED.un1_m5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_7_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17751\,
            in3 => \N__28591\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__28590\,
            in1 => \N__29112\,
            in2 => \N__28867\,
            in3 => \N__28688\,
            lcout => \POWERLED.un1_dutycycle_53_30_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__28854\,
            in1 => \N__23209\,
            in2 => \N__29145\,
            in3 => \N__26147\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_30_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_3_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17748\,
            in1 => \N__21185\,
            in2 => \N__17742\,
            in3 => \N__19422\,
            lcout => \POWERLED.dutycycle_RNI_11Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_11_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100110101"
        )
    port map (
            in0 => \N__26368\,
            in1 => \N__25544\,
            in2 => \N__26568\,
            in3 => \N__26146\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_7_a0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000010101"
        )
    port map (
            in0 => \N__26472\,
            in1 => \N__25861\,
            in2 => \N__17820\,
            in3 => \N__26565\,
            lcout => \POWERLED.un1_dutycycle_53_7_a0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__25557\,
            in1 => \N__23210\,
            in2 => \N__17817\,
            in3 => \N__28592\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_8_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__28842\,
            in1 => \N__23207\,
            in2 => \N__21186\,
            in3 => \N__29118\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_34_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \N__26566\,
            in1 => \N__17805\,
            in2 => \N__17808\,
            in3 => \N__17799\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_7_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001010"
        )
    port map (
            in0 => \N__28586\,
            in1 => \N__23204\,
            in2 => \N__25863\,
            in3 => \N__29117\,
            lcout => \POWERLED.un1_dutycycle_53_34_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_8_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__23205\,
            in1 => \_gnd_net_\,
            in2 => \N__26177\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_53_36_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_10_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__26394\,
            in1 => \N__23206\,
            in2 => \N__26478\,
            in3 => \N__26153\,
            lcout => OPEN,
            ltout => \POWERLED.un1_m2_0_a0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_7_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011010000"
        )
    port map (
            in0 => \N__21216\,
            in1 => \N__17790\,
            in2 => \N__17793\,
            in3 => \N__28588\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_7_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010101111111"
        )
    port map (
            in0 => \N__28841\,
            in1 => \N__26149\,
            in2 => \N__28593\,
            in3 => \N__29116\,
            lcout => \POWERLED.un1_m2_0_a0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010000000"
        )
    port map (
            in0 => \N__23203\,
            in1 => \N__28582\,
            in2 => \N__28690\,
            in3 => \N__28840\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18169\,
            lcout => \PCH_PWRGD.N_3120_i\,
            ltout => \PCH_PWRGD.N_3120_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__17836\,
            in1 => \N__24409\,
            in2 => \N__17958\,
            in3 => \N__17941\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38319\,
            ce => \N__35994\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__18006\,
            in1 => \N__17837\,
            in2 => \N__17946\,
            in3 => \N__18084\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIA9ET1_0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17952\,
            in2 => \N__17955\,
            in3 => \N__33263\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__17940\,
            in1 => \N__17835\,
            in2 => \N__18012\,
            in3 => \N__18083\,
            lcout => \PCH_PWRGD.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38319\,
            ce => \N__35994\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__17838\,
            in1 => \N__18081\,
            in2 => \N__24416\,
            in3 => \N__17939\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.curr_state_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIBAET1_1_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33264\,
            in1 => \_gnd_net_\,
            in2 => \N__17847\,
            in3 => \N__17844\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17823\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_3122_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__18030\,
            in1 => \N__18011\,
            in2 => \N__18024\,
            in3 => \N__36043\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38367\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18054\,
            in1 => \N__18063\,
            in2 => \_gnd_net_\,
            in3 => \N__32335\,
            lcout => \PCH_PWRGD.N_424\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIBP2A1_1_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__32336\,
            in1 => \_gnd_net_\,
            in2 => \N__18099\,
            in3 => \N__18057\,
            lcout => \PCH_PWRGD.N_278_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIBP2A1_0_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__18098\,
            in2 => \N__18174\,
            in3 => \N__32332\,
            lcout => \PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_0_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18082\,
            lcout => \PCH_PWRGD.N_413\,
            ltout => \PCH_PWRGD.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIBP2A1_0_0_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__18055\,
            in1 => \_gnd_net_\,
            in2 => \N__18033\,
            in3 => \N__32333\,
            lcout => \PCH_PWRGD.N_277_0\,
            ltout => \PCH_PWRGD.N_277_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI76R43_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__18020\,
            in1 => \N__18010\,
            in2 => \N__17991\,
            in3 => \N__36042\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.delayed_vccin_okZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17988\,
            in3 => \N__32334\,
            lcout => \N_227\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIFG4I5_0_10_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__29779\,
            in1 => \N__18228\,
            in2 => \N__18194\,
            in3 => \N__18244\,
            lcout => \PCH_PWRGD.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIFG4I5_10_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18227\,
            in1 => \_gnd_net_\,
            in2 => \N__18249\,
            in3 => \N__29777\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_10_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18245\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38396\,
            ce => \N__29897\,
            sr => \N__24296\
        );

    \PCH_PWRGD.count_1_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18137\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38396\,
            ce => \N__29897\,
            sr => \N__24296\
        );

    \PCH_PWRGD.count_12_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18218\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38396\,
            ce => \N__29897\,
            sr => \N__24296\
        );

    \PCH_PWRGD.count_RNIQRNC5_12_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18219\,
            in1 => \N__18204\,
            in2 => \_gnd_net_\,
            in3 => \N__29778\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI7H7A3_0_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__24295\,
            in1 => \N__18173\,
            in2 => \N__18150\,
            in3 => \N__32648\,
            lcout => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIMBB95_1_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18138\,
            in2 => \N__18126\,
            in3 => \N__18123\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19947\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_4_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19761\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19776\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19929\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19938\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21936\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29331\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18255\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__33185\,
            in1 => \_gnd_net_\,
            in2 => \N__19907\,
            in3 => \_gnd_net_\,
            lcout => \clk_100Khz_signalkeep_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__32211\,
            in1 => \N__19744\,
            in2 => \_gnd_net_\,
            in3 => \N__19691\,
            lcout => \RSMRST_PWRGD.N_423\,
            ltout => \RSMRST_PWRGD.N_423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18252\,
            in3 => \N__33184\,
            lcout => \RSMRST_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_1_fast_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19892\,
            in2 => \_gnd_net_\,
            in3 => \N__18488\,
            lcout => \clk_100Khz_signalkeep_4_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38413\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18300\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38515\,
            ce => \N__29874\,
            sr => \N__24353\
        );

    \PCH_PWRGD.count_14_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29927\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38515\,
            ce => \N__29874\,
            sr => \N__24353\
        );

    \POWERLED.count_off_5_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20144\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38522\,
            ce => \N__28086\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22013\,
            lcout => \POWERLED.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38522\,
            ce => \N__28086\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33148\,
            in1 => \N__18261\,
            in2 => \_gnd_net_\,
            in3 => \N__18327\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__32222\,
            in1 => \_gnd_net_\,
            in2 => \N__18267\,
            in3 => \N__19739\,
            lcout => \curr_state_RNIR5QD1_0_0\,
            ltout => \curr_state_RNIR5QD1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__19740\,
            in1 => \N__19682\,
            in2 => \N__18264\,
            in3 => \N__20509\,
            lcout => \RSMRST_PWRGD.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38489\,
            ce => \N__35999\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__20508\,
            in1 => \N__18341\,
            in2 => \N__19697\,
            in3 => \N__19741\,
            lcout => \RSMRST_PWRGD.curr_state_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38489\,
            ce => \N__35999\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__19743\,
            in1 => \N__19689\,
            in2 => \N__18544\,
            in3 => \N__20510\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.m4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18351\,
            in2 => \N__18345\,
            in3 => \N__33147\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__18342\,
            in1 => \N__19690\,
            in2 => \N__18330\,
            in3 => \N__20511\,
            lcout => \RSMRST_PWRGD.curr_state_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_fast_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__32221\,
            in1 => \_gnd_net_\,
            in2 => \N__19696\,
            in3 => \N__19742\,
            lcout => \RSMRST_PWRGD_RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38489\,
            ce => \N__35999\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIEP4G2_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__22054\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20660\,
            lcout => OPEN,
            ltout => \POWERLED.count_off_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIK80O8_0_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18438\,
            in2 => \N__18321\,
            in3 => \N__28044\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => \POWERLED.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18318\,
            in3 => \N__20008\,
            lcout => \POWERLED.count_off_RNIZ0Z_1\,
            ltout => \POWERLED.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIL90O8_1_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__20661\,
            in1 => \N__18306\,
            in2 => \N__18315\,
            in3 => \N__28043\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18312\,
            in2 => \_gnd_net_\,
            in3 => \N__20664\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => \N__28087\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFL179_3_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__20662\,
            in1 => \N__18444\,
            in2 => \N__28088\,
            in3 => \N__19982\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19983\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20665\,
            lcout => \POWERLED.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => \N__28087\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__20663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22053\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38575\,
            ce => \N__28087\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_2_1_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011111"
        )
    port map (
            in0 => \N__18811\,
            in1 => \N__23452\,
            in2 => \N__35432\,
            in3 => \N__18366\,
            lcout => \POWERLED.func_state_RNI3IN21_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0TA81_0_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18408\,
            in2 => \_gnd_net_\,
            in3 => \N__18810\,
            lcout => \POWERLED.N_425\,
            ltout => \POWERLED.N_425_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5F285_0_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__36044\,
            in1 => \N__18357\,
            in2 => \N__18372\,
            in3 => \N__22550\,
            lcout => \POWERLED.count_clk_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22750\,
            in2 => \_gnd_net_\,
            in3 => \N__18809\,
            lcout => \POWERLED.N_175\,
            ltout => \POWERLED.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_1_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18369\,
            in3 => \N__36742\,
            lcout => \POWERLED.un1_count_off_1_sqmuxa_8_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3F2B2_0_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111010"
        )
    port map (
            in0 => \N__32308\,
            in1 => \N__23422\,
            in2 => \N__19266\,
            in3 => \N__24945\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3P2F3_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__32997\,
            in1 => \N__32309\,
            in2 => \N__18360\,
            in3 => \N__20712\,
            lcout => \POWERLED.count_clk_en_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__19128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19253\,
            lcout => \POWERLED.dutycycle_1_0_iv_0_o3_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__18495\,
            in1 => \N__18461\,
            in2 => \N__18564\,
            in3 => \N__18666\,
            lcout => \POWERLED.func_state_RNI3IN21_1Z0Z_1\,
            ltout => \POWERLED.func_state_RNI3IN21_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIFJJH2_1_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__18588\,
            in1 => \N__18964\,
            in2 => \N__18657\,
            in3 => \N__36738\,
            lcout => \POWERLED.dutycycle_eena_3_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_sqmuxa_0_o2_x_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__19120\,
            in1 => \N__19233\,
            in2 => \N__33012\,
            in3 => \N__18654\,
            lcout => \POWERLED.func_state_0_sqmuxa_0_o2_xZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20592\,
            in2 => \_gnd_net_\,
            in3 => \N__22749\,
            lcout => \POWERLED.func_state_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g1_3_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__18548\,
            in1 => \N__18496\,
            in2 => \_gnd_net_\,
            in3 => \N__18462\,
            lcout => \POWERLED.g1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKBSM4_6_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111110000"
        )
    port map (
            in0 => \N__18993\,
            in1 => \N__18965\,
            in2 => \N__18720\,
            in3 => \N__29157\,
            lcout => \POWERLED.N_233_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18549\,
            in1 => \_gnd_net_\,
            in2 => \N__18500\,
            in3 => \N__18460\,
            lcout => rsmrstn,
            ltout => \rsmrstn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_0_6_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__19232\,
            in1 => \N__19119\,
            in2 => \N__18447\,
            in3 => \N__32998\,
            lcout => \POWERLED.N_388_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDUQ02_1_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001101"
        )
    port map (
            in0 => \N__19191\,
            in1 => \N__18729\,
            in2 => \N__19109\,
            in3 => \N__36727\,
            lcout => \POWERLED.un1_clk_100khz_42_and_i_o2_1_1\,
            ltout => \POWERLED.un1_clk_100khz_42_and_i_o2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIR58I4_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__18947\,
            in1 => \N__19410\,
            in2 => \N__18753\,
            in3 => \N__19326\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__19187\,
            in1 => \N__19081\,
            in2 => \_gnd_net_\,
            in3 => \N__18946\,
            lcout => \POWERLED.N_171\,
            ltout => \POWERLED.N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__19085\,
            in1 => \N__19192\,
            in2 => \N__18732\,
            in3 => \N__33141\,
            lcout => \POWERLED.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_0_1_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__19189\,
            in1 => \N__19083\,
            in2 => \N__33013\,
            in3 => \N__22748\,
            lcout => \POWERLED.N_387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_1_1_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__19084\,
            in1 => \N__19190\,
            in2 => \N__33014\,
            in3 => \N__25107\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_m1_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI98VE2_1_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__18966\,
            in1 => \N__23451\,
            in2 => \N__18723\,
            in3 => \N__36728\,
            lcout => \POWERLED.N_145_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3IN21_5_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__19082\,
            in1 => \N__19188\,
            in2 => \N__28971\,
            in3 => \N__18711\,
            lcout => \POWERLED.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNISHFV2_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111111111"
        )
    port map (
            in0 => \N__20589\,
            in1 => \N__22773\,
            in2 => \N__22808\,
            in3 => \N__22551\,
            lcout => \POWERLED.func_state_1_m2_am_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__19186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19034\,
            lcout => \POWERLED.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_0_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20588\,
            in1 => \N__19185\,
            in2 => \N__19050\,
            in3 => \N__32937\,
            lcout => \POWERLED.func_state_RNI8H551Z0Z_0\,
            ltout => \POWERLED.func_state_RNI8H551Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJK2D3_0_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18992\,
            in2 => \N__18981\,
            in3 => \N__18971\,
            lcout => \POWERLED.N_143_N\,
            ltout => \POWERLED.N_143_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIM6QF4_0_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18912\,
            in3 => \N__21024\,
            lcout => \POWERLED.N_116_f0\,
            ltout => \POWERLED.N_116_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_er_RNO_9_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100000000"
        )
    port map (
            in0 => \N__23692\,
            in1 => \_gnd_net_\,
            in2 => \N__18900\,
            in3 => \N__36053\,
            lcout => \POWERLED.dutycycle_en_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_er_9_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21002\,
            lcout => \POWERLED.dutycycle_erZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38577\,
            ce => \N__18885\,
            sr => \N__23337\
        );

    \POWERLED.func_state_RNI_2_0_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20587\,
            lcout => \POWERLED.N_3168_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIV0MP7_4_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__20882\,
            in1 => \N__23457\,
            in2 => \N__20760\,
            in3 => \N__20772\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26553\,
            in2 => \N__18756\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_7_a0_1_a1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_6_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__29151\,
            in1 => \N__21208\,
            in2 => \N__19314\,
            in3 => \N__19311\,
            lcout => \POWERLED.un1_dutycycle_53_7_a0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_7_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__21209\,
            in1 => \N__26555\,
            in2 => \N__23823\,
            in3 => \N__28589\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_13_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_13_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \N__25986\,
            in1 => \N__19290\,
            in2 => \N__19299\,
            in3 => \N__19296\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_12_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__26003\,
            in1 => \N__26554\,
            in2 => \N__28838\,
            in3 => \N__29152\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_0_0_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__19284\,
            in1 => \N__36758\,
            in2 => \_gnd_net_\,
            in3 => \N__23808\,
            lcout => \POWERLED.func_state_RNI8H551_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIANIR7_10_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__19482\,
            in1 => \N__23012\,
            in2 => \N__19467\,
            in3 => \N__26337\,
            lcout => \POWERLED.dutycycle_RNIANIR7Z0Z_10\,
            ltout => \POWERLED.dutycycle_RNIANIR7Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO3T79_10_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__19490\,
            in1 => \N__23454\,
            in2 => \N__19278\,
            in3 => \N__20984\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => \POWERLED.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_10_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19275\,
            in3 => \N__23148\,
            lcout => \POWERLED.un1_dutycycle_53_44_d_1_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNID3269_8_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__19433\,
            in1 => \N__19443\,
            in2 => \N__20838\,
            in3 => \N__23453\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => \POWERLED.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_10_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19503\,
            in3 => \N__26338\,
            lcout => \POWERLED.un1_dutycycle_53_44_d_1_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__19500\,
            in1 => \N__20985\,
            in2 => \N__19494\,
            in3 => \N__23455\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38619\,
            ce => 'H',
            sr => \N__23342\
        );

    \POWERLED.dutycycle_RNIANIR7_8_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__19481\,
            in1 => \N__23011\,
            in2 => \N__19466\,
            in3 => \N__23147\,
            lcout => \POWERLED.dutycycle_RNIANIR7Z0Z_8\,
            ltout => \POWERLED.dutycycle_RNIANIR7Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__20837\,
            in1 => \N__19434\,
            in2 => \N__19437\,
            in3 => \N__23456\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38619\,
            ce => 'H',
            sr => \N__23342\
        );

    \POWERLED.dutycycle_RNI_1_4_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000100010"
        )
    port map (
            in0 => \N__23799\,
            in1 => \N__28832\,
            in2 => \N__29156\,
            in3 => \N__26183\,
            lcout => \POWERLED.un1_dutycycle_53_39_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_3_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__23794\,
            in1 => \N__25828\,
            in2 => \N__28695\,
            in3 => \N__23164\,
            lcout => \POWERLED.dutycycle_RNI_10Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_1_0_LC_4_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__19409\,
            in1 => \N__19390\,
            in2 => \N__23807\,
            in3 => \N__19347\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_a2_6_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__23796\,
            in1 => \N__23168\,
            in2 => \N__26190\,
            in3 => \N__26356\,
            lcout => \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_6_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__25829\,
            in1 => \N__23795\,
            in2 => \_gnd_net_\,
            in3 => \N__29147\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_6\,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_8_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__26187\,
            in1 => \N__19563\,
            in2 => \N__19557\,
            in3 => \N__23170\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_10_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26355\,
            in1 => \N__29146\,
            in2 => \N__23202\,
            in3 => \N__28831\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_10\,
            ltout => \POWERLED.dutycycle_RNI_5Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_11_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__25844\,
            in1 => \N__25554\,
            in2 => \N__19554\,
            in3 => \N__23169\,
            lcout => \POWERLED.un1_dutycycle_53_44_d_c_1_s_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24057\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38133\,
            ce => \N__31953\,
            sr => \N__26806\
        );

    \VPP_VDDQ.count_2_14_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23978\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38133\,
            ce => \N__31953\,
            sr => \N__26806\
        );

    \VPP_VDDQ.count_2_4_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23910\,
            lcout => \VPP_VDDQ.count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38133\,
            ce => \N__31953\,
            sr => \N__26806\
        );

    \VPP_VDDQ.count_2_6_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23871\,
            lcout => \VPP_VDDQ.count_2_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38133\,
            ce => \N__31953\,
            sr => \N__26806\
        );

    \VPP_VDDQ.count_2_10_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24116\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38133\,
            ce => \N__31953\,
            sr => \N__26806\
        );

    \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19547\,
            in1 => \N__19518\,
            in2 => \N__30975\,
            in3 => \N__30924\,
            lcout => \N_392\,
            ltout => \N_392_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19752\,
            in2 => \N__19701\,
            in3 => \N__19698\,
            lcout => \RSMRSTn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38314\,
            ce => \N__35995\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI04B02_13_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__26790\,
            in1 => \N__31921\,
            in2 => \N__23745\,
            in3 => \N__24015\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => \VPP_VDDQ.count_2Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__31922\,
            in1 => \N__19584\,
            in2 => \N__19596\,
            in3 => \N__24056\,
            lcout => \VPP_VDDQ.un29_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI27C02_0_14_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__31830\,
            in1 => \N__21257\,
            in2 => \N__23982\,
            in3 => \N__31975\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un29_clk_100khz_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPT4L7_10_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19593\,
            in1 => \N__21483\,
            in2 => \N__19587\,
            in3 => \N__21222\,
            lcout => \VPP_VDDQ.un29_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU0A02_12_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31920\,
            in1 => \N__19583\,
            in2 => \_gnd_net_\,
            in3 => \N__24055\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011111100"
        )
    port map (
            in0 => \N__19815\,
            in1 => \N__27091\,
            in2 => \N__19802\,
            in3 => \N__26987\,
            lcout => OPEN,
            ltout => \HDA_STRAP.i4_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIT7P94_2_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19569\,
            in2 => \N__19575\,
            in3 => \N__33316\,
            lcout => \HDA_STRAP.curr_state_i_2\,
            ltout => \HDA_STRAP.curr_state_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100000011"
        )
    port map (
            in0 => \N__19817\,
            in1 => \N__27093\,
            in2 => \N__19572\,
            in3 => \N__26989\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38328\,
            ce => \N__35993\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__33322\,
            in1 => \N__19782\,
            in2 => \N__19803\,
            in3 => \N__19818\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNI_0_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27041\,
            in2 => \_gnd_net_\,
            in3 => \N__27129\,
            lcout => \HDA_STRAP.N_208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIS6P94_1_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__19824\,
            in1 => \N__27162\,
            in2 => \_gnd_net_\,
            in3 => \N__33315\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => \HDA_STRAP.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011111100"
        )
    port map (
            in0 => \N__27042\,
            in1 => \N__27092\,
            in2 => \N__19827\,
            in3 => \N__26988\,
            lcout => \HDA_STRAP.curr_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38328\,
            ce => \N__35993\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19816\,
            in2 => \_gnd_net_\,
            in3 => \N__19795\,
            lcout => \HDA_STRAP.HDA_SDO_ATP_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38328\,
            ce => \N__35993\,
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21569\,
            in1 => \N__21602\,
            in2 => \N__21588\,
            in3 => \N__21617\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21554\,
            in1 => \N__21521\,
            in2 => \N__21540\,
            in3 => \N__21758\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__21405\,
            in1 => \_gnd_net_\,
            in2 => \N__19906\,
            in3 => \N__21423\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21632\,
            in1 => \N__21286\,
            in2 => \N__21323\,
            in3 => \N__21469\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21287\,
            in1 => \N__19888\,
            in2 => \_gnd_net_\,
            in3 => \N__21273\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21441\,
            in1 => \N__21391\,
            in2 => \N__21362\,
            in3 => \N__21421\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21392\,
            in1 => \N__19886\,
            in2 => \_gnd_net_\,
            in3 => \N__21378\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19885\,
            in1 => \_gnd_net_\,
            in2 => \N__21477\,
            in3 => \N__21448\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21665\,
            in1 => \N__21650\,
            in2 => \N__21801\,
            in3 => \N__21680\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__19884\,
            in1 => \_gnd_net_\,
            in2 => \N__21449\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21695\,
            in1 => \N__21725\,
            in2 => \N__21744\,
            in3 => \N__21710\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19883\,
            in1 => \_gnd_net_\,
            in2 => \N__21339\,
            in3 => \N__21361\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__21300\,
            in1 => \N__19887\,
            in2 => \_gnd_net_\,
            in3 => \N__21322\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22064\,
            in2 => \N__20016\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNI515V2_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20668\,
            in1 => \N__20025\,
            in2 => \_gnd_net_\,
            in3 => \N__19986\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20174\,
            in2 => \_gnd_net_\,
            in3 => \N__19971\,
            lcout => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20073\,
            in3 => \N__19968\,
            lcout => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNI878V2_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20671\,
            in1 => \N__20130\,
            in2 => \_gnd_net_\,
            in3 => \N__19965\,
            lcout => \POWERLED.count_off_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNI999V2_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20669\,
            in1 => \N__21999\,
            in2 => \_gnd_net_\,
            in3 => \N__19962\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNIABAV2_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20672\,
            in1 => \_gnd_net_\,
            in2 => \N__27801\,
            in3 => \N__19959\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNIBDBV2_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20670\,
            in1 => \N__28155\,
            in2 => \_gnd_net_\,
            in3 => \N__19956\,
            lcout => \POWERLED.count_off_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNICFCV2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20673\,
            in1 => \_gnd_net_\,
            in2 => \N__21906\,
            in3 => \N__19953\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNIDHDV2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__20676\,
            in1 => \_gnd_net_\,
            in2 => \N__21888\,
            in3 => \N__19950\,
            lcout => \POWERLED.count_off_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNILNQT2_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20674\,
            in1 => \N__21857\,
            in2 => \_gnd_net_\,
            in3 => \N__20040\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNIMPRT2_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20677\,
            in1 => \N__21812\,
            in2 => \_gnd_net_\,
            in3 => \N__20037\,
            lcout => \POWERLED.count_off_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNINRST2_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20675\,
            in1 => \N__22079\,
            in2 => \_gnd_net_\,
            in3 => \N__20034\,
            lcout => \POWERLED.count_off_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNIOTTT2_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20678\,
            in1 => \N__22091\,
            in2 => \_gnd_net_\,
            in3 => \N__20031\,
            lcout => \POWERLED.count_off_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIPVUT2_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__22098\,
            in1 => \N__20679\,
            in2 => \_gnd_net_\,
            in3 => \N__20028\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNIPVUTZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21825\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38463\,
            ce => \N__28085\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20084\,
            in2 => \_gnd_net_\,
            in3 => \N__20667\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => \N__28099\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDI079_2_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20100\,
            in2 => \N__20115\,
            in3 => \N__28082\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => \POWERLED.count_offZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_1_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20009\,
            in1 => \N__20129\,
            in2 => \N__19989\,
            in3 => \N__21998\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_10_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22032\,
            in1 => \N__21894\,
            in2 => \N__20178\,
            in3 => \N__20157\,
            lcout => \POWERLED.count_off_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_3_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20069\,
            in1 => \N__27800\,
            in2 => \N__20175\,
            in3 => \N__28151\,
            lcout => \POWERLED.un34_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJR379_5_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28084\,
            in1 => \N__20151\,
            in2 => \_gnd_net_\,
            in3 => \N__20145\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20114\,
            lcout => \POWERLED.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38488\,
            ce => \N__28099\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHO279_4_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__20666\,
            in1 => \N__20094\,
            in2 => \N__20088\,
            in3 => \N__28083\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8FBJ_6_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__20055\,
            in1 => \N__25244\,
            in2 => \N__33381\,
            in3 => \N__22178\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38493\,
            ce => \N__25252\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIN1VB_10_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__22298\,
            in1 => \N__25246\,
            in2 => \N__20049\,
            in3 => \N__33348\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22299\,
            lcout => \POWERLED.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38493\,
            ce => \N__25252\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAICJ_7_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__20529\,
            in1 => \N__25245\,
            in2 => \N__33382\,
            in3 => \N__22166\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38493\,
            ce => \N__25252\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIAB7J1_0_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__20523\,
            in1 => \N__20374\,
            in2 => \_gnd_net_\,
            in3 => \N__20246\,
            lcout => \RSMRST_PWRGD.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI037J_2_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__25234\,
            in1 => \N__22199\,
            in2 => \N__20196\,
            in3 => \N__33323\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__25238\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2AHB_12_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__25236\,
            in1 => \N__22223\,
            in2 => \N__22212\,
            in3 => \N__33325\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI4DIB_13_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__20184\,
            in1 => \N__22241\,
            in2 => \N__33376\,
            in3 => \N__25237\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => \POWERLED.count_clkZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_10_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22287\,
            in1 => \N__22263\,
            in2 => \N__20187\,
            in3 => \N__22317\,
            lcout => \POWERLED.un2_count_clk_17_0_o2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22275\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__25238\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22242\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38588\,
            ce => \N__25238\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI07GB_11_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33324\,
            in1 => \N__22274\,
            in2 => \N__20739\,
            in3 => \N__25235\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__22736\,
            in1 => \N__20691\,
            in2 => \N__20706\,
            in3 => \N__20730\,
            lcout => \POWERLED.un1_func_state25_6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011011101"
        )
    port map (
            in0 => \N__20590\,
            in1 => \N__22606\,
            in2 => \_gnd_net_\,
            in3 => \N__22733\,
            lcout => \POWERLED.un1_func_state25_4_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__20823\,
            in1 => \N__24646\,
            in2 => \N__22617\,
            in3 => \N__25105\,
            lcout => \POWERLED.un1_func_state25_6_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI0TA81_7_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__24701\,
            in1 => \N__24684\,
            in2 => \N__24756\,
            in3 => \N__20697\,
            lcout => \POWERLED.count_clk_RNI0TA81Z0Z_7\,
            ltout => \POWERLED.count_clk_RNI0TA81Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIEP4G2_1_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__22734\,
            in1 => \N__22601\,
            in2 => \N__20682\,
            in3 => \N__20814\,
            lcout => \POWERLED.N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_7_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__24702\,
            in1 => \N__24685\,
            in2 => \_gnd_net_\,
            in3 => \N__24755\,
            lcout => OPEN,
            ltout => \POWERLED.N_431_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__22735\,
            in1 => \N__22825\,
            in2 => \N__20595\,
            in3 => \N__20591\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIESP71_0_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32816\,
            in1 => \N__20822\,
            in2 => \N__24648\,
            in3 => \N__22607\,
            lcout => \POWERLED.N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28649\,
            lcout => \POWERLED.un1_clk_100khz_43_and_i_0_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__23449\,
            in1 => \N__20793\,
            in2 => \N__20898\,
            in3 => \N__20799\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38594\,
            ce => 'H',
            sr => \N__23336\
        );

    \POWERLED.func_state_RNIFJJH2_0_1_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__24878\,
            in1 => \N__23448\,
            in2 => \N__23700\,
            in3 => \N__36732\,
            lcout => \POWERLED.un1_clk_100khz_40_and_i_0_0_0\,
            ltout => \POWERLED.un1_clk_100khz_40_and_i_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI41BF6_3_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__32631\,
            in1 => \N__20808\,
            in2 => \N__20802\,
            in3 => \N__22998\,
            lcout => \POWERLED.dutycycle_en_8\,
            ltout => \POWERLED.dutycycle_en_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITTKP7_3_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__20792\,
            in1 => \N__20894\,
            in2 => \N__20784\,
            in3 => \N__23447\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24876\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_40_and_i_0_d_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI41BF6_4_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__22999\,
            in1 => \N__20781\,
            in2 => \N__20775\,
            in3 => \N__32630\,
            lcout => \POWERLED.dutycycle_en_6\,
            ltout => \POWERLED.dutycycle_en_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__23450\,
            in1 => \N__20753\,
            in2 => \N__20763\,
            in3 => \N__20883\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38594\,
            ce => 'H',
            sr => \N__23336\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31376\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24999\,
            in2 => \N__36876\,
            in3 => \N__20919\,
            lcout => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36443\,
            in2 => \N__25019\,
            in3 => \N__20901\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNIZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25003\,
            in2 => \N__28650\,
            in3 => \N__20886\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25017\,
            in2 => \N__28794\,
            in3 => \N__20871\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__23529\,
            in1 => \N__25004\,
            in2 => \N__28970\,
            in3 => \N__20859\,
            lcout => \POWERLED.N_308\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29091\,
            in2 => \N__25018\,
            in3 => \N__20844\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24998\,
            in2 => \N__28569\,
            in3 => \N__20841\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25020\,
            in2 => \N__23172\,
            in3 => \N__20826\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNIECU31_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__23520\,
            in1 => \N__25005\,
            in2 => \N__26182\,
            in3 => \N__20988\,
            lcout => \POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25021\,
            in2 => \N__26367\,
            in3 => \N__20976\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__23521\,
            in1 => \N__25006\,
            in2 => \N__25528\,
            in3 => \N__20973\,
            lcout => \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HHZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__23522\,
            in1 => \N__25022\,
            in2 => \N__26539\,
            in3 => \N__20970\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25007\,
            in2 => \N__25981\,
            in3 => \N__20967\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25023\,
            in2 => \N__25751\,
            in3 => \N__20964\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__25929\,
            in1 => \N__25106\,
            in2 => \_gnd_net_\,
            in3 => \N__20961\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_6_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__26172\,
            in1 => \N__20957\,
            in2 => \N__21048\,
            in3 => \N__29142\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_10_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__26371\,
            in1 => \_gnd_net_\,
            in2 => \N__20937\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__28561\,
            in1 => \N__28674\,
            in2 => \_gnd_net_\,
            in3 => \N__28785\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_5_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__28786\,
            in1 => \N__28966\,
            in2 => \N__21051\,
            in3 => \N__23171\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_7_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26370\,
            lcout => \POWERLED.un1_dutycycle_53_axb_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011011000"
        )
    port map (
            in0 => \N__29144\,
            in1 => \N__22344\,
            in2 => \N__25860\,
            in3 => \N__26176\,
            lcout => \POWERLED.un1_i1_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__28562\,
            in1 => \N__29143\,
            in2 => \N__26188\,
            in3 => \N__28787\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_7_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__21039\,
            in1 => \N__21033\,
            in2 => \N__21027\,
            in3 => \N__23238\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_7_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28574\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3IN21_0_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__24935\,
            in1 => \N__23547\,
            in2 => \N__25848\,
            in3 => \N__36751\,
            lcout => \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__25752\,
            in1 => \_gnd_net_\,
            in2 => \N__25556\,
            in3 => \N__26357\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_10_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__26164\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21207\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_er_RNI_9_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26163\,
            lcout => \POWERLED.dutycycle_er_RNIZ0Z_9\,
            ltout => \POWERLED.dutycycle_er_RNIZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_4_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23797\,
            in2 => \N__21189\,
            in3 => \N__28795\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_4\,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_10_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__23798\,
            in1 => \N__26002\,
            in2 => \N__21162\,
            in3 => \N__21159\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_6Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_11_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011101111"
        )
    port map (
            in0 => \N__21153\,
            in1 => \N__21147\,
            in2 => \N__21141\,
            in3 => \N__21138\,
            lcout => \POWERLED.un1_dutycycle_53_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__36048\,
            in1 => \N__29213\,
            in2 => \N__21111\,
            in3 => \N__21131\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__21132\,
            in1 => \N__21110\,
            in2 => \N__29217\,
            in3 => \N__36049\,
            lcout => OPEN,
            ltout => \VPP_VDDQ_delayed_vddq_ok_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_PWRGD_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21096\,
            in3 => \N__27006\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_0_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21267\,
            in1 => \N__31913\,
            in2 => \_gnd_net_\,
            in3 => \N__23864\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__29193\,
            in1 => \N__26791\,
            in2 => \_gnd_net_\,
            in3 => \N__36047\,
            lcout => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__24117\,
            in1 => \N__21497\,
            in2 => \N__21261\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI27C02_14_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__31914\,
            in1 => \_gnd_net_\,
            in2 => \N__21258\,
            in3 => \N__23971\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__24138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26781\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38313\,
            ce => \N__31971\,
            sr => \N__26792\
        );

    \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21230\,
            in1 => \N__23842\,
            in2 => \_gnd_net_\,
            in3 => \N__31915\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38313\,
            ce => \N__31971\,
            sr => \N__26792\
        );

    \VPP_VDDQ.count_2_RNIASDQ1_9_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__26776\,
            in1 => \N__24137\,
            in2 => \N__21243\,
            in3 => \N__31916\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => \VPP_VDDQ.count_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__31918\,
            in1 => \N__23844\,
            in2 => \N__21234\,
            in3 => \N__21231\,
            lcout => \VPP_VDDQ.un29_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__24081\,
            in1 => \_gnd_net_\,
            in2 => \N__26814\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38313\,
            ce => \N__31971\,
            sr => \N__26792\
        );

    \VPP_VDDQ.count_2_RNIST802_11_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__31917\,
            in1 => \N__26777\,
            in2 => \N__21507\,
            in3 => \N__24080\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => \VPP_VDDQ.count_2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__21498\,
            in1 => \N__24115\,
            in2 => \N__21486\,
            in3 => \N__31919\,
            lcout => \VPP_VDDQ.un29_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21476\,
            in2 => \N__21453\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21422\,
            in2 => \_gnd_net_\,
            in3 => \N__21399\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21396\,
            in2 => \_gnd_net_\,
            in3 => \N__21366\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21363\,
            in2 => \_gnd_net_\,
            in3 => \N__21327\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21324\,
            in2 => \_gnd_net_\,
            in3 => \N__21291\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21288\,
            in2 => \_gnd_net_\,
            in3 => \N__21636\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21633\,
            in2 => \_gnd_net_\,
            in3 => \N__21621\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__38321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21618\,
            in2 => \_gnd_net_\,
            in3 => \N__21606\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__38321\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21603\,
            in2 => \_gnd_net_\,
            in3 => \N__21591\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21587\,
            in2 => \_gnd_net_\,
            in3 => \N__21573\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21570\,
            in2 => \_gnd_net_\,
            in3 => \N__21558\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21555\,
            in2 => \_gnd_net_\,
            in3 => \N__21543\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21539\,
            in2 => \_gnd_net_\,
            in3 => \N__21525\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21522\,
            in2 => \_gnd_net_\,
            in3 => \N__21510\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21759\,
            in2 => \_gnd_net_\,
            in3 => \N__21747\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21743\,
            in2 => \_gnd_net_\,
            in3 => \N__21729\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__38315\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21726\,
            in2 => \_gnd_net_\,
            in3 => \N__21714\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21711\,
            in2 => \_gnd_net_\,
            in3 => \N__21699\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21696\,
            in2 => \_gnd_net_\,
            in3 => \N__21684\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21681\,
            in2 => \_gnd_net_\,
            in3 => \N__21669\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21666\,
            in2 => \_gnd_net_\,
            in3 => \N__21654\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21651\,
            in2 => \_gnd_net_\,
            in3 => \N__21639\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21800\,
            in2 => \_gnd_net_\,
            in3 => \N__21786\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21948\,
            in2 => \_gnd_net_\,
            in3 => \N__21783\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__38340\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21959\,
            in2 => \_gnd_net_\,
            in3 => \N__21780\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21984\,
            in3 => \N__21777\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21972\,
            in3 => \N__21774\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29345\,
            in2 => \_gnd_net_\,
            in3 => \N__21771\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29384\,
            in2 => \_gnd_net_\,
            in3 => \N__21768\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29363\,
            in2 => \_gnd_net_\,
            in3 => \N__21765\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29402\,
            in2 => \_gnd_net_\,
            in3 => \N__21762\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38262\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21980\,
            in1 => \N__21968\,
            in2 => \N__21960\,
            in3 => \N__21947\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21915\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38123\,
            ce => \N__28107\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIR7879_9_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21921\,
            in1 => \N__21914\,
            in2 => \_gnd_net_\,
            in3 => \N__28103\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => \POWERLED.count_offZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_10_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21813\,
            in1 => \N__21887\,
            in2 => \N__21897\,
            in3 => \N__21858\,
            lcout => \POWERLED.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI4ID59_10_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21864\,
            in1 => \N__28104\,
            in2 => \_gnd_net_\,
            in3 => \N__21872\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21873\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38123\,
            ce => \N__28107\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDPQ39_11_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21837\,
            in1 => \N__28105\,
            in2 => \_gnd_net_\,
            in3 => \N__21845\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38123\,
            ce => \N__28107\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIFSR39_12_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21831\,
            in1 => \N__28106\,
            in2 => \_gnd_net_\,
            in3 => \N__21824\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22112\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38263\,
            ce => \N__28080\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHVS39_13_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28069\,
            in1 => \N__22137\,
            in2 => \_gnd_net_\,
            in3 => \N__22145\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22149\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38263\,
            ce => \N__28080\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJ2U39_14_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28070\,
            in1 => \N__22119\,
            in2 => \_gnd_net_\,
            in3 => \N__22127\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22131\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38263\,
            ce => \N__28080\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIL5V39_15_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22113\,
            in1 => \N__22104\,
            in2 => \_gnd_net_\,
            in3 => \N__28081\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => \POWERLED.count_offZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22092\,
            in1 => \N__22080\,
            in2 => \N__22068\,
            in3 => \N__22065\,
            lcout => \POWERLED.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILU479_6_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28068\,
            in1 => \N__22026\,
            in2 => \_gnd_net_\,
            in3 => \N__22014\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25426\,
            in2 => \N__24808\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25386\,
            in1 => \N__22438\,
            in2 => \_gnd_net_\,
            in3 => \N__22191\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25390\,
            in1 => \N__22383\,
            in2 => \_gnd_net_\,
            in3 => \N__22188\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25387\,
            in1 => \_gnd_net_\,
            in2 => \N__24550\,
            in3 => \N__22185\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25391\,
            in1 => \_gnd_net_\,
            in2 => \N__24602\,
            in3 => \N__22182\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25388\,
            in1 => \N__22418\,
            in2 => \_gnd_net_\,
            in3 => \N__22170\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25392\,
            in1 => \N__24667\,
            in2 => \_gnd_net_\,
            in3 => \N__22158\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25389\,
            in1 => \N__22458\,
            in2 => \_gnd_net_\,
            in3 => \N__22155\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25393\,
            in1 => \N__24728\,
            in2 => \_gnd_net_\,
            in3 => \N__22152\,
            lcout => \POWERLED.count_clk_1_9\,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__25397\,
            in1 => \_gnd_net_\,
            in2 => \N__22316\,
            in3 => \N__22290\,
            lcout => \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9\,
            carryout => \POWERLED.un1_count_clk_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25394\,
            in1 => \N__22286\,
            in2 => \_gnd_net_\,
            in3 => \N__22266\,
            lcout => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10\,
            carryout => \POWERLED.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25398\,
            in1 => \N__22262\,
            in2 => \_gnd_net_\,
            in3 => \N__22251\,
            lcout => \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11\,
            carryout => \POWERLED.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25395\,
            in1 => \N__22248\,
            in2 => \_gnd_net_\,
            in3 => \N__22233\,
            lcout => \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12\,
            carryout => \POWERLED.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25399\,
            in1 => \N__24470\,
            in2 => \_gnd_net_\,
            in3 => \N__22230\,
            lcout => \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__25396\,
            in1 => \N__24513\,
            in2 => \_gnd_net_\,
            in3 => \N__22227\,
            lcout => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22224\,
            lcout => \POWERLED.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38309\,
            ce => \N__25302\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_2_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__22457\,
            in1 => \N__22381\,
            in2 => \N__22467\,
            in3 => \N__22439\,
            lcout => \POWERLED.N_385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38421\,
            ce => \N__25285\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_4_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24551\,
            in1 => \N__22424\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNICLDJ_8_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33363\,
            in1 => \N__22364\,
            in2 => \N__22353\,
            in3 => \N__25284\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => \POWERLED.count_clkZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_2_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__24552\,
            in1 => \N__22382\,
            in2 => \N__22443\,
            in3 => \N__22440\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_6_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__22425\,
            in1 => \N__24740\,
            in2 => \N__22407\,
            in3 => \N__24687\,
            lcout => \POWERLED.count_clk_RNIZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI268J_3_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__25283\,
            in1 => \N__22403\,
            in2 => \N__22392\,
            in3 => \N__33362\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22365\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38421\,
            ce => \N__25285\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__28856\,
            in1 => \N__23208\,
            in2 => \_gnd_net_\,
            in3 => \N__28631\,
            lcout => \POWERLED.un1_N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_3_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__28632\,
            in1 => \N__31419\,
            in2 => \N__28869\,
            in3 => \N__36630\,
            lcout => \POWERLED.g3_0_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__31418\,
            in1 => \_gnd_net_\,
            in2 => \N__28868\,
            in3 => \N__36859\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_1_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__32976\,
            in1 => \N__35513\,
            in2 => \N__22616\,
            in3 => \N__24647\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_1_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__36678\,
            in1 => \N__22826\,
            in2 => \N__22782\,
            in3 => \N__22751\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI43L44_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22779\,
            in1 => \N__22772\,
            in2 => \N__22755\,
            in3 => \N__22533\,
            lcout => \POWERLED.func_state_RNI43L44_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22752\,
            in2 => \_gnd_net_\,
            in3 => \N__22602\,
            lcout => \POWERLED.func_state_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__22475\,
            in1 => \N__22497\,
            in2 => \N__22491\,
            in3 => \N__23537\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38564\,
            ce => 'H',
            sr => \N__23341\
        );

    \POWERLED.dutycycle_RNI28MU5_7_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111111111"
        )
    port map (
            in0 => \N__23535\,
            in1 => \N__23022\,
            in2 => \N__28573\,
            in3 => \N__23686\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_5_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIB8FGC_7_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__23684\,
            in1 => \N__32638\,
            in2 => \N__22512\,
            in3 => \N__22509\,
            lcout => \POWERLED.dutycycle_RNIB8FGCZ0Z_7\,
            ltout => \POWERLED.dutycycle_RNIB8FGCZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNICHTQD_7_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__23538\,
            in1 => \N__22487\,
            in2 => \N__22479\,
            in3 => \N__22476\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1BA98_14_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__23527\,
            in1 => \N__22925\,
            in2 => \N__22959\,
            in3 => \N__22946\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM6QF4_14_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23528\,
            in2 => \N__22965\,
            in3 => \N__23021\,
            lcout => OPEN,
            ltout => \POWERLED.N_158_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI41BF6_14_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__23685\,
            in1 => \N__24948\,
            in2 => \N__22962\,
            in3 => \N__32639\,
            lcout => \POWERLED.dutycycle_en_11\,
            ltout => \POWERLED.dutycycle_en_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__23536\,
            in1 => \N__22935\,
            in2 => \N__22950\,
            in3 => \N__22947\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38564\,
            ce => 'H',
            sr => \N__23341\
        );

    \POWERLED.dutycycle_11_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__22890\,
            in1 => \N__22901\,
            in2 => \N__22914\,
            in3 => \N__32647\,
            lcout => \POWERLED.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38612\,
            ce => 'H',
            sr => \N__23335\
        );

    \POWERLED.dutycycle_RNI8D4S4_11_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__32645\,
            in1 => \N__22910\,
            in2 => \N__22902\,
            in3 => \N__22889\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => \POWERLED.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_11_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22878\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__32646\,
            in1 => \N__22875\,
            in2 => \N__22851\,
            in3 => \N__22866\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38612\,
            ce => 'H',
            sr => \N__23335\
        );

    \POWERLED.dutycycle_RNIAG5S4_12_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__22874\,
            in1 => \N__22865\,
            in2 => \N__32649\,
            in3 => \N__22847\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => \POWERLED.dutycycleZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25527\,
            in2 => \N__23100\,
            in3 => \N__25916\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_6_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100001111"
        )
    port map (
            in0 => \N__23097\,
            in1 => \N__23091\,
            in2 => \N__23079\,
            in3 => \N__23076\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23070\,
            in3 => \N__25917\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIV7998_13_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__23523\,
            in1 => \N__23036\,
            in2 => \N__23061\,
            in3 => \N__23048\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => \POWERLED.dutycycleZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM6QF4_13_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23524\,
            in2 => \N__23067\,
            in3 => \N__23013\,
            lcout => OPEN,
            ltout => \POWERLED.N_156_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI41BF6_13_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__23698\,
            in1 => \N__24946\,
            in2 => \N__23064\,
            in3 => \N__32643\,
            lcout => \POWERLED.dutycycle_en_10\,
            ltout => \POWERLED.dutycycle_en_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__23534\,
            in1 => \N__23037\,
            in2 => \N__23052\,
            in3 => \N__23049\,
            lcout => \POWERLED.dutycycleZ1Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__23343\
        );

    \POWERLED.dutycycle_RNI3EB98_15_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__23351\,
            in1 => \N__23533\,
            in2 => \N__23565\,
            in3 => \N__23555\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => \POWERLED.dutycycleZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM6QF4_15_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23525\,
            in2 => \N__23025\,
            in3 => \N__23014\,
            lcout => OPEN,
            ltout => \POWERLED.N_161_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI41BF6_15_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__23699\,
            in1 => \N__24947\,
            in2 => \N__23568\,
            in3 => \N__32644\,
            lcout => \POWERLED.dutycycle_en_12\,
            ltout => \POWERLED.dutycycle_en_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__23556\,
            in1 => \N__23526\,
            in2 => \N__23355\,
            in3 => \N__23352\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38613\,
            ce => 'H',
            sr => \N__23343\
        );

    \POWERLED.dutycycle_RNI_3_6_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29141\,
            in1 => \N__23790\,
            in2 => \N__26470\,
            in3 => \N__25852\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_8_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__23791\,
            in1 => \N__23211\,
            in2 => \N__25862\,
            in3 => \N__28863\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_49_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_10_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__26453\,
            in1 => \N__23231\,
            in2 => \N__23241\,
            in3 => \N__26392\,
            lcout => \POWERLED.un1_dutycycle_53_49_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__26393\,
            in1 => \N__25970\,
            in2 => \N__26471\,
            in3 => \N__26559\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_8_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__23220\,
            in1 => \N__23232\,
            in2 => \N__23223\,
            in3 => \N__26178\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_8_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011111111"
        )
    port map (
            in0 => \N__23793\,
            in1 => \N__23213\,
            in2 => \N__28866\,
            in3 => \N__26454\,
            lcout => \POWERLED.un1_dutycycle_53_2_1_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__23212\,
            in1 => \N__23792\,
            in2 => \N__26567\,
            in3 => \N__26391\,
            lcout => \POWERLED.un1_dutycycle_53_axb_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_3_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28694\,
            in2 => \N__23806\,
            in3 => \N__28864\,
            lcout => \POWERLED.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__26803\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24014\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37881\,
            ce => \N__31977\,
            sr => \N__26805\
        );

    \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31887\,
            in1 => \_gnd_net_\,
            in2 => \N__23906\,
            in3 => \N__23730\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => \VPP_VDDQ.count_2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26932\,
            in1 => \N__23940\,
            in2 => \N__23721\,
            in3 => \N__23883\,
            lcout => \VPP_VDDQ.un29_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINUSC_0_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32765\,
            in1 => \N__26930\,
            in2 => \_gnd_net_\,
            in3 => \N__26801\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIC4UI1_0_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__26907\,
            in1 => \_gnd_net_\,
            in2 => \N__23718\,
            in3 => \N__31886\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINUSC_1_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23939\,
            in2 => \N__23715\,
            in3 => \N__26802\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID5UI1_1_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23706\,
            in2 => \N__23712\,
            in3 => \N__31885\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => \VPP_VDDQ.count_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26931\,
            in2 => \N__23709\,
            in3 => \N__26804\,
            lcout => \VPP_VDDQ.count_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37881\,
            ce => \N__31977\,
            sr => \N__26805\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23938\,
            in2 => \N__26934\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26270\,
            in2 => \_gnd_net_\,
            in3 => \N__23922\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26236\,
            in2 => \_gnd_net_\,
            in3 => \N__23919\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26783\,
            in1 => \N__23916\,
            in2 => \_gnd_net_\,
            in3 => \N__23889\,
            lcout => \VPP_VDDQ.count_2_rst_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26581\,
            in2 => \_gnd_net_\,
            in3 => \N__23886\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26784\,
            in1 => \N__23882\,
            in2 => \_gnd_net_\,
            in3 => \N__23853\,
            lcout => \VPP_VDDQ.count_2_rst_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26775\,
            in1 => \N__23850\,
            in2 => \_gnd_net_\,
            in3 => \N__23829\,
            lcout => \VPP_VDDQ.count_2_rst_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26850\,
            in3 => \N__23826\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24144\,
            in2 => \_gnd_net_\,
            in3 => \N__24129\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26795\,
            in1 => \N__24126\,
            in2 => \_gnd_net_\,
            in3 => \N__24090\,
            lcout => \VPP_VDDQ.count_2_rst_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24087\,
            in2 => \_gnd_net_\,
            in3 => \N__24072\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26793\,
            in1 => \N__24069\,
            in2 => \_gnd_net_\,
            in3 => \N__24030\,
            lcout => \VPP_VDDQ.count_2_rst_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24027\,
            in2 => \_gnd_net_\,
            in3 => \N__23994\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26794\,
            in1 => \N__23991\,
            in2 => \_gnd_net_\,
            in3 => \N__23946\,
            lcout => \VPP_VDDQ.count_2_rst_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31826\,
            in1 => \N__26796\,
            in2 => \_gnd_net_\,
            in3 => \N__23943\,
            lcout => \VPP_VDDQ.count_2_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32003\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37968\,
            ce => \N__31965\,
            sr => \N__26800\
        );

    \POWERLED.count_4_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29696\,
            lcout => \POWERLED.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38260\,
            ce => \N__35992\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27276\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38260\,
            ce => \N__35992\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI5S8O_15_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24168\,
            in1 => \N__33310\,
            in2 => \_gnd_net_\,
            in3 => \N__27323\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27327\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38075\,
            ce => \N__35988\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI7UKN_7_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24162\,
            in1 => \_gnd_net_\,
            in2 => \N__27261\,
            in3 => \N__33311\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27260\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38075\,
            ce => \N__35988\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI91MN_8_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24156\,
            in1 => \N__33313\,
            in2 => \_gnd_net_\,
            in3 => \N__27242\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27246\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38075\,
            ce => \N__35988\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIB4NN_9_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24150\,
            in1 => \N__33312\,
            in2 => \_gnd_net_\,
            in3 => \N__27227\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27231\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38075\,
            ce => \N__35988\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI1M6O_13_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33289\,
            in1 => \N__24423\,
            in2 => \_gnd_net_\,
            in3 => \N__27357\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_13_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27356\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38261\,
            ce => \N__35991\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__33286\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24417\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI3OIN_5_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24189\,
            in1 => \N__33288\,
            in2 => \_gnd_net_\,
            in3 => \N__27287\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27291\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38261\,
            ce => \N__35991\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI3P7O_14_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27342\,
            in1 => \N__24183\,
            in2 => \_gnd_net_\,
            in3 => \N__33290\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27341\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38261\,
            ce => \N__35991\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI5RJN_6_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24177\,
            in1 => \N__33287\,
            in2 => \_gnd_net_\,
            in3 => \N__27275\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNITF4O_11_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27213\,
            in1 => \N__24441\,
            in2 => \_gnd_net_\,
            in3 => \N__33292\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27212\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38122\,
            ce => \N__35990\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIVHGN_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24435\,
            in2 => \N__27183\,
            in3 => \N__33291\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27182\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38122\,
            ce => \N__35990\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIVI5O_12_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27369\,
            in1 => \N__24429\,
            in2 => \_gnd_net_\,
            in3 => \N__33293\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27368\,
            lcout => \POWERLED.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38122\,
            ce => \N__35990\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__25442\,
            in1 => \_gnd_net_\,
            in2 => \N__25404\,
            in3 => \N__24810\,
            lcout => \POWERLED.count_clk_RNIZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25441\,
            in2 => \_gnd_net_\,
            in3 => \N__25400\,
            lcout => \POWERLED.count_clk_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29272\,
            in2 => \_gnd_net_\,
            in3 => \N__36202\,
            lcout => \VPP_VDDQ.N_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27759\,
            lcout => \POWERLED.mult1_un103_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27488\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27659\,
            lcout => \POWERLED.un85_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30045\,
            lcout => \POWERLED.un85_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI499J_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33284\,
            in1 => \N__24519\,
            in2 => \N__24531\,
            in3 => \N__25303\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24530\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38076\,
            ce => \N__25295\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24480\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38076\,
            ce => \N__25295\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8JKB_15_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__24447\,
            in1 => \N__33285\,
            in2 => \N__25311\,
            in3 => \N__24459\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => \POWERLED.count_clkZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_15_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24471\,
            in1 => \N__24501\,
            in2 => \N__24489\,
            in3 => \N__25425\,
            lcout => \POWERLED.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI6GJB_14_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25304\,
            in1 => \N__24486\,
            in2 => \N__33359\,
            in3 => \N__24479\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24458\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38076\,
            ce => \N__25295\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI9LLG_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__25308\,
            in1 => \N__25320\,
            in2 => \N__33358\,
            in3 => \N__24765\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__24729\,
            in1 => \N__24801\,
            in2 => \N__24603\,
            in3 => \N__24713\,
            lcout => \POWERLED.N_193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24612\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38308\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIEOEJ_9_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__33361\,
            in1 => \N__24573\,
            in2 => \N__25279\,
            in3 => \N__24581\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => \POWERLED.count_clkZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_5_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__24714\,
            in1 => \_gnd_net_\,
            in2 => \N__24705\,
            in3 => \N__24598\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24700\,
            in1 => \N__24686\,
            in2 => \N__24651\,
            in3 => \N__24800\,
            lcout => \POWERLED.count_clk_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI6CAJ_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__24618\,
            in1 => \N__25254\,
            in2 => \N__33388\,
            in3 => \N__24611\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24582\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38308\,
            ce => \N__25310\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAMLG_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__24774\,
            in1 => \N__33360\,
            in2 => \N__24567\,
            in3 => \N__25253\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27828\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24821\,
            in2 => \N__33885\,
            in3 => \N__24843\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27714\,
            in2 => \N__24825\,
            in3 => \N__24840\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27705\,
            in2 => \N__30738\,
            in3 => \N__24837\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27696\,
            in2 => \N__30737\,
            in3 => \N__24834\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__33707\,
            in1 => \N__24820\,
            in2 => \N__27687\,
            in3 => \N__24831\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27675\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24828\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30730\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000101000"
        )
    port map (
            in0 => \N__25379\,
            in1 => \N__24809\,
            in2 => \N__25443\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38420\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25437\,
            in2 => \_gnd_net_\,
            in3 => \N__25380\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38420\,
            ce => \N__25309\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNI_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27072\,
            lcout => \HDA_STRAP.N_3252_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_6_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25138\,
            lcout => \POWERLED.N_203_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25118\,
            lcout => \POWERLED.N_175_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24936\,
            lcout => \POWERLED.func_state_RNI_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27924\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27614\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28689\,
            in2 => \N__31417\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31400\,
            in2 => \N__24855\,
            in3 => \N__24846\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36464\,
            in2 => \N__28884\,
            in3 => \N__25614\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26199\,
            in2 => \N__36475\,
            in3 => \N__25611\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28983\,
            in2 => \N__28485\,
            in3 => \N__25608\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25605\,
            in2 => \N__28969\,
            in3 => \N__25593\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28959\,
            in2 => \N__25590\,
            in3 => \N__25578\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26397\,
            in2 => \N__25575\,
            in3 => \N__25560\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25543\,
            in2 => \N__25485\,
            in3 => \N__25467\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26538\,
            in2 => \N__25464\,
            in3 => \N__25446\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25973\,
            in2 => \N__26070\,
            in3 => \N__25689\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25747\,
            in2 => \N__26031\,
            in3 => \N__25686\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25918\,
            in2 => \N__25683\,
            in3 => \N__25674\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25671\,
            in2 => \N__25982\,
            in3 => \N__25662\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26049\,
            in2 => \N__25760\,
            in3 => \N__25659\,
            lcout => \POWERLED.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26019\,
            in2 => \N__25930\,
            in3 => \N__25656\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25695\,
            in2 => \N__25931\,
            in3 => \N__25653\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25650\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100101101"
        )
    port map (
            in0 => \N__36879\,
            in1 => \N__25647\,
            in2 => \N__28353\,
            in3 => \N__28855\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_2_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26202\,
            in3 => \N__36463\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__25977\,
            in1 => \N__26189\,
            in2 => \N__26085\,
            in3 => \N__26396\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27923\,
            in2 => \N__27951\,
            in3 => \N__27895\,
            lcout => \POWERLED.mult1_un40_sum_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \N__25758\,
            in1 => \N__26289\,
            in2 => \N__26061\,
            in3 => \N__25971\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26040\,
            in2 => \_gnd_net_\,
            in3 => \N__25753\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__25925\,
            in1 => \_gnd_net_\,
            in2 => \N__25707\,
            in3 => \N__25754\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_13_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__26010\,
            in1 => \N__25972\,
            in2 => \N__25932\,
            in3 => \N__25874\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_a2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_14_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25856\,
            in2 => \N__25785\,
            in3 => \N__25759\,
            lcout => \POWERLED.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25761\,
            in3 => \N__25706\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26560\,
            in2 => \N__26477\,
            in3 => \N__26395\,
            lcout => \POWERLED.un1_m2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS66Q1_2_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26249\,
            in1 => \N__26280\,
            in2 => \_gnd_net_\,
            in3 => \N__31923\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_2\,
            ltout => \VPP_VDDQ.un1_count_2_1_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__32758\,
            in1 => \N__26258\,
            in2 => \N__26283\,
            in3 => \N__26807\,
            lcout => \VPP_VDDQ.count_2_rst_6\,
            ltout => \VPP_VDDQ.count_2_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__26250\,
            in1 => \N__26238\,
            in2 => \N__26274\,
            in3 => \N__31925\,
            lcout => \VPP_VDDQ.un29_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__26271\,
            in1 => \N__26259\,
            in2 => \N__32776\,
            in3 => \N__26812\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37883\,
            ce => \N__31936\,
            sr => \N__26813\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__26222\,
            in1 => \N__26237\,
            in2 => \N__26817\,
            in3 => \N__32759\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU97Q1_3_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31924\,
            in1 => \_gnd_net_\,
            in2 => \N__26241\,
            in3 => \N__26208\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => \VPP_VDDQ.count_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__26223\,
            in1 => \N__26816\,
            in2 => \N__26211\,
            in3 => \N__32764\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37883\,
            ce => \N__31936\,
            sr => \N__26813\
        );

    \VPP_VDDQ.count_2_0_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32760\,
            in1 => \N__26933\,
            in2 => \_gnd_net_\,
            in3 => \N__26811\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__37883\,
            ce => \N__31936\,
            sr => \N__26813\
        );

    \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31964\,
            in1 => \N__26898\,
            in2 => \_gnd_net_\,
            in3 => \N__26604\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => \VPP_VDDQ.count_2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__26828\,
            in1 => \N__32768\,
            in2 => \N__26901\,
            in3 => \N__26785\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38354\,
            ce => \N__31969\,
            sr => \N__26782\
        );

    \VPP_VDDQ.count_2_5_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__26582\,
            in1 => \N__32769\,
            in2 => \N__26815\,
            in3 => \N__26891\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38354\,
            ce => \N__31969\,
            sr => \N__26782\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__26892\,
            in1 => \N__26583\,
            in2 => \N__32777\,
            in3 => \N__26789\,
            lcout => \VPP_VDDQ.count_2_rst_3\,
            ltout => \VPP_VDDQ.count_2_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__31970\,
            in1 => \N__26597\,
            in2 => \N__26883\,
            in3 => \N__26845\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un29_clk_100khz_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINKK9B_2_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26880\,
            in1 => \N__26868\,
            in2 => \N__26859\,
            in3 => \N__26856\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => \VPP_VDDQ.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__26849\,
            in1 => \N__26829\,
            in2 => \N__26820\,
            in3 => \N__26763\,
            lcout => \VPP_VDDQ.count_2_rst_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26598\,
            in1 => \N__26589\,
            in2 => \_gnd_net_\,
            in3 => \N__31963\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIR99J4_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__26940\,
            in1 => \N__27153\,
            in2 => \_gnd_net_\,
            in3 => \N__33314\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => \HDA_STRAP.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m8_i_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111001100"
        )
    port map (
            in0 => \N__27004\,
            in1 => \N__27090\,
            in2 => \N__27165\,
            in3 => \N__27065\,
            lcout => \HDA_STRAP.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m6_i_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__38712\,
            in1 => \_gnd_net_\,
            in2 => \N__26955\,
            in3 => \N__26964\,
            lcout => \HDA_STRAP.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_en_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26950\,
            in2 => \_gnd_net_\,
            in3 => \N__36045\,
            lcout => \HDA_STRAP.count_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27033\,
            in2 => \_gnd_net_\,
            in3 => \N__27125\,
            lcout => \N_414\,
            ltout => \N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27096\,
            in3 => \N__38710\,
            lcout => \HDA_STRAP.N_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010011011"
        )
    port map (
            in0 => \N__27064\,
            in1 => \N__27034\,
            in2 => \N__27018\,
            in3 => \N__27003\,
            lcout => \HDA_STRAP.m6_i_0\,
            ltout => \HDA_STRAP.m6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38711\,
            in2 => \N__26958\,
            in3 => \N__26951\,
            lcout => \HDA_STRAP.curr_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38457\,
            ce => \N__35998\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_2_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__30370\,
            in1 => \_gnd_net_\,
            in2 => \N__30340\,
            in3 => \N__30297\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_5_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__30227\,
            in1 => \N__30190\,
            in2 => \N__27201\,
            in3 => \N__30260\,
            lcout => \POWERLED.un79_clk_100khzlto15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__33386\,
            in1 => \_gnd_net_\,
            in2 => \N__32118\,
            in3 => \N__32075\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_15_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30479\,
            in1 => \N__27315\,
            in2 => \_gnd_net_\,
            in3 => \N__30430\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_8_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__30127\,
            in1 => \N__30622\,
            in2 => \N__27198\,
            in3 => \N__27195\,
            lcout => \POWERLED.count_RNIZ0Z_8\,
            ltout => \POWERLED.count_RNIZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIHU1M_0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__32116\,
            in1 => \N__36052\,
            in2 => \N__27189\,
            in3 => \N__33387\,
            lcout => \POWERLED.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30003\,
            in2 => \N__30404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIB209_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29646\,
            in1 => \N__30371\,
            in2 => \_gnd_net_\,
            in3 => \N__27186\,
            lcout => \POWERLED.count_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIC419_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29649\,
            in1 => \N__30341\,
            in2 => \_gnd_net_\,
            in3 => \N__27168\,
            lcout => \POWERLED.count_1_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2\,
            carryout => \POWERLED.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNID629_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29645\,
            in1 => \N__30295\,
            in2 => \_gnd_net_\,
            in3 => \N__27294\,
            lcout => \POWERLED.count_1_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3\,
            carryout => \POWERLED.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNIE839_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29650\,
            in1 => \N__30256\,
            in2 => \_gnd_net_\,
            in3 => \N__27279\,
            lcout => \POWERLED.count_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNIFA49_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29647\,
            in1 => \N__30223\,
            in2 => \_gnd_net_\,
            in3 => \N__27264\,
            lcout => \POWERLED.count_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIGC59_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29651\,
            in1 => \N__30191\,
            in2 => \_gnd_net_\,
            in3 => \N__27249\,
            lcout => \POWERLED.count_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIHE69_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29648\,
            in1 => \N__30128\,
            in2 => \_gnd_net_\,
            in3 => \N__27234\,
            lcout => \POWERLED.count_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNIIG79_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29652\,
            in1 => \N__30623\,
            in2 => \_gnd_net_\,
            in3 => \N__27219\,
            lcout => \POWERLED.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNIJI89_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__29657\,
            in1 => \_gnd_net_\,
            in2 => \N__30596\,
            in3 => \N__27216\,
            lcout => \POWERLED.count_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__29653\,
            in1 => \_gnd_net_\,
            in2 => \N__30563\,
            in3 => \N__27204\,
            lcout => \POWERLED.count_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNISEH7_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29655\,
            in1 => \N__30530\,
            in2 => \_gnd_net_\,
            in3 => \N__27360\,
            lcout => \POWERLED.count_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNITGI7_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29654\,
            in1 => \N__30503\,
            in2 => \_gnd_net_\,
            in3 => \N__27345\,
            lcout => \POWERLED.count_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29656\,
            in1 => \N__30475\,
            in2 => \_gnd_net_\,
            in3 => \N__27333\,
            lcout => \POWERLED.count_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__30437\,
            in1 => \N__29658\,
            in2 => \_gnd_net_\,
            in3 => \N__27330\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30502\,
            in1 => \N__30529\,
            in2 => \N__30595\,
            in3 => \N__30556\,
            lcout => \POWERLED.un79_clk_100khzlto15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_1_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100001010"
        )
    port map (
            in0 => \N__32456\,
            in1 => \N__34274\,
            in2 => \N__32412\,
            in3 => \N__32495\,
            lcout => \DSW_PWRGD.curr_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38486\,
            ce => \N__36002\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_7_1_0__m6_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011100"
        )
    port map (
            in0 => \N__34272\,
            in1 => \N__32458\,
            in2 => \N__32502\,
            in3 => \N__32398\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.curr_state_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNIMJ7I_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33330\,
            in1 => \_gnd_net_\,
            in2 => \N__27306\,
            in3 => \N__27303\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_1\,
            ltout => \DSW_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010100000"
        )
    port map (
            in0 => \N__34273\,
            in1 => \N__32455\,
            in2 => \N__27297\,
            in3 => \N__32403\,
            lcout => \DSW_PWRGD.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38486\,
            ce => \N__36002\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_7_1_0__m4_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010100000"
        )
    port map (
            in0 => \N__32457\,
            in1 => \N__34271\,
            in2 => \N__32413\,
            in3 => \N__32496\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNILI7I_0_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27405\,
            in2 => \N__27399\,
            in3 => \N__33329\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_0\,
            ltout => \DSW_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNIIJFC_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33331\,
            in1 => \N__32459\,
            in2 => \N__27396\,
            in3 => \N__32493\,
            lcout => \DSW_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.DSW_PWROK_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__32494\,
            in1 => \N__32454\,
            in2 => \_gnd_net_\,
            in3 => \N__32402\,
            lcout => \DSW_PWRGD.DSW_PWROK_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38486\,
            ce => \N__36002\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33827\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27502\,
            in2 => \N__27393\,
            in3 => \N__27381\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27456\,
            in2 => \N__27507\,
            in3 => \N__27378\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27655\,
            in2 => \N__27447\,
            in3 => \N__27375\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27435\,
            in2 => \N__27660\,
            in3 => \N__27372\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30044\,
            in1 => \N__27506\,
            in2 => \N__27426\,
            in3 => \N__27513\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27414\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27510\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27654\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27492\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_9_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27628\,
            in2 => \N__27471\,
            in3 => \N__27450\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2_c\,
            carryout => \POWERLED.mult1_un110_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27597\,
            in2 => \N__27633\,
            in3 => \N__27438\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3_c\,
            carryout => \POWERLED.mult1_un110_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27751\,
            in2 => \N__27582\,
            in3 => \N__27429\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4_c\,
            carryout => \POWERLED.mult1_un110_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27561\,
            in2 => \N__27758\,
            in3 => \N__27417\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5_c\,
            carryout => \POWERLED.mult1_un110_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__27653\,
            in1 => \N__27632\,
            in2 => \N__27546\,
            in3 => \N__27408\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6_c\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27522\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27663\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27750\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27618\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27724\,
            in2 => \N__27813\,
            in3 => \N__27591\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27588\,
            in2 => \N__27729\,
            in3 => \N__27573\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33708\,
            in2 => \N__27570\,
            in3 => \N__27555\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27552\,
            in2 => \N__33716\,
            in3 => \N__27537\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__27749\,
            in1 => \N__27728\,
            in2 => \N__27534\,
            in3 => \N__27516\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__27768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27762\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33712\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33902\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33642\,
            in2 => \N__27866\,
            in3 => \N__27708\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27862\,
            in2 => \N__30675\,
            in3 => \N__27699\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30822\,
            in2 => \N__30663\,
            in3 => \N__27690\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30651\,
            in2 => \N__30828\,
            in3 => \N__27678\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30729\,
            in1 => \N__30852\,
            in2 => \N__27867\,
            in3 => \N__27669\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30843\,
            in3 => \N__27666\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30821\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31005\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27849\,
            in3 => \N__27840\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27879\,
            in3 => \N__27837\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28291\,
            in2 => \N__27933\,
            in3 => \N__27834\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27831\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27827\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__28327\,
            in1 => \N__28328\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIN1679_7_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__28042\,
            in1 => \N__28161\,
            in2 => \_gnd_net_\,
            in3 => \N__28178\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38614\,
            ce => \N__28089\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIP4779_8_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__28131\,
            in1 => \_gnd_net_\,
            in2 => \N__28116\,
            in3 => \N__28041\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28130\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38614\,
            ce => \N__28089\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000101"
        )
    port map (
            in0 => \N__27922\,
            in1 => \_gnd_net_\,
            in2 => \N__27900\,
            in3 => \N__27950\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27921\,
            in2 => \_gnd_net_\,
            in3 => \N__27896\,
            lcout => \POWERLED.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28238\,
            in2 => \_gnd_net_\,
            in3 => \N__28250\,
            lcout => \POWERLED.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30884\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30984\,
            in3 => \N__27870\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28344\,
            in2 => \N__28335\,
            in3 => \N__28311\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28292\,
            in2 => \N__28308\,
            in3 => \N__28296\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28293\,
            in2 => \N__28272\,
            in3 => \N__28260\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28406\,
            in1 => \N__28218\,
            in2 => \N__28203\,
            in3 => \N__28257\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28254\,
            in2 => \N__28239\,
            in3 => \N__28221\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__28216\,
            in1 => \N__28217\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28364\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30867\,
            in2 => \N__28385\,
            in3 => \N__28194\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28381\,
            in2 => \N__28191\,
            in3 => \N__28182\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28402\,
            in2 => \N__28449\,
            in3 => \N__28440\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28437\,
            in2 => \N__28407\,
            in3 => \N__28431\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31465\,
            in1 => \N__28428\,
            in2 => \N__28386\,
            in3 => \N__28422\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28419\,
            in3 => \N__28410\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28401\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36866\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28368\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__28675\,
            in1 => \N__36468\,
            in2 => \_gnd_net_\,
            in3 => \N__29122\,
            lcout => \POWERLED.un1_dutycycle_53_axb_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__36863\,
            in1 => \N__28676\,
            in2 => \_gnd_net_\,
            in3 => \N__29124\,
            lcout => \POWERLED.d_i3_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_3_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__28677\,
            in1 => \N__29123\,
            in2 => \N__28865\,
            in3 => \N__36864\,
            lcout => OPEN,
            ltout => \POWERLED.un1_i3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_5_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__28478\,
            in1 => \N__28968\,
            in2 => \N__28992\,
            in3 => \N__28989\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__28967\,
            in1 => \N__36865\,
            in2 => \N__36476\,
            in3 => \N__28846\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28847\,
            in1 => \N__28678\,
            in2 => \_gnd_net_\,
            in3 => \N__28587\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28458\,
            in1 => \N__29289\,
            in2 => \_gnd_net_\,
            in3 => \N__33374\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28464\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_3140_i\,
            ltout => \VPP_VDDQ.N_3140_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__32767\,
            in1 => \N__29207\,
            in2 => \N__28461\,
            in3 => \N__33622\,
            lcout => \VPP_VDDQ.m4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__29273\,
            in1 => \N__29282\,
            in2 => \_gnd_net_\,
            in3 => \N__29437\,
            lcout => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0\,
            ltout => \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__29178\,
            in1 => \N__33602\,
            in2 => \N__28452\,
            in3 => \N__33375\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__29206\,
            in1 => \N__32766\,
            in2 => \N__29319\,
            in3 => \N__29303\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38206\,
            ce => \N__35989\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__29283\,
            in1 => \_gnd_net_\,
            in2 => \N__29444\,
            in3 => \N__29274\,
            lcout => \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_1_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__33603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29192\,
            lcout => \VPP_VDDQ.curr_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38206\,
            ce => \N__35989\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_6_c_RNI2H3S_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__34964\,
            in1 => \N__31577\,
            in2 => \N__31610\,
            in3 => \N__34297\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIU43Q1_7_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34725\,
            in1 => \_gnd_net_\,
            in2 => \N__29172\,
            in3 => \N__31482\,
            lcout => \DSW_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIQU0Q1_5_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29471\,
            in1 => \N__34724\,
            in2 => \_gnd_net_\,
            in3 => \N__29166\,
            lcout => \DSW_PWRGD.un2_count_1_axb_5\,
            ltout => \DSW_PWRGD.un2_count_1_axb_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_4_c_RNI0D1S_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__34296\,
            in1 => \N__31643\,
            in2 => \N__29169\,
            in3 => \N__34963\,
            lcout => \DSW_PWRGD.count_rst_9\,
            ltout => \DSW_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIQU0Q1_0_5_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__29472\,
            in1 => \N__34727\,
            in2 => \N__29160\,
            in3 => \N__31602\,
            lcout => \DSW_PWRGD.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_5_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__31658\,
            in1 => \N__31644\,
            in2 => \N__34315\,
            in3 => \N__35014\,
            lcout => \DSW_PWRGD.count_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38355\,
            ce => \N__34733\,
            sr => \N__35013\
        );

    \DSW_PWRGD.un2_count_1_cry_9_c_RNI5N6S_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__34965\,
            in1 => \N__34298\,
            in2 => \N__31802\,
            in3 => \N__31769\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIBAB22_10_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34726\,
            in1 => \_gnd_net_\,
            in2 => \N__29463\,
            in3 => \N__29541\,
            lcout => \DSW_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33626\,
            lcout => \VPP_VDDQ.N_3160_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_1_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34542\,
            lcout => \DSW_PWRGD.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38182\,
            ce => \N__34729\,
            sr => \N__34968\
        );

    \DSW_PWRGD.un2_count_1_cry_7_c_RNI3J4S_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31553\,
            in1 => \N__34966\,
            in2 => \N__31539\,
            in3 => \N__34269\,
            lcout => \DSW_PWRGD.count_rst_6\,
            ltout => \DSW_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNI084Q1_0_8_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__34708\,
            in1 => \N__29559\,
            in2 => \N__29421\,
            in3 => \N__31800\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.un12_clk_100khz_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNI227D7_2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34194\,
            in1 => \N__31278\,
            in2 => \N__29418\,
            in3 => \N__29415\,
            lcout => \DSW_PWRGD.un12_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29406\,
            in1 => \N__29388\,
            in2 => \N__29370\,
            in3 => \N__29349\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNI084Q1_8_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29558\,
            in1 => \N__34707\,
            in2 => \_gnd_net_\,
            in3 => \N__29568\,
            lcout => \DSW_PWRGD.un2_count_1_axb_8\,
            ltout => \DSW_PWRGD.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_8_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__34270\,
            in1 => \N__34980\,
            in2 => \N__29562\,
            in3 => \N__31538\,
            lcout => \DSW_PWRGD.count_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38359\,
            ce => \N__34734\,
            sr => \N__34981\
        );

    \DSW_PWRGD.count_RNIHLBVB_4_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34755\,
            in1 => \N__29550\,
            in2 => \N__34386\,
            in3 => \N__34449\,
            lcout => \DSW_PWRGD.N_1_i\,
            ltout => \DSW_PWRGD.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_10_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__34967\,
            in1 => \N__31801\,
            in2 => \N__29544\,
            in3 => \N__31770\,
            lcout => \DSW_PWRGD.count_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38359\,
            ce => \N__34734\,
            sr => \N__34981\
        );

    \POWERLED.curr_state_RNI2PKG_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36054\,
            in2 => \_gnd_net_\,
            in3 => \N__32111\,
            lcout => \POWERLED.g0_i_o3_0\,
            ltout => \POWERLED.g0_i_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101110"
        )
    port map (
            in0 => \N__29507\,
            in1 => \N__32047\,
            in2 => \N__29532\,
            in3 => \N__29516\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38456\,
            ce => 'H',
            sr => \N__29529\
        );

    \POWERLED.pwm_out_RNIEHDM1_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010100"
        )
    port map (
            in0 => \N__29517\,
            in1 => \N__29508\,
            in2 => \N__32054\,
            in3 => \N__29499\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__32112\,
            in1 => \N__32074\,
            in2 => \_gnd_net_\,
            in3 => \N__32046\,
            lcout => OPEN,
            ltout => \POWERLED.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI3P6L_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32019\,
            in2 => \N__29475\,
            in3 => \N__33300\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => \POWERLED.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIF5D5_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__33301\,
            in1 => \_gnd_net_\,
            in2 => \N__29682\,
            in3 => \N__32073\,
            lcout => \POWERLED.count_0_sqmuxa_i\,
            ltout => \POWERLED.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__30004\,
            in1 => \_gnd_net_\,
            in2 => \N__29679\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGAFE_0_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33302\,
            in1 => \_gnd_net_\,
            in2 => \N__29676\,
            in3 => \N__29592\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__29661\,
            in1 => \N__30400\,
            in2 => \_gnd_net_\,
            in3 => \N__29998\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIHBFE_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29667\,
            in2 => \N__29673\,
            in3 => \N__33377\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => \POWERLED.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30002\,
            in2 => \N__29670\,
            in3 => \N__29659\,
            lcout => \POWERLED.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38352\,
            ce => \N__35996\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__29660\,
            in1 => \_gnd_net_\,
            in2 => \N__30008\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38352\,
            ce => \N__35996\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIKKSP_10_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33379\,
            in1 => \_gnd_net_\,
            in2 => \N__29586\,
            in3 => \N__29574\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29582\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38352\,
            ce => \N__35996\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNITEFN_2_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33378\,
            in1 => \N__29955\,
            in2 => \_gnd_net_\,
            in3 => \N__29963\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29967\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38352\,
            ce => \N__35996\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIS12Q1_6_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29949\,
            in1 => \N__34706\,
            in2 => \_gnd_net_\,
            in3 => \N__31628\,
            lcout => \DSW_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_6_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.count_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38487\,
            ce => \N__34728\,
            sr => \N__34937\
        );

    \HDA_STRAP.count_RNID9AT_4_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37771\,
            in1 => \N__33858\,
            in2 => \_gnd_net_\,
            in3 => \N__33981\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIF61V_14_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33873\,
            in1 => \N__34041\,
            in2 => \_gnd_net_\,
            in3 => \N__37770\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIJIDT_7_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37772\,
            in1 => \N__33843\,
            in2 => \_gnd_net_\,
            in3 => \N__33951\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIU1QC5_14_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29943\,
            in1 => \N__29931\,
            in2 => \_gnd_net_\,
            in3 => \N__29895\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI1LHN_4_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29709\,
            in1 => \N__33380\,
            in2 => \_gnd_net_\,
            in3 => \N__29697\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33764\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30019\,
            in2 => \N__33804\,
            in3 => \N__30105\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30102\,
            in2 => \N__30024\,
            in3 => \N__30096\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30047\,
            in2 => \N__30093\,
            in3 => \N__30084\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30081\,
            in2 => \N__30051\,
            in3 => \N__30075\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__33484\,
            in1 => \N__30023\,
            in2 => \N__30072\,
            in3 => \N__30063\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__30060\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30054\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30046\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30009\,
            in1 => \N__29973\,
            in2 => \N__31296\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33675\,
            in2 => \N__30381\,
            in3 => \N__30405\,
            lcout => \POWERLED.N_6478_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30372\,
            in1 => \N__30348\,
            in2 => \N__33921\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6479_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36489\,
            in2 => \N__30306\,
            in3 => \N__30342\,
            lcout => \POWERLED.N_6480_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30296\,
            in1 => \N__30270\,
            in2 => \N__33738\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6481_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30264\,
            in1 => \N__30237\,
            in2 => \N__33417\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6482_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30231\,
            in1 => \N__30204\,
            in2 => \N__32796\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6483_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30198\,
            in1 => \N__30159\,
            in2 => \N__30174\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6484_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30111\,
            in2 => \N__30153\,
            in3 => \N__30138\,
            lcout => \POWERLED.N_6485_i\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30642\,
            in2 => \N__30606\,
            in3 => \N__30630\,
            lcout => \POWERLED.N_6486_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30597\,
            in1 => \N__30573\,
            in2 => \N__33687\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_6487_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30543\,
            in2 => \N__30705\,
            in3 => \N__30567\,
            lcout => \POWERLED.N_6488_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30516\,
            in2 => \N__30684\,
            in3 => \N__30537\,
            lcout => \POWERLED.N_6489_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30690\,
            in2 => \N__30489\,
            in3 => \N__30510\,
            lcout => \POWERLED.N_6490_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30696\,
            in2 => \N__30453\,
            in3 => \N__30480\,
            lcout => \POWERLED.N_6491_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30861\,
            in2 => \N__30414\,
            in3 => \N__30444\,
            lcout => \POWERLED.N_6492_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30741\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30728\,
            lcout => \POWERLED.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31124\,
            lcout => \POWERLED.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31074\,
            lcout => \POWERLED.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30827\,
            lcout => \POWERLED.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33659\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31029\,
            in2 => \N__30800\,
            in3 => \N__30666\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30796\,
            in2 => \N__30783\,
            in3 => \N__30654\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31065\,
            in2 => \N__30771\,
            in3 => \N__30645\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30759\,
            in2 => \N__31073\,
            in3 => \N__30846\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__30826\,
            in1 => \N__30750\,
            in2 => \N__30801\,
            in3 => \N__30834\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31089\,
            in3 => \N__30831\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31064\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31043\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31266\,
            in2 => \N__31022\,
            in3 => \N__30774\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31018\,
            in2 => \N__31236\,
            in3 => \N__30762\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31212\,
            in2 => \N__31125\,
            in3 => \N__30753\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31123\,
            in2 => \N__31191\,
            in3 => \N__30744\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31069\,
            in1 => \N__31170\,
            in2 => \N__31023\,
            in3 => \N__31080\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31152\,
            in3 => \N__31077\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31110\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31004\,
            lcout => \POWERLED.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30952\,
            in2 => \_gnd_net_\,
            in3 => \N__30911\,
            lcout => v1p8a_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30885\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31466\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31259\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31260\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31242\,
            in2 => \N__31439\,
            in3 => \N__31224\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31435\,
            in2 => \N__31221\,
            in3 => \N__31203\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31461\,
            in2 => \N__31200\,
            in3 => \N__31179\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31176\,
            in2 => \N__31467\,
            in3 => \N__31161\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31111\,
            in1 => \N__31158\,
            in2 => \N__31440\,
            in3 => \N__31140\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31137\,
            in3 => \N__31128\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31460\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31420\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31309\,
            in2 => \N__31326\,
            in3 => \N__37087\,
            lcout => \G_3119\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36603\,
            in2 => \N__31314\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37088\,
            in2 => \N__37197\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37167\,
            in2 => \N__37092\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31313\,
            in2 => \N__37143\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37116\,
            in2 => \_gnd_net_\,
            in3 => \N__31299\,
            lcout => \POWERLED.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIKLTP1_0_2_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__34683\,
            in1 => \N__31515\,
            in2 => \N__31694\,
            in3 => \N__31503\,
            lcout => \DSW_PWRGD.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_1_c_RNIT6UR_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__31706\,
            in1 => \N__31719\,
            in2 => \N__34316\,
            in3 => \N__34955\,
            lcout => \DSW_PWRGD.count_rst_12\,
            ltout => \DSW_PWRGD.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIKLTP1_2_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34681\,
            in1 => \_gnd_net_\,
            in2 => \N__31509\,
            in3 => \N__31502\,
            lcout => \DSW_PWRGD.un2_count_1_axb_2\,
            ltout => \DSW_PWRGD.un2_count_1_axb_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_2_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31707\,
            in1 => \N__34314\,
            in2 => \N__31506\,
            in3 => \N__34956\,
            lcout => \DSW_PWRGD.count_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38366\,
            ce => \N__34722\,
            sr => \N__35023\
        );

    \DSW_PWRGD.un2_count_1_cry_2_c_RNIU8VR_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__34312\,
            in1 => \N__31673\,
            in2 => \N__31695\,
            in3 => \N__34958\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIMOUP1_3_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31488\,
            in2 => \N__31494\,
            in3 => \N__34682\,
            lcout => \DSW_PWRGD.countZ0Z_3\,
            ltout => \DSW_PWRGD.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_3_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__34313\,
            in1 => \N__31674\,
            in2 => \N__31491\,
            in3 => \N__34959\,
            lcout => \DSW_PWRGD.count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38366\,
            ce => \N__34722\,
            sr => \N__35023\
        );

    \DSW_PWRGD.count_7_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__31611\,
            in1 => \N__31578\,
            in2 => \N__34317\,
            in3 => \N__34957\,
            lcout => \DSW_PWRGD.count_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38366\,
            ce => \N__34722\,
            sr => \N__35023\
        );

    \DSW_PWRGD.un2_count_1_cry_0_c_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34062\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \DSW_PWRGD.un2_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_0_c_RNIS4TR_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35015\,
            in1 => \N__34517\,
            in2 => \_gnd_net_\,
            in3 => \N__31470\,
            lcout => \DSW_PWRGD.count_rst_13\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_0\,
            carryout => \DSW_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_1_THRU_LUT4_0_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31718\,
            in2 => \_gnd_net_\,
            in3 => \N__31698\,
            lcout => \DSW_PWRGD.un2_count_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_1\,
            carryout => \DSW_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31687\,
            in2 => \_gnd_net_\,
            in3 => \N__31665\,
            lcout => \DSW_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_2\,
            carryout => \DSW_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_3_c_RNIVA0S_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35016\,
            in1 => \N__34437\,
            in2 => \_gnd_net_\,
            in3 => \N__31662\,
            lcout => \DSW_PWRGD.count_rst_10\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_3\,
            carryout => \DSW_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31659\,
            in2 => \_gnd_net_\,
            in3 => \N__31632\,
            lcout => \DSW_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_4\,
            carryout => \DSW_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_5_c_RNI1F2S_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35017\,
            in1 => \N__34406\,
            in2 => \_gnd_net_\,
            in3 => \N__31614\,
            lcout => \DSW_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_5\,
            carryout => \DSW_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31606\,
            in2 => \_gnd_net_\,
            in3 => \N__31560\,
            lcout => \DSW_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_6\,
            carryout => \DSW_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31557\,
            in2 => \_gnd_net_\,
            in3 => \N__31521\,
            lcout => \DSW_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \DSW_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_8_c_RNI4L5S_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35018\,
            in1 => \N__34182\,
            in2 => \_gnd_net_\,
            in3 => \N__31518\,
            lcout => \DSW_PWRGD.count_rst_5\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_8\,
            carryout => \DSW_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31803\,
            in2 => \_gnd_net_\,
            in3 => \N__31749\,
            lcout => \DSW_PWRGD.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_9\,
            carryout => \DSW_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34335\,
            in3 => \N__31746\,
            lcout => \DSW_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_10\,
            carryout => \DSW_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_11_c_RNIEJ0P_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35020\,
            in1 => \N__34479\,
            in2 => \_gnd_net_\,
            in3 => \N__31743\,
            lcout => \DSW_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_11\,
            carryout => \DSW_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_12_c_RNIFL1P_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35019\,
            in1 => \N__34766\,
            in2 => \_gnd_net_\,
            in3 => \N__31740\,
            lcout => \DSW_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_12\,
            carryout => \DSW_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_13_c_RNIGN2P_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__35022\,
            in1 => \N__34782\,
            in2 => \_gnd_net_\,
            in3 => \N__31737\,
            lcout => \DSW_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un2_count_1_cry_13\,
            carryout => \DSW_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_14_c_RNIHP3P_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34806\,
            in1 => \N__35021\,
            in2 => \_gnd_net_\,
            in3 => \N__31734\,
            lcout => \DSW_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_15_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35129\,
            in1 => \N__35655\,
            in2 => \N__35175\,
            in3 => \N__35628\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un13_clk_100khz_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIU55T1_11_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__32151\,
            in1 => \N__35688\,
            in2 => \N__31731\,
            in3 => \N__31725\,
            lcout => \VPP_VDDQ.un13_clk_100khz_i\,
            ltout => \VPP_VDDQ.un13_clk_100khz_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__35128\,
            in1 => \_gnd_net_\,
            in2 => \N__31728\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__35901\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_3_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35067\,
            in1 => \N__35357\,
            in2 => \N__35085\,
            in3 => \N__35099\,
            lcout => \VPP_VDDQ.un13_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNINRAO_0_11_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__35333\,
            in1 => \N__35204\,
            in2 => \N__35309\,
            in3 => \N__35144\,
            lcout => \VPP_VDDQ.un13_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_0_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35127\,
            in2 => \_gnd_net_\,
            in3 => \N__35255\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI513Q_0_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32145\,
            in2 => \N__32139\,
            in3 => \N__35877\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => \VPP_VDDQ.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_1_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__35145\,
            in1 => \_gnd_net_\,
            in2 => \N__32136\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38441\,
            ce => \N__35901\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI623Q_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32133\,
            in1 => \N__32124\,
            in2 => \_gnd_net_\,
            in3 => \N__35878\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => \VPP_VDDQ.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__35123\,
            in1 => \_gnd_net_\,
            in2 => \N__32127\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32117\,
            in2 => \N__32085\,
            in3 => \N__32055\,
            lcout => \POWERLED.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38445\,
            ce => \N__35997\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI4AD02_15_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32010\,
            in1 => \N__31992\,
            in2 => \_gnd_net_\,
            in3 => \N__31976\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI95OO_12_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35571\,
            in1 => \N__35583\,
            in2 => \_gnd_net_\,
            in3 => \N__35879\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI9DR41_3_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35880\,
            in1 => \N__35547\,
            in2 => \_gnd_net_\,
            in3 => \N__35558\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIB8PO_13_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35601\,
            in1 => \N__35589\,
            in2 => \_gnd_net_\,
            in3 => \N__35881\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIBGS41_4_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__35882\,
            in1 => \N__35537\,
            in2 => \_gnd_net_\,
            in3 => \N__35523\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIDBQO_14_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32169\,
            in1 => \N__35640\,
            in2 => \_gnd_net_\,
            in3 => \N__35885\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_14_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38449\,
            ce => \N__35897\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIDJT41_5_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32163\,
            in1 => \N__35051\,
            in2 => \_gnd_net_\,
            in3 => \N__35884\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_5_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38449\,
            ce => \N__35897\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFERO_15_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32157\,
            in1 => \N__35609\,
            in2 => \_gnd_net_\,
            in3 => \N__35886\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_15_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35610\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38449\,
            ce => \N__35897\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFMU41_6_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35373\,
            in1 => \N__32712\,
            in2 => \_gnd_net_\,
            in3 => \N__35883\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_6_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35372\,
            lcout => \VPP_VDDQ.count_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38449\,
            ce => \N__35897\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.DSW_PWROK_RNIH6QL_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32706\,
            in1 => \_gnd_net_\,
            in2 => \N__33389\,
            in3 => \N__32379\,
            lcout => dsw_pwrok,
            ltout => \dsw_pwrok_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__32679\,
            in1 => \_gnd_net_\,
            in2 => \N__32667\,
            in3 => \N__32175\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNI57NN_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__32414\,
            in1 => \N__32500\,
            in2 => \N__32469\,
            in3 => \N__32635\,
            lcout => \DSW_PWRGD.curr_state_RNI57NNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNI3E27_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__32501\,
            in1 => \N__32465\,
            in2 => \_gnd_net_\,
            in3 => \N__32415\,
            lcout => \DSW_PWRGD.curr_state_RNI3E27Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32373\,
            in1 => \N__32358\,
            in2 => \N__32346\,
            in3 => \N__32226\,
            lcout => \VCCIN_PWRGD.un10_outputZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI67MK_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__35256\,
            in1 => \N__36075\,
            in2 => \N__33399\,
            in3 => \N__33369\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => \VPP_VDDQ.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__33036\,
            in1 => \N__36117\,
            in2 => \N__33402\,
            in3 => \N__35257\,
            lcout => \VPP_VDDQ.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38548\,
            ce => \N__36000\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNO_0_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36090\,
            in2 => \_gnd_net_\,
            in3 => \N__33370\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIUHA31_10_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35277\,
            in1 => \N__33030\,
            in2 => \_gnd_net_\,
            in3 => \N__35819\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_10_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35276\,
            lcout => \VPP_VDDQ.count_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38547\,
            ce => \N__35876\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32928\,
            in2 => \_gnd_net_\,
            in3 => \N__32892\,
            lcout => \POWERLED.N_388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33560\,
            lcout => \POWERLED.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33497\,
            lcout => \POWERLED.un85_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33500\,
            in2 => \_gnd_net_\,
            in3 => \N__33455\,
            lcout => \POWERLED.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32778\,
            in2 => \_gnd_net_\,
            in3 => \N__33633\,
            lcout => \VPP_VDDQ.m4_0_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33789\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33744\,
            in2 => \N__33585\,
            in3 => \N__33576\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33573\,
            in2 => \N__33567\,
            in3 => \N__33543\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33506\,
            in2 => \N__33540\,
            in3 => \N__33525\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33522\,
            in2 => \N__33510\,
            in3 => \N__33471\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36282\,
            in1 => \N__33468\,
            in2 => \N__33462\,
            in3 => \N__33438\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33435\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33423\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => \POWERLED.mult1_un131_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33420\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33828\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33768\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35672\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33720\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36569\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37076\,
            lcout => \POWERLED.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33663\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37053\,
            lcout => \POWERLED.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33906\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__36248\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34040\,
            lcout => \HDA_STRAP.count_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__37695\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33974\,
            lcout => \HDA_STRAP.count_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__37695\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33947\,
            lcout => \HDA_STRAP.count_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__37695\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37367\,
            lcout => \HDA_STRAP.count_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__37695\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34002\,
            lcout => \HDA_STRAP.count_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38623\,
            ce => \N__37695\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_1_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37347\,
            in2 => \N__37488\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \HDA_STRAP.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37614\,
            in2 => \_gnd_net_\,
            in3 => \N__33987\,
            lcout => \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_1\,
            carryout => \HDA_STRAP.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37017\,
            in2 => \_gnd_net_\,
            in3 => \N__33984\,
            lcout => \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_2\,
            carryout => \HDA_STRAP.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37010\,
            in2 => \_gnd_net_\,
            in3 => \N__33960\,
            lcout => \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_3\,
            carryout => \HDA_STRAP.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37416\,
            in2 => \_gnd_net_\,
            in3 => \N__33957\,
            lcout => \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_4\,
            carryout => \HDA_STRAP.un2_count_1_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38701\,
            in1 => \N__34149\,
            in2 => \_gnd_net_\,
            in3 => \N__33954\,
            lcout => \HDA_STRAP.count_1_6\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_5_cZ0\,
            carryout => \HDA_STRAP.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37250\,
            in2 => \_gnd_net_\,
            in3 => \N__33933\,
            lcout => \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_6\,
            carryout => \HDA_STRAP.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38702\,
            in1 => \N__37638\,
            in2 => \_gnd_net_\,
            in3 => \N__33930\,
            lcout => \HDA_STRAP.count_1_8\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_7\,
            carryout => \HDA_STRAP.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37224\,
            in2 => \_gnd_net_\,
            in3 => \N__33927\,
            lcout => \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \HDA_STRAP.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38690\,
            in1 => \N__37532\,
            in2 => \_gnd_net_\,
            in3 => \N__33924\,
            lcout => \HDA_STRAP.count_1_10\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_9\,
            carryout => \HDA_STRAP.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38692\,
            in1 => \N__37563\,
            in2 => \_gnd_net_\,
            in3 => \N__34050\,
            lcout => \HDA_STRAP.count_1_11\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_10\,
            carryout => \HDA_STRAP.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37455\,
            in2 => \_gnd_net_\,
            in3 => \N__34047\,
            lcout => \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_11\,
            carryout => \HDA_STRAP.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37257\,
            in2 => \_gnd_net_\,
            in3 => \N__34044\,
            lcout => \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_12\,
            carryout => \HDA_STRAP.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37322\,
            in2 => \_gnd_net_\,
            in3 => \N__34023\,
            lcout => \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_13\,
            carryout => \HDA_STRAP.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34176\,
            in2 => \_gnd_net_\,
            in3 => \N__34020\,
            lcout => \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_14\,
            carryout => \HDA_STRAP.un2_count_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__38691\,
            in1 => \N__34113\,
            in2 => \_gnd_net_\,
            in3 => \N__34017\,
            lcout => \HDA_STRAP.count_1_16\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un2_count_1_cry_15\,
            carryout => \HDA_STRAP.un2_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__34074\,
            in1 => \N__38686\,
            in2 => \_gnd_net_\,
            in3 => \N__34014\,
            lcout => \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNILF4V_17_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34011\,
            in1 => \N__33998\,
            in2 => \_gnd_net_\,
            in3 => \N__37780\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34166\,
            lcout => \HDA_STRAP.count_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38635\,
            ce => \N__37696\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34130\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38635\,
            ce => \N__37696\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDB8R_15_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34139\,
            in1 => \N__34129\,
            in2 => \_gnd_net_\,
            in3 => \N__37773\,
            lcout => \HDA_STRAP.un2_count_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIHFCT_6_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__34155\,
            in2 => \N__37785\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => \HDA_STRAP.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDB8R_0_15_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001010000"
        )
    port map (
            in0 => \N__34140\,
            in1 => \N__34131\,
            in2 => \N__34116\,
            in3 => \N__37775\,
            lcout => \HDA_STRAP.un25_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIEC8R_16_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37776\,
            in1 => \N__34104\,
            in2 => \_gnd_net_\,
            in3 => \N__34094\,
            lcout => \HDA_STRAP.un2_count_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34090\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38635\,
            ce => \N__37696\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIEC8R_0_16_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__37774\,
            in1 => \N__34103\,
            in2 => \N__34095\,
            in3 => \N__34073\,
            lcout => \HDA_STRAP.un25_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.un2_count_1_cry_0_c_RNO_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34350\,
            in1 => \N__34675\,
            in2 => \_gnd_net_\,
            in3 => \N__34056\,
            lcout => \DSW_PWRGD.un2_count_1_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNI70FA1_0_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__34938\,
            in1 => \N__34302\,
            in2 => \_gnd_net_\,
            in3 => \N__34793\,
            lcout => \DSW_PWRGD.count_rst_14\,
            ltout => \DSW_PWRGD.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNILCVT_0_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34349\,
            in2 => \N__34356\,
            in3 => \N__34674\,
            lcout => \DSW_PWRGD.count_i_0\,
            ltout => \DSW_PWRGD.count_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_0_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35025\,
            in2 => \N__34353\,
            in3 => \N__34305\,
            lcout => \DSW_PWRGD.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38485\,
            ce => \N__34723\,
            sr => \N__35024\
        );

    \DSW_PWRGD.un2_count_1_cry_10_c_RNIDHVO_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__34303\,
            in1 => \N__34220\,
            in2 => \N__35010\,
            in3 => \N__34331\,
            lcout => \DSW_PWRGD.count_rst_3\,
            ltout => \DSW_PWRGD.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIK54V1_11_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34676\,
            in1 => \_gnd_net_\,
            in2 => \N__34338\,
            in3 => \N__34202\,
            lcout => \DSW_PWRGD.un2_count_1_axb_11\,
            ltout => \DSW_PWRGD.un2_count_1_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_11_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__34304\,
            in1 => \N__34939\,
            in2 => \N__34224\,
            in3 => \N__34221\,
            lcout => \DSW_PWRGD.count_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38485\,
            ce => \N__34723\,
            sr => \N__35024\
        );

    \DSW_PWRGD.count_RNIK54V1_0_11_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__34677\,
            in1 => \N__34209\,
            in2 => \N__34524\,
            in3 => \N__34203\,
            lcout => \DSW_PWRGD.un12_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_12_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.count_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__34718\,
            sr => \N__35012\
        );

    \DSW_PWRGD.count_RNI2B5Q1_9_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34460\,
            in1 => \N__34685\,
            in2 => \_gnd_net_\,
            in3 => \N__34471\,
            lcout => \DSW_PWRGD.un2_count_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_9_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.count_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__34718\,
            sr => \N__35012\
        );

    \DSW_PWRGD.count_RNIM85V1_12_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34494\,
            in1 => \N__34686\,
            in2 => \_gnd_net_\,
            in3 => \N__34487\,
            lcout => \DSW_PWRGD.countZ0Z_12\,
            ltout => \DSW_PWRGD.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNI2B5Q1_0_9_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__34472\,
            in1 => \N__34461\,
            in2 => \N__34452\,
            in3 => \N__34688\,
            lcout => \DSW_PWRGD.un12_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIORVP1_4_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34415\,
            in1 => \N__34684\,
            in2 => \_gnd_net_\,
            in3 => \N__34429\,
            lcout => \DSW_PWRGD.un2_count_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_4_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.count_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38432\,
            ce => \N__34718\,
            sr => \N__35012\
        );

    \DSW_PWRGD.count_RNIORVP1_0_4_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100111"
        )
    port map (
            in0 => \N__34687\,
            in1 => \N__34430\,
            in2 => \N__34419\,
            in3 => \N__34407\,
            lcout => \DSW_PWRGD.un12_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_15_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34820\,
            lcout => \DSW_PWRGD.count_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38353\,
            ce => \N__34689\,
            sr => \N__35011\
        );

    \DSW_PWRGD.count_RNIOB6V1_13_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34362\,
            in1 => \N__34679\,
            in2 => \_gnd_net_\,
            in3 => \N__34370\,
            lcout => \DSW_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_13_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.count_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38353\,
            ce => \N__34689\,
            sr => \N__35011\
        );

    \DSW_PWRGD.count_RNIQE7V1_14_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35040\,
            in1 => \N__34690\,
            in2 => \_gnd_net_\,
            in3 => \N__35031\,
            lcout => \DSW_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_14_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35039\,
            lcout => \DSW_PWRGD.count_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38353\,
            ce => \N__34689\,
            sr => \N__35011\
        );

    \DSW_PWRGD.count_RNISH8V1_15_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__34821\,
            in1 => \N__34680\,
            in2 => \_gnd_net_\,
            in3 => \N__34812\,
            lcout => \DSW_PWRGD.countZ0Z_15\,
            ltout => \DSW_PWRGD.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNILCVT_0_0_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__34797\,
            in1 => \N__34781\,
            in2 => \N__34770\,
            in3 => \N__34767\,
            lcout => \DSW_PWRGD.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIIISP1_1_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34743\,
            in1 => \N__34678\,
            in2 => \_gnd_net_\,
            in3 => \N__34535\,
            lcout => \DSW_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIHPV41_7_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34506\,
            in1 => \N__35345\,
            in2 => \_gnd_net_\,
            in3 => \N__35890\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_7_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38419\,
            ce => \N__35891\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIJS051_8_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34500\,
            in1 => \N__35321\,
            in2 => \_gnd_net_\,
            in3 => \N__35887\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_8_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38419\,
            ce => \N__35891\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNILV151_9_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35291\,
            in1 => \N__35157\,
            in2 => \_gnd_net_\,
            in3 => \N__35889\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_9_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35292\,
            lcout => \VPP_VDDQ.count_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38419\,
            ce => \N__35891\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNINRAO_11_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35151\,
            in1 => \N__35192\,
            in2 => \_gnd_net_\,
            in3 => \N__35888\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_11_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35193\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38419\,
            ce => \N__35891\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_1_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35143\,
            in2 => \N__35130\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => \VPP_VDDQ.un4_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36084\,
            in2 => \_gnd_net_\,
            in3 => \N__35103\,
            lcout => \VPP_VDDQ.count_rst_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_1\,
            carryout => \VPP_VDDQ.un4_count_1_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35252\,
            in1 => \N__35100\,
            in2 => \_gnd_net_\,
            in3 => \N__35088\,
            lcout => \VPP_VDDQ.count_rst_8\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_2_cZ0\,
            carryout => \VPP_VDDQ.un4_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35254\,
            in1 => \N__35081\,
            in2 => \_gnd_net_\,
            in3 => \N__35070\,
            lcout => \VPP_VDDQ.count_rst_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_3\,
            carryout => \VPP_VDDQ.un4_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35250\,
            in1 => \N__35066\,
            in2 => \_gnd_net_\,
            in3 => \N__35043\,
            lcout => \VPP_VDDQ.count_rst_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_4\,
            carryout => \VPP_VDDQ.un4_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35706\,
            in3 => \N__35364\,
            lcout => \VPP_VDDQ.count_rst_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_5\,
            carryout => \VPP_VDDQ.un4_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__35251\,
            in1 => \_gnd_net_\,
            in2 => \N__35361\,
            in3 => \N__35337\,
            lcout => \VPP_VDDQ.count_rst_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_6\,
            carryout => \VPP_VDDQ.un4_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35253\,
            in1 => \N__35334\,
            in2 => \_gnd_net_\,
            in3 => \N__35313\,
            lcout => \VPP_VDDQ.count_rst_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_7\,
            carryout => \VPP_VDDQ.un4_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35258\,
            in1 => \N__35310\,
            in2 => \_gnd_net_\,
            in3 => \N__35280\,
            lcout => \VPP_VDDQ.count_rst_14\,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \VPP_VDDQ.un4_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35724\,
            in2 => \_gnd_net_\,
            in3 => \N__35262\,
            lcout => \VPP_VDDQ.count_rst\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_9\,
            carryout => \VPP_VDDQ.un4_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_10_c_RNI72NO_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__35259\,
            in1 => \N__35208\,
            in2 => \_gnd_net_\,
            in3 => \N__35181\,
            lcout => \VPP_VDDQ.count_rst_0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_10\,
            carryout => \VPP_VDDQ.un4_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35738\,
            in2 => \_gnd_net_\,
            in3 => \N__35178\,
            lcout => \VPP_VDDQ.count_rst_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_11\,
            carryout => \VPP_VDDQ.un4_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35171\,
            in2 => \_gnd_net_\,
            in3 => \N__35160\,
            lcout => \VPP_VDDQ.count_rst_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_12\,
            carryout => \VPP_VDDQ.un4_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35651\,
            in2 => \_gnd_net_\,
            in3 => \N__35631\,
            lcout => \VPP_VDDQ.count_rst_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un4_count_1_cry_13\,
            carryout => \VPP_VDDQ.un4_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__35627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35613\,
            lcout => \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_13_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35600\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38534\,
            ce => \N__35892\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_12_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35582\,
            lcout => \VPP_VDDQ.count_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38549\,
            ce => \N__35893\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35760\,
            lcout => \VPP_VDDQ.count_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38549\,
            ce => \N__35893\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_3_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35562\,
            lcout => \VPP_VDDQ.count_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38549\,
            ce => \N__35893\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__35538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38549\,
            ce => \N__35893\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIU6GQ_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__35514\,
            in1 => \N__35475\,
            in2 => \N__36212\,
            in3 => \N__35428\,
            lcout => \POWERLED.un1_clk_100khz_51_and_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100101111"
        )
    port map (
            in0 => \N__36123\,
            in1 => \N__36051\,
            in2 => \N__36213\,
            in3 => \N__36074\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__36073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36113\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38595\,
            ce => \N__36001\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__36112\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36072\,
            lcout => \VPP_VDDQ.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38595\,
            ce => \N__36001\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI7AQ41_0_2_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35771\,
            in1 => \N__35759\,
            in2 => \_gnd_net_\,
            in3 => \N__35818\,
            lcout => \VPP_VDDQ.un4_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI2PKG_1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36071\,
            in2 => \_gnd_net_\,
            in3 => \N__36050\,
            lcout => \VPP_VDDQ.count_en\,
            ltout => \VPP_VDDQ.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI7AQ41_2_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__35772\,
            in1 => \_gnd_net_\,
            in2 => \N__35763\,
            in3 => \N__35758\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.countZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI7AQ41_2_2_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__35739\,
            in1 => \N__35720\,
            in2 => \N__35709\,
            in3 => \N__35705\,
            lcout => \VPP_VDDQ.un13_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35676\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36262\,
            in2 => \N__36354\,
            in3 => \N__36345\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36342\,
            in2 => \N__36267\,
            in3 => \N__36336\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36284\,
            in2 => \N__36333\,
            in3 => \N__36324\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36321\,
            in2 => \N__36288\,
            in3 => \N__36315\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36563\,
            in1 => \N__36266\,
            in2 => \N__36312\,
            in3 => \N__36300\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36297\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36291\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36283\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36252\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36523\,
            in2 => \N__36225\,
            in3 => \N__36216\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36588\,
            in2 => \N__36528\,
            in3 => \N__36582\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36579\,
            in2 => \N__36570\,
            in3 => \N__36573\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36567\,
            in2 => \N__36543\,
            in3 => \N__36531\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36909\,
            in1 => \N__36527\,
            in2 => \N__36513\,
            in3 => \N__36504\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36501\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36495\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => \POWERLED.mult1_un145_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36492\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36477\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36889\,
            in2 => \N__36366\,
            in3 => \N__36357\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36966\,
            in2 => \N__36894\,
            in3 => \N__36960\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36911\,
            in2 => \N__36957\,
            in3 => \N__36948\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36945\,
            in2 => \N__36915\,
            in3 => \N__36939\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__37052\,
            in1 => \N__36893\,
            in2 => \N__36936\,
            in3 => \N__36927\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__36924\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36918\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36910\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36877\,
            in2 => \_gnd_net_\,
            in3 => \N__36716\,
            lcout => \POWERLED.g0_9_0\,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37027\,
            in2 => \N__36618\,
            in3 => \N__36591\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37203\,
            in2 => \N__37032\,
            in3 => \N__37179\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37055\,
            in2 => \N__37176\,
            in3 => \N__37152\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37149\,
            in2 => \N__37059\,
            in3 => \N__37128\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__37075\,
            in1 => \N__37031\,
            in2 => \N__37125\,
            in3 => \N__37104\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__37101\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37095\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37054\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB69T_3_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36986\,
            in1 => \N__37766\,
            in2 => \_gnd_net_\,
            in3 => \N__36976\,
            lcout => \HDA_STRAP.un2_count_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__37692\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB69T_0_3_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000101"
        )
    port map (
            in0 => \N__37011\,
            in1 => \N__37769\,
            in2 => \N__36990\,
            in3 => \N__36977\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un25_clk_100khz_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIUE4N3_3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37293\,
            in1 => \N__37425\,
            in2 => \N__37326\,
            in3 => \N__37230\,
            lcout => \HDA_STRAP.un25_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNID30V_0_13_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000011"
        )
    port map (
            in0 => \N__37271\,
            in1 => \N__37323\,
            in2 => \N__37287\,
            in3 => \N__37768\,
            lcout => \HDA_STRAP.un25_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37272\,
            lcout => \HDA_STRAP.count_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38634\,
            ce => \N__37692\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNID30V_13_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37283\,
            in1 => \N__37270\,
            in2 => \_gnd_net_\,
            in3 => \N__37765\,
            lcout => \HDA_STRAP.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIFCBT_0_5_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100011"
        )
    port map (
            in0 => \N__37767\,
            in1 => \N__37251\,
            in2 => \N__37395\,
            in3 => \N__37410\,
            lcout => \HDA_STRAP.un25_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37212\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38624\,
            ce => \N__37694\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38624\,
            ce => \N__37694\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNINOFT_9_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37448\,
            in1 => \N__37438\,
            in2 => \_gnd_net_\,
            in3 => \N__37760\,
            lcout => \HDA_STRAP.un2_count_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB0VU_12_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37761\,
            in1 => \N__37218\,
            in2 => \_gnd_net_\,
            in3 => \N__37211\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => \HDA_STRAP.countZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNINOFT_0_9_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__37449\,
            in1 => \N__37439\,
            in2 => \N__37428\,
            in3 => \N__37763\,
            lcout => \HDA_STRAP.un25_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIFCBT_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37762\,
            in1 => \N__37391\,
            in2 => \_gnd_net_\,
            in3 => \N__37408\,
            lcout => \HDA_STRAP.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37409\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38624\,
            ce => \N__37694\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI0THV_10_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__37764\,
            in1 => \N__37380\,
            in2 => \N__37368\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI938T_2_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37782\,
            in1 => \N__37587\,
            in2 => \_gnd_net_\,
            in3 => \N__37598\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIOR6P_1_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__37625\,
            in1 => \N__37781\,
            in2 => \_gnd_net_\,
            in3 => \N__37332\,
            lcout => \HDA_STRAP.un2_count_1_axb_1\,
            ltout => \HDA_STRAP.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__37476\,
            in1 => \_gnd_net_\,
            in2 => \N__37350\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38637\,
            ce => \N__37693\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI_1_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__37346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37475\,
            lcout => \HDA_STRAP.count_RNIZ0Z_1\,
            ltout => \HDA_STRAP.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIOR6P_0_1_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__37784\,
            in1 => \N__37626\,
            in2 => \N__37617\,
            in3 => \N__37613\,
            lcout => \HDA_STRAP.un25_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37599\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.count_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38637\,
            ce => \N__37693\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI9TTU_11_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__37783\,
            in1 => \N__37569\,
            in2 => \_gnd_net_\,
            in3 => \N__37581\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37580\,
            lcout => \HDA_STRAP.count_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38637\,
            ce => \N__37693\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI68FK1_1_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__37562\,
            in1 => \N__37551\,
            in2 => \N__37487\,
            in3 => \N__37545\,
            lcout => \HDA_STRAP.un25_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNILLET_0_8_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__37813\,
            in1 => \N__37539\,
            in2 => \N__37800\,
            in3 => \N__37759\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un25_clk_100khz_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI6OA47_8_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37521\,
            in1 => \N__37512\,
            in2 => \N__37503\,
            in3 => \N__37500\,
            lcout => \HDA_STRAP.count_RNI6OA47Z0Z_8\,
            ltout => \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI_0_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37494\,
            in3 => \N__37483\,
            lcout => OPEN,
            ltout => \HDA_STRAP.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNINQ6P_0_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__37758\,
            in1 => \_gnd_net_\,
            in2 => \N__37491\,
            in3 => \N__38643\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => \HDA_STRAP.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38715\,
            in3 => \N__38685\,
            lcout => \HDA_STRAP.count_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38636\,
            ce => \N__37697\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37814\,
            lcout => \HDA_STRAP.count_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__38636\,
            ce => \N__37697\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNILLET_8_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37815\,
            in1 => \N__37796\,
            in2 => \_gnd_net_\,
            in3 => \N__37757\,
            lcout => \HDA_STRAP.un2_count_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
