// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 7 2022 10:06:34

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    output SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__35432;
    wire N__35431;
    wire N__35430;
    wire N__35423;
    wire N__35422;
    wire N__35421;
    wire N__35414;
    wire N__35413;
    wire N__35412;
    wire N__35405;
    wire N__35404;
    wire N__35403;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35387;
    wire N__35386;
    wire N__35385;
    wire N__35378;
    wire N__35377;
    wire N__35376;
    wire N__35369;
    wire N__35368;
    wire N__35367;
    wire N__35360;
    wire N__35359;
    wire N__35358;
    wire N__35351;
    wire N__35350;
    wire N__35349;
    wire N__35342;
    wire N__35341;
    wire N__35340;
    wire N__35333;
    wire N__35332;
    wire N__35331;
    wire N__35324;
    wire N__35323;
    wire N__35322;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35288;
    wire N__35287;
    wire N__35286;
    wire N__35279;
    wire N__35278;
    wire N__35277;
    wire N__35270;
    wire N__35269;
    wire N__35268;
    wire N__35261;
    wire N__35260;
    wire N__35259;
    wire N__35252;
    wire N__35251;
    wire N__35250;
    wire N__35243;
    wire N__35242;
    wire N__35241;
    wire N__35234;
    wire N__35233;
    wire N__35232;
    wire N__35225;
    wire N__35224;
    wire N__35223;
    wire N__35216;
    wire N__35215;
    wire N__35214;
    wire N__35207;
    wire N__35206;
    wire N__35205;
    wire N__35198;
    wire N__35197;
    wire N__35196;
    wire N__35189;
    wire N__35188;
    wire N__35187;
    wire N__35180;
    wire N__35179;
    wire N__35178;
    wire N__35171;
    wire N__35170;
    wire N__35169;
    wire N__35162;
    wire N__35161;
    wire N__35160;
    wire N__35153;
    wire N__35152;
    wire N__35151;
    wire N__35144;
    wire N__35143;
    wire N__35142;
    wire N__35135;
    wire N__35134;
    wire N__35133;
    wire N__35126;
    wire N__35125;
    wire N__35124;
    wire N__35117;
    wire N__35116;
    wire N__35115;
    wire N__35108;
    wire N__35107;
    wire N__35106;
    wire N__35099;
    wire N__35098;
    wire N__35097;
    wire N__35090;
    wire N__35089;
    wire N__35088;
    wire N__35081;
    wire N__35080;
    wire N__35079;
    wire N__35072;
    wire N__35071;
    wire N__35070;
    wire N__35063;
    wire N__35062;
    wire N__35061;
    wire N__35054;
    wire N__35053;
    wire N__35052;
    wire N__35045;
    wire N__35044;
    wire N__35043;
    wire N__35036;
    wire N__35035;
    wire N__35034;
    wire N__35027;
    wire N__35026;
    wire N__35025;
    wire N__35018;
    wire N__35017;
    wire N__35016;
    wire N__35009;
    wire N__35008;
    wire N__35007;
    wire N__35000;
    wire N__34999;
    wire N__34998;
    wire N__34991;
    wire N__34990;
    wire N__34989;
    wire N__34982;
    wire N__34981;
    wire N__34980;
    wire N__34973;
    wire N__34972;
    wire N__34971;
    wire N__34964;
    wire N__34963;
    wire N__34962;
    wire N__34955;
    wire N__34954;
    wire N__34953;
    wire N__34946;
    wire N__34945;
    wire N__34944;
    wire N__34937;
    wire N__34936;
    wire N__34935;
    wire N__34928;
    wire N__34927;
    wire N__34926;
    wire N__34919;
    wire N__34918;
    wire N__34917;
    wire N__34910;
    wire N__34909;
    wire N__34908;
    wire N__34891;
    wire N__34890;
    wire N__34889;
    wire N__34888;
    wire N__34887;
    wire N__34886;
    wire N__34885;
    wire N__34884;
    wire N__34883;
    wire N__34882;
    wire N__34881;
    wire N__34880;
    wire N__34879;
    wire N__34878;
    wire N__34877;
    wire N__34876;
    wire N__34875;
    wire N__34874;
    wire N__34873;
    wire N__34872;
    wire N__34871;
    wire N__34870;
    wire N__34869;
    wire N__34868;
    wire N__34867;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34863;
    wire N__34862;
    wire N__34861;
    wire N__34860;
    wire N__34859;
    wire N__34858;
    wire N__34857;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34850;
    wire N__34849;
    wire N__34848;
    wire N__34847;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34842;
    wire N__34841;
    wire N__34840;
    wire N__34839;
    wire N__34830;
    wire N__34821;
    wire N__34812;
    wire N__34805;
    wire N__34798;
    wire N__34789;
    wire N__34780;
    wire N__34771;
    wire N__34762;
    wire N__34759;
    wire N__34754;
    wire N__34745;
    wire N__34736;
    wire N__34729;
    wire N__34726;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34714;
    wire N__34713;
    wire N__34712;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34706;
    wire N__34703;
    wire N__34700;
    wire N__34697;
    wire N__34696;
    wire N__34693;
    wire N__34690;
    wire N__34689;
    wire N__34688;
    wire N__34687;
    wire N__34684;
    wire N__34681;
    wire N__34678;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34654;
    wire N__34651;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34562;
    wire N__34561;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34538;
    wire N__34537;
    wire N__34534;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34506;
    wire N__34501;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34489;
    wire N__34486;
    wire N__34477;
    wire N__34474;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34462;
    wire N__34461;
    wire N__34460;
    wire N__34459;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34451;
    wire N__34450;
    wire N__34449;
    wire N__34446;
    wire N__34445;
    wire N__34444;
    wire N__34441;
    wire N__34440;
    wire N__34439;
    wire N__34438;
    wire N__34435;
    wire N__34434;
    wire N__34433;
    wire N__34432;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34426;
    wire N__34425;
    wire N__34422;
    wire N__34421;
    wire N__34418;
    wire N__34417;
    wire N__34416;
    wire N__34413;
    wire N__34412;
    wire N__34409;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34394;
    wire N__34391;
    wire N__34390;
    wire N__34389;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34378;
    wire N__34375;
    wire N__34374;
    wire N__34373;
    wire N__34372;
    wire N__34369;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34361;
    wire N__34358;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34350;
    wire N__34349;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34332;
    wire N__34329;
    wire N__34328;
    wire N__34325;
    wire N__34324;
    wire N__34323;
    wire N__34322;
    wire N__34321;
    wire N__34318;
    wire N__34311;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34294;
    wire N__34293;
    wire N__34292;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34275;
    wire N__34272;
    wire N__34271;
    wire N__34268;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34241;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34233;
    wire N__34230;
    wire N__34225;
    wire N__34224;
    wire N__34223;
    wire N__34222;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34185;
    wire N__34182;
    wire N__34171;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34163;
    wire N__34162;
    wire N__34161;
    wire N__34158;
    wire N__34153;
    wire N__34148;
    wire N__34145;
    wire N__34144;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34126;
    wire N__34119;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34086;
    wire N__34085;
    wire N__34084;
    wire N__34081;
    wire N__34080;
    wire N__34073;
    wire N__34070;
    wire N__34069;
    wire N__34064;
    wire N__34059;
    wire N__34056;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34013;
    wire N__34010;
    wire N__34003;
    wire N__34000;
    wire N__33999;
    wire N__33998;
    wire N__33997;
    wire N__33996;
    wire N__33993;
    wire N__33984;
    wire N__33983;
    wire N__33980;
    wire N__33975;
    wire N__33970;
    wire N__33963;
    wire N__33960;
    wire N__33955;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33937;
    wire N__33932;
    wire N__33929;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33906;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33876;
    wire N__33875;
    wire N__33872;
    wire N__33869;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33853;
    wire N__33850;
    wire N__33843;
    wire N__33830;
    wire N__33825;
    wire N__33820;
    wire N__33815;
    wire N__33804;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33758;
    wire N__33751;
    wire N__33746;
    wire N__33739;
    wire N__33730;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33705;
    wire N__33704;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33683;
    wire N__33680;
    wire N__33673;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33661;
    wire N__33658;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33646;
    wire N__33643;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33631;
    wire N__33628;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33616;
    wire N__33613;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33598;
    wire N__33595;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33583;
    wire N__33580;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33568;
    wire N__33565;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33543;
    wire N__33540;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33489;
    wire N__33488;
    wire N__33487;
    wire N__33486;
    wire N__33485;
    wire N__33484;
    wire N__33483;
    wire N__33480;
    wire N__33477;
    wire N__33476;
    wire N__33475;
    wire N__33472;
    wire N__33471;
    wire N__33470;
    wire N__33469;
    wire N__33466;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33455;
    wire N__33454;
    wire N__33453;
    wire N__33444;
    wire N__33437;
    wire N__33434;
    wire N__33429;
    wire N__33424;
    wire N__33419;
    wire N__33418;
    wire N__33417;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33411;
    wire N__33408;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33392;
    wire N__33383;
    wire N__33370;
    wire N__33355;
    wire N__33354;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33333;
    wire N__33332;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33324;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33318;
    wire N__33317;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33271;
    wire N__33268;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33257;
    wire N__33254;
    wire N__33247;
    wire N__33238;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33211;
    wire N__33206;
    wire N__33201;
    wire N__33194;
    wire N__33175;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33160;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33145;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33133;
    wire N__33130;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33118;
    wire N__33115;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33100;
    wire N__33097;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33085;
    wire N__33082;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33070;
    wire N__33067;
    wire N__33066;
    wire N__33061;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33043;
    wire N__33040;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33025;
    wire N__33024;
    wire N__33021;
    wire N__33020;
    wire N__33019;
    wire N__33018;
    wire N__33015;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32970;
    wire N__32969;
    wire N__32968;
    wire N__32967;
    wire N__32966;
    wire N__32965;
    wire N__32964;
    wire N__32963;
    wire N__32960;
    wire N__32957;
    wire N__32956;
    wire N__32953;
    wire N__32952;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32939;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32901;
    wire N__32898;
    wire N__32893;
    wire N__32886;
    wire N__32883;
    wire N__32882;
    wire N__32877;
    wire N__32874;
    wire N__32867;
    wire N__32862;
    wire N__32859;
    wire N__32854;
    wire N__32849;
    wire N__32842;
    wire N__32841;
    wire N__32840;
    wire N__32837;
    wire N__32832;
    wire N__32829;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32818;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32752;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32736;
    wire N__32735;
    wire N__32732;
    wire N__32729;
    wire N__32728;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32700;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32669;
    wire N__32666;
    wire N__32659;
    wire N__32658;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32617;
    wire N__32614;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32607;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32587;
    wire N__32584;
    wire N__32581;
    wire N__32580;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32556;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32544;
    wire N__32541;
    wire N__32540;
    wire N__32537;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32521;
    wire N__32518;
    wire N__32515;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32485;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32473;
    wire N__32470;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32455;
    wire N__32454;
    wire N__32449;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32434;
    wire N__32433;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32419;
    wire N__32418;
    wire N__32415;
    wire N__32414;
    wire N__32413;
    wire N__32410;
    wire N__32407;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32389;
    wire N__32388;
    wire N__32383;
    wire N__32380;
    wire N__32377;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32364;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32350;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32338;
    wire N__32335;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32316;
    wire N__32311;
    wire N__32308;
    wire N__32305;
    wire N__32304;
    wire N__32301;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32283;
    wire N__32280;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32256;
    wire N__32251;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32228;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32216;
    wire N__32213;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32190;
    wire N__32185;
    wire N__32182;
    wire N__32181;
    wire N__32178;
    wire N__32177;
    wire N__32174;
    wire N__32173;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32169;
    wire N__32168;
    wire N__32167;
    wire N__32166;
    wire N__32165;
    wire N__32164;
    wire N__32155;
    wire N__32154;
    wire N__32153;
    wire N__32152;
    wire N__32151;
    wire N__32150;
    wire N__32149;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32143;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32107;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32091;
    wire N__32090;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32083;
    wire N__32074;
    wire N__32073;
    wire N__32070;
    wire N__32069;
    wire N__32068;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32044;
    wire N__32033;
    wire N__32030;
    wire N__32021;
    wire N__32002;
    wire N__32001;
    wire N__31998;
    wire N__31993;
    wire N__31990;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31984;
    wire N__31983;
    wire N__31982;
    wire N__31981;
    wire N__31980;
    wire N__31979;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31973;
    wire N__31972;
    wire N__31971;
    wire N__31968;
    wire N__31957;
    wire N__31954;
    wire N__31953;
    wire N__31952;
    wire N__31951;
    wire N__31950;
    wire N__31949;
    wire N__31948;
    wire N__31947;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31936;
    wire N__31931;
    wire N__31928;
    wire N__31927;
    wire N__31926;
    wire N__31925;
    wire N__31922;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31910;
    wire N__31909;
    wire N__31908;
    wire N__31907;
    wire N__31906;
    wire N__31903;
    wire N__31902;
    wire N__31901;
    wire N__31898;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31876;
    wire N__31871;
    wire N__31866;
    wire N__31861;
    wire N__31856;
    wire N__31845;
    wire N__31836;
    wire N__31829;
    wire N__31824;
    wire N__31815;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31795;
    wire N__31794;
    wire N__31793;
    wire N__31792;
    wire N__31791;
    wire N__31790;
    wire N__31787;
    wire N__31786;
    wire N__31785;
    wire N__31784;
    wire N__31783;
    wire N__31782;
    wire N__31781;
    wire N__31780;
    wire N__31779;
    wire N__31778;
    wire N__31777;
    wire N__31776;
    wire N__31775;
    wire N__31774;
    wire N__31771;
    wire N__31770;
    wire N__31767;
    wire N__31766;
    wire N__31765;
    wire N__31764;
    wire N__31763;
    wire N__31762;
    wire N__31749;
    wire N__31748;
    wire N__31747;
    wire N__31746;
    wire N__31745;
    wire N__31744;
    wire N__31743;
    wire N__31742;
    wire N__31739;
    wire N__31730;
    wire N__31721;
    wire N__31710;
    wire N__31707;
    wire N__31702;
    wire N__31699;
    wire N__31690;
    wire N__31687;
    wire N__31680;
    wire N__31671;
    wire N__31664;
    wire N__31661;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31632;
    wire N__31631;
    wire N__31628;
    wire N__31627;
    wire N__31626;
    wire N__31623;
    wire N__31622;
    wire N__31621;
    wire N__31620;
    wire N__31619;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31607;
    wire N__31606;
    wire N__31605;
    wire N__31604;
    wire N__31601;
    wire N__31598;
    wire N__31595;
    wire N__31594;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31584;
    wire N__31577;
    wire N__31570;
    wire N__31569;
    wire N__31568;
    wire N__31567;
    wire N__31566;
    wire N__31559;
    wire N__31556;
    wire N__31553;
    wire N__31552;
    wire N__31551;
    wire N__31550;
    wire N__31549;
    wire N__31548;
    wire N__31547;
    wire N__31542;
    wire N__31535;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31517;
    wire N__31510;
    wire N__31507;
    wire N__31502;
    wire N__31495;
    wire N__31480;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31429;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31353;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31263;
    wire N__31258;
    wire N__31255;
    wire N__31254;
    wire N__31253;
    wire N__31250;
    wire N__31245;
    wire N__31240;
    wire N__31237;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31180;
    wire N__31177;
    wire N__31176;
    wire N__31173;
    wire N__31168;
    wire N__31167;
    wire N__31166;
    wire N__31165;
    wire N__31164;
    wire N__31163;
    wire N__31160;
    wire N__31159;
    wire N__31158;
    wire N__31155;
    wire N__31154;
    wire N__31153;
    wire N__31150;
    wire N__31149;
    wire N__31148;
    wire N__31147;
    wire N__31146;
    wire N__31145;
    wire N__31142;
    wire N__31141;
    wire N__31140;
    wire N__31139;
    wire N__31134;
    wire N__31133;
    wire N__31132;
    wire N__31129;
    wire N__31124;
    wire N__31121;
    wire N__31120;
    wire N__31117;
    wire N__31116;
    wire N__31115;
    wire N__31114;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31090;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31068;
    wire N__31065;
    wire N__31060;
    wire N__31055;
    wire N__31050;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31032;
    wire N__31029;
    wire N__31028;
    wire N__31027;
    wire N__31026;
    wire N__31019;
    wire N__31016;
    wire N__31013;
    wire N__31006;
    wire N__31001;
    wire N__30998;
    wire N__30991;
    wire N__30984;
    wire N__30981;
    wire N__30972;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30952;
    wire N__30951;
    wire N__30950;
    wire N__30947;
    wire N__30942;
    wire N__30941;
    wire N__30940;
    wire N__30939;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30923;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30880;
    wire N__30879;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30825;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30810;
    wire N__30809;
    wire N__30808;
    wire N__30807;
    wire N__30804;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30789;
    wire N__30786;
    wire N__30785;
    wire N__30784;
    wire N__30783;
    wire N__30782;
    wire N__30781;
    wire N__30780;
    wire N__30779;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30726;
    wire N__30721;
    wire N__30718;
    wire N__30717;
    wire N__30716;
    wire N__30713;
    wire N__30708;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30660;
    wire N__30657;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30636;
    wire N__30633;
    wire N__30632;
    wire N__30631;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30620;
    wire N__30617;
    wire N__30616;
    wire N__30615;
    wire N__30614;
    wire N__30613;
    wire N__30612;
    wire N__30607;
    wire N__30606;
    wire N__30605;
    wire N__30604;
    wire N__30603;
    wire N__30602;
    wire N__30601;
    wire N__30600;
    wire N__30599;
    wire N__30596;
    wire N__30589;
    wire N__30580;
    wire N__30579;
    wire N__30578;
    wire N__30577;
    wire N__30576;
    wire N__30575;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30558;
    wire N__30549;
    wire N__30548;
    wire N__30547;
    wire N__30546;
    wire N__30539;
    wire N__30532;
    wire N__30531;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30511;
    wire N__30508;
    wire N__30503;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30491;
    wire N__30490;
    wire N__30485;
    wire N__30482;
    wire N__30477;
    wire N__30474;
    wire N__30469;
    wire N__30466;
    wire N__30465;
    wire N__30462;
    wire N__30457;
    wire N__30454;
    wire N__30447;
    wire N__30444;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30411;
    wire N__30410;
    wire N__30407;
    wire N__30406;
    wire N__30403;
    wire N__30402;
    wire N__30401;
    wire N__30400;
    wire N__30399;
    wire N__30396;
    wire N__30389;
    wire N__30380;
    wire N__30375;
    wire N__30372;
    wire N__30371;
    wire N__30370;
    wire N__30365;
    wire N__30360;
    wire N__30359;
    wire N__30358;
    wire N__30353;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30327;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30292;
    wire N__30289;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30274;
    wire N__30273;
    wire N__30266;
    wire N__30261;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30238;
    wire N__30237;
    wire N__30234;
    wire N__30233;
    wire N__30230;
    wire N__30229;
    wire N__30228;
    wire N__30225;
    wire N__30222;
    wire N__30219;
    wire N__30218;
    wire N__30215;
    wire N__30214;
    wire N__30213;
    wire N__30212;
    wire N__30209;
    wire N__30206;
    wire N__30201;
    wire N__30194;
    wire N__30191;
    wire N__30190;
    wire N__30189;
    wire N__30188;
    wire N__30185;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30165;
    wire N__30164;
    wire N__30161;
    wire N__30160;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30149;
    wire N__30144;
    wire N__30141;
    wire N__30136;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30108;
    wire N__30097;
    wire N__30096;
    wire N__30095;
    wire N__30094;
    wire N__30089;
    wire N__30084;
    wire N__30079;
    wire N__30076;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30051;
    wire N__30050;
    wire N__30049;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30038;
    wire N__30037;
    wire N__30032;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30013;
    wire N__30004;
    wire N__30003;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29995;
    wire N__29994;
    wire N__29993;
    wire N__29992;
    wire N__29991;
    wire N__29990;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29986;
    wire N__29985;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29981;
    wire N__29978;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29958;
    wire N__29953;
    wire N__29948;
    wire N__29945;
    wire N__29944;
    wire N__29943;
    wire N__29940;
    wire N__29939;
    wire N__29936;
    wire N__29931;
    wire N__29928;
    wire N__29923;
    wire N__29918;
    wire N__29917;
    wire N__29916;
    wire N__29915;
    wire N__29914;
    wire N__29913;
    wire N__29908;
    wire N__29905;
    wire N__29900;
    wire N__29897;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29880;
    wire N__29875;
    wire N__29872;
    wire N__29867;
    wire N__29864;
    wire N__29857;
    wire N__29854;
    wire N__29833;
    wire N__29830;
    wire N__29829;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29825;
    wire N__29822;
    wire N__29821;
    wire N__29820;
    wire N__29817;
    wire N__29816;
    wire N__29813;
    wire N__29812;
    wire N__29811;
    wire N__29810;
    wire N__29809;
    wire N__29808;
    wire N__29807;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29790;
    wire N__29781;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29773;
    wire N__29772;
    wire N__29763;
    wire N__29760;
    wire N__29759;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29745;
    wire N__29744;
    wire N__29743;
    wire N__29738;
    wire N__29735;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29717;
    wire N__29714;
    wire N__29713;
    wire N__29712;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29697;
    wire N__29694;
    wire N__29689;
    wire N__29682;
    wire N__29679;
    wire N__29678;
    wire N__29675;
    wire N__29672;
    wire N__29669;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29626;
    wire N__29625;
    wire N__29622;
    wire N__29621;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29593;
    wire N__29592;
    wire N__29591;
    wire N__29590;
    wire N__29589;
    wire N__29588;
    wire N__29587;
    wire N__29584;
    wire N__29583;
    wire N__29582;
    wire N__29575;
    wire N__29574;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29564;
    wire N__29557;
    wire N__29554;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29525;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29505;
    wire N__29504;
    wire N__29501;
    wire N__29496;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29481;
    wire N__29480;
    wire N__29479;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29473;
    wire N__29470;
    wire N__29469;
    wire N__29466;
    wire N__29461;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29455;
    wire N__29452;
    wire N__29451;
    wire N__29448;
    wire N__29447;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29426;
    wire N__29425;
    wire N__29424;
    wire N__29419;
    wire N__29412;
    wire N__29409;
    wire N__29398;
    wire N__29393;
    wire N__29392;
    wire N__29389;
    wire N__29384;
    wire N__29383;
    wire N__29382;
    wire N__29375;
    wire N__29372;
    wire N__29371;
    wire N__29366;
    wire N__29361;
    wire N__29358;
    wire N__29353;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29334;
    wire N__29333;
    wire N__29332;
    wire N__29331;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29322;
    wire N__29319;
    wire N__29318;
    wire N__29317;
    wire N__29316;
    wire N__29315;
    wire N__29314;
    wire N__29313;
    wire N__29308;
    wire N__29307;
    wire N__29306;
    wire N__29305;
    wire N__29304;
    wire N__29303;
    wire N__29302;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29246;
    wire N__29241;
    wire N__29236;
    wire N__29229;
    wire N__29224;
    wire N__29223;
    wire N__29220;
    wire N__29215;
    wire N__29210;
    wire N__29203;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29188;
    wire N__29185;
    wire N__29176;
    wire N__29173;
    wire N__29166;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29127;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29115;
    wire N__29110;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29067;
    wire N__29066;
    wire N__29063;
    wire N__29062;
    wire N__29061;
    wire N__29060;
    wire N__29055;
    wire N__29052;
    wire N__29051;
    wire N__29050;
    wire N__29049;
    wire N__29044;
    wire N__29041;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29026;
    wire N__29021;
    wire N__29018;
    wire N__29011;
    wire N__29008;
    wire N__29003;
    wire N__29000;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28984;
    wire N__28983;
    wire N__28982;
    wire N__28981;
    wire N__28980;
    wire N__28979;
    wire N__28974;
    wire N__28971;
    wire N__28966;
    wire N__28963;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28955;
    wire N__28950;
    wire N__28945;
    wire N__28942;
    wire N__28941;
    wire N__28932;
    wire N__28927;
    wire N__28924;
    wire N__28917;
    wire N__28914;
    wire N__28913;
    wire N__28912;
    wire N__28911;
    wire N__28910;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28901;
    wire N__28898;
    wire N__28893;
    wire N__28886;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28871;
    wire N__28868;
    wire N__28861;
    wire N__28858;
    wire N__28847;
    wire N__28842;
    wire N__28839;
    wire N__28836;
    wire N__28831;
    wire N__28828;
    wire N__28827;
    wire N__28824;
    wire N__28821;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28755;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28693;
    wire N__28690;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28656;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28644;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28600;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28578;
    wire N__28575;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28509;
    wire N__28506;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28473;
    wire N__28470;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28444;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28362;
    wire N__28357;
    wire N__28354;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28332;
    wire N__28327;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28299;
    wire N__28294;
    wire N__28291;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28279;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28271;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28253;
    wire N__28246;
    wire N__28243;
    wire N__28242;
    wire N__28241;
    wire N__28240;
    wire N__28239;
    wire N__28236;
    wire N__28235;
    wire N__28234;
    wire N__28229;
    wire N__28228;
    wire N__28227;
    wire N__28226;
    wire N__28225;
    wire N__28224;
    wire N__28223;
    wire N__28222;
    wire N__28219;
    wire N__28218;
    wire N__28217;
    wire N__28216;
    wire N__28213;
    wire N__28212;
    wire N__28211;
    wire N__28210;
    wire N__28209;
    wire N__28208;
    wire N__28207;
    wire N__28206;
    wire N__28205;
    wire N__28204;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28182;
    wire N__28179;
    wire N__28174;
    wire N__28171;
    wire N__28170;
    wire N__28169;
    wire N__28168;
    wire N__28167;
    wire N__28166;
    wire N__28163;
    wire N__28160;
    wire N__28151;
    wire N__28140;
    wire N__28131;
    wire N__28128;
    wire N__28121;
    wire N__28114;
    wire N__28107;
    wire N__28098;
    wire N__28095;
    wire N__28084;
    wire N__28083;
    wire N__28080;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28064;
    wire N__28061;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28023;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28002;
    wire N__28001;
    wire N__27998;
    wire N__27993;
    wire N__27990;
    wire N__27985;
    wire N__27984;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27966;
    wire N__27965;
    wire N__27962;
    wire N__27957;
    wire N__27952;
    wire N__27949;
    wire N__27948;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27910;
    wire N__27909;
    wire N__27906;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27898;
    wire N__27895;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27853;
    wire N__27852;
    wire N__27851;
    wire N__27850;
    wire N__27849;
    wire N__27846;
    wire N__27845;
    wire N__27844;
    wire N__27839;
    wire N__27838;
    wire N__27835;
    wire N__27834;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27822;
    wire N__27821;
    wire N__27820;
    wire N__27815;
    wire N__27812;
    wire N__27811;
    wire N__27810;
    wire N__27809;
    wire N__27808;
    wire N__27807;
    wire N__27806;
    wire N__27805;
    wire N__27804;
    wire N__27803;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27784;
    wire N__27781;
    wire N__27780;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27755;
    wire N__27750;
    wire N__27743;
    wire N__27732;
    wire N__27727;
    wire N__27722;
    wire N__27703;
    wire N__27702;
    wire N__27701;
    wire N__27700;
    wire N__27699;
    wire N__27698;
    wire N__27697;
    wire N__27696;
    wire N__27695;
    wire N__27694;
    wire N__27693;
    wire N__27692;
    wire N__27691;
    wire N__27686;
    wire N__27685;
    wire N__27674;
    wire N__27671;
    wire N__27670;
    wire N__27659;
    wire N__27656;
    wire N__27653;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27633;
    wire N__27628;
    wire N__27625;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27610;
    wire N__27607;
    wire N__27606;
    wire N__27605;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27576;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27552;
    wire N__27551;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27526;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27508;
    wire N__27505;
    wire N__27502;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27477;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27465;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27429;
    wire N__27428;
    wire N__27425;
    wire N__27424;
    wire N__27423;
    wire N__27422;
    wire N__27421;
    wire N__27420;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27412;
    wire N__27411;
    wire N__27408;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27392;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27349;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27340;
    wire N__27339;
    wire N__27336;
    wire N__27335;
    wire N__27334;
    wire N__27333;
    wire N__27326;
    wire N__27323;
    wire N__27320;
    wire N__27319;
    wire N__27316;
    wire N__27315;
    wire N__27312;
    wire N__27307;
    wire N__27304;
    wire N__27303;
    wire N__27302;
    wire N__27299;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27281;
    wire N__27278;
    wire N__27277;
    wire N__27274;
    wire N__27269;
    wire N__27266;
    wire N__27265;
    wire N__27264;
    wire N__27259;
    wire N__27254;
    wire N__27251;
    wire N__27248;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27223;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27162;
    wire N__27161;
    wire N__27160;
    wire N__27155;
    wire N__27154;
    wire N__27153;
    wire N__27152;
    wire N__27151;
    wire N__27146;
    wire N__27145;
    wire N__27144;
    wire N__27143;
    wire N__27142;
    wire N__27141;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27110;
    wire N__27105;
    wire N__27102;
    wire N__27097;
    wire N__27094;
    wire N__27089;
    wire N__27086;
    wire N__27079;
    wire N__27078;
    wire N__27073;
    wire N__27070;
    wire N__27069;
    wire N__27066;
    wire N__27055;
    wire N__27054;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27032;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27014;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26982;
    wire N__26981;
    wire N__26974;
    wire N__26971;
    wire N__26970;
    wire N__26969;
    wire N__26966;
    wire N__26963;
    wire N__26960;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26946;
    wire N__26943;
    wire N__26942;
    wire N__26939;
    wire N__26934;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26920;
    wire N__26919;
    wire N__26918;
    wire N__26917;
    wire N__26916;
    wire N__26915;
    wire N__26914;
    wire N__26913;
    wire N__26912;
    wire N__26911;
    wire N__26910;
    wire N__26909;
    wire N__26908;
    wire N__26907;
    wire N__26906;
    wire N__26905;
    wire N__26896;
    wire N__26887;
    wire N__26880;
    wire N__26875;
    wire N__26868;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26862;
    wire N__26861;
    wire N__26856;
    wire N__26853;
    wire N__26848;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26828;
    wire N__26825;
    wire N__26820;
    wire N__26815;
    wire N__26814;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26769;
    wire N__26768;
    wire N__26767;
    wire N__26766;
    wire N__26765;
    wire N__26760;
    wire N__26759;
    wire N__26756;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26742;
    wire N__26741;
    wire N__26738;
    wire N__26733;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26717;
    wire N__26716;
    wire N__26715;
    wire N__26712;
    wire N__26701;
    wire N__26700;
    wire N__26695;
    wire N__26694;
    wire N__26693;
    wire N__26692;
    wire N__26691;
    wire N__26690;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26682;
    wire N__26679;
    wire N__26678;
    wire N__26677;
    wire N__26674;
    wire N__26667;
    wire N__26660;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26644;
    wire N__26639;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26604;
    wire N__26603;
    wire N__26602;
    wire N__26601;
    wire N__26600;
    wire N__26599;
    wire N__26596;
    wire N__26595;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26583;
    wire N__26580;
    wire N__26579;
    wire N__26578;
    wire N__26577;
    wire N__26576;
    wire N__26575;
    wire N__26574;
    wire N__26571;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26545;
    wire N__26540;
    wire N__26535;
    wire N__26532;
    wire N__26527;
    wire N__26522;
    wire N__26517;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26494;
    wire N__26491;
    wire N__26476;
    wire N__26475;
    wire N__26474;
    wire N__26471;
    wire N__26470;
    wire N__26469;
    wire N__26468;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26456;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26432;
    wire N__26427;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26412;
    wire N__26411;
    wire N__26408;
    wire N__26405;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26387;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26355;
    wire N__26354;
    wire N__26353;
    wire N__26352;
    wire N__26351;
    wire N__26348;
    wire N__26341;
    wire N__26338;
    wire N__26333;
    wire N__26328;
    wire N__26325;
    wire N__26318;
    wire N__26311;
    wire N__26308;
    wire N__26305;
    wire N__26304;
    wire N__26299;
    wire N__26296;
    wire N__26295;
    wire N__26290;
    wire N__26287;
    wire N__26286;
    wire N__26285;
    wire N__26282;
    wire N__26277;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26263;
    wire N__26260;
    wire N__26259;
    wire N__26254;
    wire N__26251;
    wire N__26250;
    wire N__26249;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26239;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26223;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26211;
    wire N__26210;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26164;
    wire N__26163;
    wire N__26158;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26152;
    wire N__26151;
    wire N__26148;
    wire N__26147;
    wire N__26144;
    wire N__26141;
    wire N__26138;
    wire N__26135;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26070;
    wire N__26069;
    wire N__26068;
    wire N__26065;
    wire N__26060;
    wire N__26057;
    wire N__26050;
    wire N__26049;
    wire N__26048;
    wire N__26047;
    wire N__26046;
    wire N__26043;
    wire N__26038;
    wire N__26037;
    wire N__26036;
    wire N__26031;
    wire N__26026;
    wire N__26021;
    wire N__26018;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26002;
    wire N__26001;
    wire N__25998;
    wire N__25997;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25975;
    wire N__25970;
    wire N__25963;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25942;
    wire N__25939;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25918;
    wire N__25915;
    wire N__25914;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25896;
    wire N__25895;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25883;
    wire N__25876;
    wire N__25873;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25865;
    wire N__25864;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25849;
    wire N__25848;
    wire N__25843;
    wire N__25840;
    wire N__25837;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25817;
    wire N__25814;
    wire N__25809;
    wire N__25804;
    wire N__25801;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25735;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25713;
    wire N__25708;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25669;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25597;
    wire N__25596;
    wire N__25593;
    wire N__25592;
    wire N__25591;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25583;
    wire N__25580;
    wire N__25579;
    wire N__25578;
    wire N__25575;
    wire N__25574;
    wire N__25571;
    wire N__25570;
    wire N__25569;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25558;
    wire N__25557;
    wire N__25554;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25541;
    wire N__25538;
    wire N__25531;
    wire N__25528;
    wire N__25523;
    wire N__25518;
    wire N__25517;
    wire N__25514;
    wire N__25505;
    wire N__25502;
    wire N__25497;
    wire N__25496;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25474;
    wire N__25469;
    wire N__25456;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25431;
    wire N__25428;
    wire N__25427;
    wire N__25426;
    wire N__25423;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25408;
    wire N__25407;
    wire N__25406;
    wire N__25405;
    wire N__25400;
    wire N__25395;
    wire N__25390;
    wire N__25387;
    wire N__25378;
    wire N__25377;
    wire N__25376;
    wire N__25375;
    wire N__25372;
    wire N__25371;
    wire N__25370;
    wire N__25367;
    wire N__25366;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25345;
    wire N__25342;
    wire N__25341;
    wire N__25338;
    wire N__25331;
    wire N__25328;
    wire N__25323;
    wire N__25320;
    wire N__25313;
    wire N__25306;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25285;
    wire N__25282;
    wire N__25279;
    wire N__25276;
    wire N__25273;
    wire N__25272;
    wire N__25271;
    wire N__25270;
    wire N__25269;
    wire N__25268;
    wire N__25267;
    wire N__25266;
    wire N__25263;
    wire N__25252;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25234;
    wire N__25233;
    wire N__25232;
    wire N__25229;
    wire N__25222;
    wire N__25221;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25210;
    wire N__25209;
    wire N__25208;
    wire N__25207;
    wire N__25204;
    wire N__25191;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25173;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25165;
    wire N__25162;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25122;
    wire N__25121;
    wire N__25120;
    wire N__25119;
    wire N__25118;
    wire N__25117;
    wire N__25114;
    wire N__25111;
    wire N__25110;
    wire N__25107;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25099;
    wire N__25098;
    wire N__25097;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25062;
    wire N__25051;
    wire N__25048;
    wire N__25043;
    wire N__25040;
    wire N__25035;
    wire N__25032;
    wire N__25027;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25013;
    wire N__25010;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24961;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24935;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24904;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24859;
    wire N__24856;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24818;
    wire N__24815;
    wire N__24810;
    wire N__24805;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24784;
    wire N__24781;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24741;
    wire N__24738;
    wire N__24735;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24720;
    wire N__24715;
    wire N__24712;
    wire N__24711;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24678;
    wire N__24673;
    wire N__24670;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24658;
    wire N__24655;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24643;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24631;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24619;
    wire N__24616;
    wire N__24615;
    wire N__24612;
    wire N__24609;
    wire N__24604;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24592;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24582;
    wire N__24577;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24547;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24535;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24520;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24492;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24477;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24456;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24442;
    wire N__24439;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24418;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24387;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24366;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24331;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24312;
    wire N__24307;
    wire N__24306;
    wire N__24305;
    wire N__24302;
    wire N__24297;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24235;
    wire N__24234;
    wire N__24233;
    wire N__24230;
    wire N__24229;
    wire N__24228;
    wire N__24221;
    wire N__24218;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24197;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24141;
    wire N__24140;
    wire N__24135;
    wire N__24132;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24088;
    wire N__24085;
    wire N__24084;
    wire N__24083;
    wire N__24082;
    wire N__24079;
    wire N__24074;
    wire N__24071;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24052;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24040;
    wire N__24037;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24019;
    wire N__24018;
    wire N__24015;
    wire N__24010;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23931;
    wire N__23930;
    wire N__23927;
    wire N__23922;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23880;
    wire N__23879;
    wire N__23876;
    wire N__23875;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23859;
    wire N__23856;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23813;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23796;
    wire N__23793;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23786;
    wire N__23783;
    wire N__23778;
    wire N__23775;
    wire N__23770;
    wire N__23765;
    wire N__23762;
    wire N__23761;
    wire N__23760;
    wire N__23759;
    wire N__23758;
    wire N__23757;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23730;
    wire N__23719;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23696;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23685;
    wire N__23682;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23665;
    wire N__23664;
    wire N__23661;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23617;
    wire N__23616;
    wire N__23615;
    wire N__23612;
    wire N__23607;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23578;
    wire N__23577;
    wire N__23576;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23535;
    wire N__23534;
    wire N__23533;
    wire N__23532;
    wire N__23529;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23463;
    wire N__23462;
    wire N__23461;
    wire N__23460;
    wire N__23459;
    wire N__23458;
    wire N__23457;
    wire N__23452;
    wire N__23449;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23427;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23408;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23391;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23366;
    wire N__23361;
    wire N__23358;
    wire N__23353;
    wire N__23350;
    wire N__23347;
    wire N__23346;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23314;
    wire N__23311;
    wire N__23310;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23298;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23286;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23274;
    wire N__23273;
    wire N__23270;
    wire N__23269;
    wire N__23268;
    wire N__23267;
    wire N__23266;
    wire N__23265;
    wire N__23262;
    wire N__23261;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23230;
    wire N__23229;
    wire N__23224;
    wire N__23219;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23172;
    wire N__23167;
    wire N__23166;
    wire N__23163;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23146;
    wire N__23143;
    wire N__23142;
    wire N__23137;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23129;
    wire N__23126;
    wire N__23121;
    wire N__23116;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23088;
    wire N__23085;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23072;
    wire N__23071;
    wire N__23070;
    wire N__23069;
    wire N__23068;
    wire N__23065;
    wire N__23060;
    wire N__23057;
    wire N__23052;
    wire N__23047;
    wire N__23044;
    wire N__23037;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23025;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23013;
    wire N__23012;
    wire N__23011;
    wire N__23010;
    wire N__23009;
    wire N__23008;
    wire N__23007;
    wire N__23006;
    wire N__23005;
    wire N__23004;
    wire N__23003;
    wire N__23002;
    wire N__23001;
    wire N__22994;
    wire N__22987;
    wire N__22978;
    wire N__22969;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22839;
    wire N__22838;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22826;
    wire N__22823;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22782;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22764;
    wire N__22763;
    wire N__22758;
    wire N__22755;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22740;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22716;
    wire N__22711;
    wire N__22708;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22696;
    wire N__22693;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22660;
    wire N__22659;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22602;
    wire N__22601;
    wire N__22600;
    wire N__22593;
    wire N__22590;
    wire N__22585;
    wire N__22584;
    wire N__22581;
    wire N__22580;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22524;
    wire N__22523;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22461;
    wire N__22460;
    wire N__22459;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22441;
    wire N__22438;
    wire N__22437;
    wire N__22434;
    wire N__22433;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22383;
    wire N__22382;
    wire N__22379;
    wire N__22378;
    wire N__22377;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22366;
    wire N__22361;
    wire N__22358;
    wire N__22357;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22343;
    wire N__22342;
    wire N__22339;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22314;
    wire N__22309;
    wire N__22306;
    wire N__22301;
    wire N__22298;
    wire N__22289;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22224;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22179;
    wire N__22176;
    wire N__22175;
    wire N__22172;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22146;
    wire N__22145;
    wire N__22144;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22140;
    wire N__22139;
    wire N__22136;
    wire N__22133;
    wire N__22130;
    wire N__22129;
    wire N__22126;
    wire N__22121;
    wire N__22118;
    wire N__22113;
    wire N__22112;
    wire N__22107;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22095;
    wire N__22094;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22069;
    wire N__22064;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22033;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22014;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22002;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21966;
    wire N__21965;
    wire N__21958;
    wire N__21955;
    wire N__21954;
    wire N__21953;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21926;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21900;
    wire N__21897;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21891;
    wire N__21890;
    wire N__21889;
    wire N__21888;
    wire N__21885;
    wire N__21880;
    wire N__21875;
    wire N__21870;
    wire N__21865;
    wire N__21858;
    wire N__21847;
    wire N__21840;
    wire N__21835;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21810;
    wire N__21809;
    wire N__21808;
    wire N__21807;
    wire N__21806;
    wire N__21805;
    wire N__21804;
    wire N__21803;
    wire N__21802;
    wire N__21801;
    wire N__21800;
    wire N__21797;
    wire N__21796;
    wire N__21793;
    wire N__21788;
    wire N__21785;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21775;
    wire N__21772;
    wire N__21767;
    wire N__21766;
    wire N__21763;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21730;
    wire N__21729;
    wire N__21728;
    wire N__21723;
    wire N__21720;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21694;
    wire N__21689;
    wire N__21684;
    wire N__21681;
    wire N__21676;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21617;
    wire N__21612;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21582;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21567;
    wire N__21566;
    wire N__21563;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21555;
    wire N__21552;
    wire N__21551;
    wire N__21548;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21530;
    wire N__21529;
    wire N__21528;
    wire N__21525;
    wire N__21518;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21493;
    wire N__21492;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21480;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21462;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21450;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21439;
    wire N__21438;
    wire N__21435;
    wire N__21434;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21404;
    wire N__21401;
    wire N__21388;
    wire N__21387;
    wire N__21386;
    wire N__21385;
    wire N__21382;
    wire N__21381;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21369;
    wire N__21362;
    wire N__21361;
    wire N__21360;
    wire N__21359;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21340;
    wire N__21335;
    wire N__21328;
    wire N__21327;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21307;
    wire N__21302;
    wire N__21301;
    wire N__21300;
    wire N__21299;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21280;
    wire N__21279;
    wire N__21278;
    wire N__21275;
    wire N__21268;
    wire N__21267;
    wire N__21264;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21242;
    wire N__21241;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21223;
    wire N__21218;
    wire N__21213;
    wire N__21204;
    wire N__21199;
    wire N__21184;
    wire N__21183;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21169;
    wire N__21166;
    wire N__21163;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21138;
    wire N__21137;
    wire N__21132;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21126;
    wire N__21125;
    wire N__21124;
    wire N__21123;
    wire N__21122;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21110;
    wire N__21109;
    wire N__21108;
    wire N__21107;
    wire N__21106;
    wire N__21105;
    wire N__21104;
    wire N__21103;
    wire N__21102;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21078;
    wire N__21073;
    wire N__21068;
    wire N__21067;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21040;
    wire N__21035;
    wire N__21030;
    wire N__21023;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21003;
    wire N__20986;
    wire N__20985;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20965;
    wire N__20964;
    wire N__20963;
    wire N__20962;
    wire N__20959;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20949;
    wire N__20944;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20921;
    wire N__20920;
    wire N__20919;
    wire N__20914;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20882;
    wire N__20877;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20854;
    wire N__20847;
    wire N__20830;
    wire N__20829;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20814;
    wire N__20813;
    wire N__20812;
    wire N__20811;
    wire N__20810;
    wire N__20809;
    wire N__20808;
    wire N__20807;
    wire N__20806;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20794;
    wire N__20785;
    wire N__20780;
    wire N__20777;
    wire N__20776;
    wire N__20775;
    wire N__20774;
    wire N__20773;
    wire N__20772;
    wire N__20771;
    wire N__20768;
    wire N__20765;
    wire N__20764;
    wire N__20763;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20751;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20722;
    wire N__20713;
    wire N__20710;
    wire N__20695;
    wire N__20694;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20682;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20664;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20607;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20592;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20542;
    wire N__20539;
    wire N__20538;
    wire N__20535;
    wire N__20532;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20484;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20472;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20454;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20436;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20406;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20391;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20328;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20305;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20266;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20213;
    wire N__20212;
    wire N__20211;
    wire N__20208;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20092;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19944;
    wire N__19943;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19861;
    wire N__19858;
    wire N__19857;
    wire N__19856;
    wire N__19853;
    wire N__19852;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19836;
    wire N__19833;
    wire N__19832;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19812;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19711;
    wire N__19708;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19500;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19485;
    wire N__19480;
    wire N__19477;
    wire N__19476;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19448;
    wire N__19443;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19344;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19332;
    wire N__19327;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19314;
    wire N__19313;
    wire N__19310;
    wire N__19307;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19297;
    wire N__19294;
    wire N__19289;
    wire N__19286;
    wire N__19283;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19266;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19201;
    wire N__19200;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19177;
    wire N__19176;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19105;
    wire N__19104;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19078;
    wire N__19075;
    wire N__19074;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19039;
    wire N__19038;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19011;
    wire N__19008;
    wire N__19005;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18987;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18949;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18937;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18922;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18889;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18877;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18862;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18829;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18817;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18802;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18757;
    wire N__18754;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18731;
    wire N__18726;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18685;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18673;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18658;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18646;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18634;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18622;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18607;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18595;
    wire N__18592;
    wire N__18589;
    wire N__18586;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18540;
    wire N__18533;
    wire N__18530;
    wire N__18523;
    wire N__18522;
    wire N__18519;
    wire N__18518;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18467;
    wire N__18466;
    wire N__18465;
    wire N__18462;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18442;
    wire N__18439;
    wire N__18438;
    wire N__18435;
    wire N__18434;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18393;
    wire N__18390;
    wire N__18389;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18267;
    wire N__18264;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18252;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18219;
    wire N__18218;
    wire N__18215;
    wire N__18214;
    wire N__18211;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18193;
    wire N__18192;
    wire N__18189;
    wire N__18188;
    wire N__18185;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18136;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18079;
    wire N__18078;
    wire N__18075;
    wire N__18074;
    wire N__18071;
    wire N__18070;
    wire N__18067;
    wire N__18062;
    wire N__18059;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18033;
    wire N__18030;
    wire N__18029;
    wire N__18026;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18003;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17887;
    wire N__17884;
    wire N__17883;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17872;
    wire N__17869;
    wire N__17862;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17844;
    wire N__17843;
    wire N__17840;
    wire N__17839;
    wire N__17836;
    wire N__17833;
    wire N__17830;
    wire N__17827;
    wire N__17818;
    wire N__17815;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17808;
    wire N__17803;
    wire N__17798;
    wire N__17795;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17731;
    wire N__17728;
    wire N__17727;
    wire N__17724;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17703;
    wire N__17702;
    wire N__17697;
    wire N__17694;
    wire N__17689;
    wire N__17686;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17628;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17604;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17577;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17562;
    wire N__17557;
    wire N__17554;
    wire N__17553;
    wire N__17548;
    wire N__17545;
    wire N__17544;
    wire N__17541;
    wire N__17538;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17526;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17439;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17409;
    wire N__17408;
    wire N__17405;
    wire N__17400;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17310;
    wire N__17309;
    wire N__17306;
    wire N__17301;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17280;
    wire N__17279;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17261;
    wire N__17260;
    wire N__17257;
    wire N__17252;
    wire N__17249;
    wire N__17242;
    wire N__17241;
    wire N__17240;
    wire N__17237;
    wire N__17232;
    wire N__17227;
    wire N__17224;
    wire N__17223;
    wire N__17220;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17212;
    wire N__17209;
    wire N__17204;
    wire N__17201;
    wire N__17194;
    wire N__17193;
    wire N__17192;
    wire N__17189;
    wire N__17184;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17169;
    wire N__17168;
    wire N__17165;
    wire N__17160;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17145;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17106;
    wire N__17105;
    wire N__17104;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17094;
    wire N__17087;
    wire N__17084;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__17001;
    wire N__16998;
    wire N__16997;
    wire N__16990;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16978;
    wire N__16977;
    wire N__16974;
    wire N__16973;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16744;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16693;
    wire N__16690;
    wire N__16689;
    wire N__16684;
    wire N__16681;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16641;
    wire N__16640;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16628;
    wire N__16625;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16585;
    wire N__16582;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16552;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16516;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16483;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16459;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16428;
    wire N__16425;
    wire N__16424;
    wire N__16423;
    wire N__16420;
    wire N__16415;
    wire N__16412;
    wire N__16405;
    wire N__16402;
    wire N__16401;
    wire N__16398;
    wire N__16397;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16376;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16354;
    wire N__16351;
    wire N__16350;
    wire N__16347;
    wire N__16346;
    wire N__16343;
    wire N__16336;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16254;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16243;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16216;
    wire N__16215;
    wire N__16214;
    wire N__16211;
    wire N__16208;
    wire N__16205;
    wire N__16202;
    wire N__16197;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16086;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16071;
    wire N__16068;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16051;
    wire N__16048;
    wire N__16047;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16019;
    wire N__16014;
    wire N__16011;
    wire N__16006;
    wire N__16005;
    wire N__16002;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15975;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15960;
    wire N__15955;
    wire N__15954;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15942;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15918;
    wire N__15913;
    wire N__15912;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15897;
    wire N__15894;
    wire N__15893;
    wire N__15890;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15876;
    wire N__15871;
    wire N__15870;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15855;
    wire N__15852;
    wire N__15851;
    wire N__15850;
    wire N__15849;
    wire N__15848;
    wire N__15847;
    wire N__15846;
    wire N__15845;
    wire N__15844;
    wire N__15843;
    wire N__15842;
    wire N__15841;
    wire N__15840;
    wire N__15839;
    wire N__15838;
    wire N__15837;
    wire N__15830;
    wire N__15821;
    wire N__15814;
    wire N__15807;
    wire N__15798;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15757;
    wire N__15754;
    wire N__15753;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15743;
    wire N__15736;
    wire N__15735;
    wire N__15732;
    wire N__15731;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15715;
    wire N__15712;
    wire N__15711;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15687;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15677;
    wire N__15670;
    wire N__15669;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15654;
    wire N__15649;
    wire N__15646;
    wire N__15645;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15630;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15620;
    wire N__15615;
    wire N__15610;
    wire N__15607;
    wire N__15606;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15579;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15562;
    wire N__15559;
    wire N__15558;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15520;
    wire N__15517;
    wire N__15516;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15480;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15463;
    wire N__15462;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15439;
    wire N__15436;
    wire N__15427;
    wire N__15424;
    wire N__15423;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15408;
    wire N__15403;
    wire N__15402;
    wire N__15399;
    wire N__15394;
    wire N__15391;
    wire N__15388;
    wire N__15387;
    wire N__15384;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15369;
    wire N__15364;
    wire N__15361;
    wire N__15360;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15346;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15330;
    wire N__15327;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15300;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15274;
    wire N__15273;
    wire N__15268;
    wire N__15265;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15253;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15226;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15196;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15184;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15169;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15136;
    wire N__15135;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15121;
    wire N__15118;
    wire N__15117;
    wire N__15116;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15087;
    wire N__15086;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15075;
    wire N__15072;
    wire N__15063;
    wire N__15058;
    wire N__15055;
    wire N__15054;
    wire N__15053;
    wire N__15050;
    wire N__15045;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15027;
    wire N__15024;
    wire N__15023;
    wire N__15022;
    wire N__15021;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15015;
    wire N__15014;
    wire N__15007;
    wire N__15006;
    wire N__15003;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14941;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14929;
    wire N__14928;
    wire N__14925;
    wire N__14924;
    wire N__14923;
    wire N__14918;
    wire N__14915;
    wire N__14908;
    wire N__14907;
    wire N__14900;
    wire N__14891;
    wire N__14884;
    wire N__14881;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14854;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14842;
    wire N__14839;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14824;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14812;
    wire N__14809;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14797;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14782;
    wire N__14779;
    wire N__14776;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14719;
    wire N__14716;
    wire N__14715;
    wire N__14714;
    wire N__14713;
    wire N__14712;
    wire N__14711;
    wire N__14710;
    wire N__14709;
    wire N__14708;
    wire N__14705;
    wire N__14694;
    wire N__14687;
    wire N__14684;
    wire N__14677;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14629;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14617;
    wire N__14614;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14602;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14542;
    wire N__14539;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14473;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14449;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14434;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14305;
    wire N__14302;
    wire N__14299;
    wire N__14296;
    wire N__14293;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14221;
    wire N__14218;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14196;
    wire N__14191;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14167;
    wire N__14164;
    wire N__14163;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14106;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire VCCG0;
    wire bfn_1_1_0_;
    wire \HDA_STRAP.un1_count_1_cry_0 ;
    wire \HDA_STRAP.un1_count_1_cry_1 ;
    wire \HDA_STRAP.un1_count_1_cry_2 ;
    wire \HDA_STRAP.un1_count_1_cry_3 ;
    wire \HDA_STRAP.un1_count_1_cry_4 ;
    wire \HDA_STRAP.un1_count_1_cry_5 ;
    wire \HDA_STRAP.un1_count_1_cry_6 ;
    wire \HDA_STRAP.un1_count_1_cry_7 ;
    wire bfn_1_2_0_;
    wire \HDA_STRAP.un1_count_1_cry_8 ;
    wire \HDA_STRAP.un1_count_1_cry_9 ;
    wire \HDA_STRAP.un1_count_1_cry_10 ;
    wire \HDA_STRAP.un1_count_1_cry_11 ;
    wire \HDA_STRAP.un1_count_1_cry_12 ;
    wire \HDA_STRAP.un1_count_1_cry_13 ;
    wire \HDA_STRAP.un1_count_1_cry_14 ;
    wire \HDA_STRAP.un1_count_1_cry_15 ;
    wire bfn_1_3_0_;
    wire \HDA_STRAP.un1_count_1_cry_16 ;
    wire \HDA_STRAP.curr_state_RNIH91AZ0Z_1 ;
    wire bfn_1_5_0_;
    wire \DSW_PWRGD.un1_count_1_cry_0 ;
    wire \DSW_PWRGD.un1_count_1_cry_1 ;
    wire \DSW_PWRGD.un1_count_1_cry_2 ;
    wire \DSW_PWRGD.un1_count_1_cry_3 ;
    wire \DSW_PWRGD.un1_count_1_cry_4 ;
    wire \DSW_PWRGD.un1_count_1_cry_5 ;
    wire \DSW_PWRGD.un1_count_1_cry_6 ;
    wire \DSW_PWRGD.un1_count_1_cry_7 ;
    wire bfn_1_6_0_;
    wire \DSW_PWRGD.un1_count_1_cry_8 ;
    wire \DSW_PWRGD.un1_count_1_cry_9 ;
    wire \DSW_PWRGD.un1_count_1_cry_10 ;
    wire \DSW_PWRGD.un1_count_1_cry_11 ;
    wire \DSW_PWRGD.un1_count_1_cry_12 ;
    wire \DSW_PWRGD.un1_count_1_cry_13 ;
    wire \DSW_PWRGD.un1_count_1_cry_14 ;
    wire \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_1_7_0_;
    wire \POWERLED.count_0_4 ;
    wire \POWERLED.count_0_13 ;
    wire \POWERLED.count_0_5 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.count_1_1_cascade_ ;
    wire \POWERLED.countZ0Z_1_cascade_ ;
    wire \POWERLED.count_0_1 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.count_0_12 ;
    wire pwrbtn_led;
    wire \POWERLED.curr_state_3_0_cascade_ ;
    wire \POWERLED.curr_stateZ0Z_0_cascade_ ;
    wire \POWERLED.count_0_sqmuxa_i_cascade_ ;
    wire \POWERLED.count_1_0_cascade_ ;
    wire \POWERLED.count_0_0 ;
    wire \POWERLED.pwm_outZ0 ;
    wire \POWERLED.g0_i_o3_0 ;
    wire \POWERLED.un79_clk_100khzlt6_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_5_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_7_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_3 ;
    wire \POWERLED.count_RNIZ0Z_8_cascade_ ;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \POWERLED.N_8 ;
    wire \POWERLED.un1_count_cry_0_i ;
    wire bfn_1_13_0_;
    wire \POWERLED.N_5110_i ;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.N_5111_i ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.N_5112_i ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.N_5113_i ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.N_5114_i ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.N_5115_i ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.N_5116_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.N_5117_i ;
    wire bfn_1_14_0_;
    wire \POWERLED.N_5118_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.N_5119_i ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.N_5120_i ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.N_5121_i ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.N_5122_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.N_5123_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.N_5124_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_1_15_0_;
    wire \POWERLED.mult1_un82_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_5 ;
    wire \POWERLED.un85_clk_100khz_9 ;
    wire \POWERLED.un85_clk_100khz_8 ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_10 ;
    wire \POWERLED.mult1_un89_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_3 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_0 ;
    wire \HDA_STRAP.un4_count_cascade_ ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.countZ0Z_3 ;
    wire \HDA_STRAP.countZ0Z_5 ;
    wire \HDA_STRAP.un4_count_10 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_17 ;
    wire \HDA_STRAP.countZ0Z_1 ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \HDA_STRAP.un4_count_9_cascade_ ;
    wire \HDA_STRAP.un4_count_13 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_16 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_10 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.countZ0Z_9 ;
    wire \HDA_STRAP.countZ0Z_13 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un4_count_11 ;
    wire \HDA_STRAP.countZ0Z_15 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.un4_count_12 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_6 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_8 ;
    wire \HDA_STRAP.countZ0Z_8 ;
    wire \HDA_STRAP.count_RNO_0Z0Z_11 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.N_14_cascade_ ;
    wire \HDA_STRAP.un4_count ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire hda_sdo_atp;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_ ;
    wire \HDA_STRAP.curr_state_RNO_0Z0Z_0 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.N_5_0 ;
    wire \DSW_PWRGD.countZ0Z_14 ;
    wire \DSW_PWRGD.countZ0Z_13 ;
    wire \DSW_PWRGD.countZ0Z_15 ;
    wire \DSW_PWRGD.countZ0Z_12 ;
    wire \DSW_PWRGD.un4_count_9_cascade_ ;
    wire \DSW_PWRGD.countZ0Z_2 ;
    wire \DSW_PWRGD.countZ0Z_5 ;
    wire \DSW_PWRGD.countZ0Z_7 ;
    wire \DSW_PWRGD.countZ0Z_3 ;
    wire \DSW_PWRGD.un4_count_10 ;
    wire \DSW_PWRGD.countZ0Z_11 ;
    wire \DSW_PWRGD.countZ0Z_10 ;
    wire \DSW_PWRGD.countZ0Z_8 ;
    wire \DSW_PWRGD.countZ0Z_0 ;
    wire \DSW_PWRGD.un4_count_11 ;
    wire \DSW_PWRGD.un1_curr_state10_0 ;
    wire \DSW_PWRGD.curr_stateZ0Z_1 ;
    wire v33dsw_ok;
    wire \DSW_PWRGD.curr_stateZ0Z_0 ;
    wire \DSW_PWRGD.N_1_i ;
    wire DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_;
    wire G_27;
    wire G_27_cascade_;
    wire \DSW_PWRGD.N_29_1 ;
    wire \POWERLED.d_i1_mux_cascade_ ;
    wire \POWERLED.dutycycle_RNI_16Z0Z_9_cascade_ ;
    wire \POWERLED.d_i3_mux_cascade_ ;
    wire \POWERLED.un1_i3_mux ;
    wire \POWERLED.dutycycle_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_3_1 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_ ;
    wire \POWERLED.count_0_10 ;
    wire \POWERLED.count_0_2 ;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.countZ0Z_0 ;
    wire bfn_2_10_0_;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.count_1_2 ;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.count_1_3 ;
    wire \POWERLED.un1_count_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.count_1_4 ;
    wire \POWERLED.un1_count_cry_3 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.count_1_5 ;
    wire \POWERLED.un1_count_cry_4 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire bfn_2_11_0_;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.count_1_10 ;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.count_1_11 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.count_1_12 ;
    wire \POWERLED.un1_count_cry_11_cZ0 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.count_1_13 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ;
    wire \POWERLED.un1_count_cry_13_cZ0 ;
    wire \POWERLED.count_0_sqmuxa_i ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.count_1_9 ;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.count_1_6 ;
    wire \POWERLED.count_0_6 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ;
    wire \POWERLED.count_0_15 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.count_1_7 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.count_1_8 ;
    wire \POWERLED.count_0_8 ;
    wire bfn_2_13_0_;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8_cascade_ ;
    wire \POWERLED.un85_clk_100khz_7 ;
    wire bfn_2_14_0_;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire bfn_2_15_0_;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire bfn_2_16_0_;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_2_c ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_3_c ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_4_c ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_cry_5_c ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6_c ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.count_off_0_8 ;
    wire \POWERLED.count_offZ0Z_8_cascade_ ;
    wire \POWERLED.count_off_0_3 ;
    wire \POWERLED.count_off_0_7 ;
    wire \DSW_PWRGD.countZ0Z_1 ;
    wire \DSW_PWRGD.countZ0Z_6 ;
    wire \DSW_PWRGD.countZ0Z_9 ;
    wire \DSW_PWRGD.countZ0Z_4 ;
    wire \DSW_PWRGD.un4_count_8 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_3_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_20_0_0 ;
    wire \POWERLED.o2_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_7_1 ;
    wire \POWERLED.un1_dutycycle_53_axb_7_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_10 ;
    wire \POWERLED.un1_dutycycle_53_axb_4_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_8_2_0 ;
    wire \POWERLED.un1_dutycycle_53_8_2_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_8_5_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_12_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_8_3 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_3 ;
    wire \POWERLED.un1_dutycycle_53_56_a0_1 ;
    wire \POWERLED.un1_dutycycle_53_56_a1_1 ;
    wire \POWERLED.un1_clk_100khz_45_and_i_i_a3_0_0_cascade_ ;
    wire \POWERLED.N_4_cascade_ ;
    wire \POWERLED.dutycycle_eena_3_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_3 ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \POWERLED.dutycycle_eena_3_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_2_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_4_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_4_3_1 ;
    wire \POWERLED.un2_count_clk_17_0_a2_1_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_a2_5_cascade_ ;
    wire bfn_4_10_0_;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire v5s_enn;
    wire \POWERLED.mult1_un47_sum_i ;
    wire \POWERLED.mult1_un103_sum_i ;
    wire v33a_enn;
    wire \POWERLED.un85_clk_100khz_6 ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire bfn_4_13_0_;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire bfn_4_14_0_;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_7_l_fx ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire vpp_ok;
    wire vddq_en;
    wire \POWERLED.mult1_un75_sum_i_8 ;
    wire bfn_4_16_0_;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire bfn_5_1_0_;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_5_2_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_5_3_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_5_4_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \POWERLED.count_off_0_9 ;
    wire \POWERLED.count_offZ0Z_9_cascade_ ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_off_0_11 ;
    wire \POWERLED.dutycycle_eena_8_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_8_cascade_ ;
    wire \POWERLED.dutycycle_eena_8 ;
    wire \POWERLED.dutycycleZ1Z_3 ;
    wire \POWERLED.dutycycleZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_eena_4_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_4 ;
    wire \POWERLED.dutycycle_eena_4_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \POWERLED.dutycycle_eena_5_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_5_cascade_ ;
    wire \POWERLED.dutycycle_eena_5_1 ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \POWERLED.dutycycle_eena_6_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_6 ;
    wire \POWERLED.dutycycle_eena_6_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire \POWERLED.dutycycle_eena_5 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.N_4_0_cascade_ ;
    wire \POWERLED.dutycycle_en_12_cascade_ ;
    wire \POWERLED.un1_clk_100khz_48_and_i_i_a3_0_0 ;
    wire \POWERLED.dutycycle_en_12 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.dutycycleZ0Z_13_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_12_cascade_ ;
    wire bfn_5_9_0_;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un47_sum_cry_5_THRU_CO ;
    wire \POWERLED.un1_dutycycle_53_4_3 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.count_RNIZ0Z_8 ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.curr_state_1_0 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_10 ;
    wire \POWERLED.dutycycle_RNI_9Z0Z_9 ;
    wire \POWERLED.mult1_un40_sum_i_5 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_s_6 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire \POWERLED.mult1_un47_sum_s_4_sf ;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire bfn_5_11_0_;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8_cascade_ ;
    wire bfn_5_12_0_;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire bfn_5_13_0_;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire bfn_5_14_0_;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire bfn_5_15_0_;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8_cascade_ ;
    wire \POWERLED.un85_clk_100khz_4 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_6_2_0_;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire COUNTER_un4_counter_7;
    wire bfn_6_3_0_;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.un4_counter_4_and ;
    wire pch_pwrok;
    wire vccst_pwrgd;
    wire bfn_6_4_0_;
    wire \POWERLED.un3_count_off_1_cry_1 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.count_off_1_8 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_off_1_9 ;
    wire bfn_6_5_0_;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_off_1_10 ;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.count_off_1_12 ;
    wire \POWERLED.count_off_0_12 ;
    wire \POWERLED.dutycycleZ1Z_14 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_13Z0Z_9 ;
    wire \POWERLED.un1_dutycycle_53_2_0 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_11_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_4 ;
    wire \POWERLED.dutycycle_en_7_cascade_ ;
    wire \POWERLED.un1_clk_100khz_39_and_i_0_0 ;
    wire \POWERLED.un1_clk_100khz_30_and_i_0_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI4J2O7Z0Z_9 ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.dutycycle_RNI4J2O7Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_11 ;
    wire \POWERLED.dutycycle_en_7 ;
    wire \POWERLED.un1_dutycycle_53_20_1 ;
    wire \POWERLED.un1_dutycycle_53_3_2_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_3_2_cascade_ ;
    wire \POWERLED.dutycycle_en_10 ;
    wire \POWERLED.dutycycleZ1Z_13 ;
    wire \POWERLED.un1_dutycycle_53_50_0 ;
    wire \POWERLED.dutycycle_RNI_12Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_15Z0Z_9 ;
    wire \POWERLED.dutycycle_RNI_11Z0Z_9 ;
    wire bfn_6_9_0_;
    wire \POWERLED.dutycycle_RNI_1Z0Z_0 ;
    wire \POWERLED.un1_dutycycle_53_cry_0_cZ0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_2 ;
    wire \POWERLED.un1_dutycycle_53_cry_1_cZ0 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_2 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_2_cZ0 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_3 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_3 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_3_cZ0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_4 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_4_cZ0 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_9 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_5_cZ0 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_10 ;
    wire \POWERLED.un1_dutycycle_53_cry_6 ;
    wire \POWERLED.un1_dutycycle_53_cry_7 ;
    wire \POWERLED.dutycycle_RNIZ0Z_11 ;
    wire bfn_6_10_0_;
    wire \POWERLED.dutycycle_RNI_1Z0Z_12 ;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_8 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_9 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.dutycycle_RNIZ0Z_15 ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.mult1_un47_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire bfn_6_11_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.g2_1 ;
    wire \POWERLED.g2_5 ;
    wire \POWERLED.g0_4_4 ;
    wire \POWERLED.g0_4_5_cascade_ ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.g3_1_0 ;
    wire \POWERLED.g3_1_4_cascade_ ;
    wire \POWERLED.g3_1_6_cascade_ ;
    wire \POWERLED.un2_count_clk_17_0_a2_5 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_i_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un85_clk_100khz_2 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un145_sum ;
    wire bfn_6_14_0_;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un89_sum ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \PCH_PWRGD.count_0_15 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \PCH_PWRGD.countZ0Z_15_cascade_ ;
    wire \PCH_PWRGD.count_rst_10_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_4_cascade_ ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.countZ0Z_14_cascade_ ;
    wire \PCH_PWRGD.count_0_12 ;
    wire PCH_PWRGD_delayed_vccin_ok;
    wire \PCH_PWRGD.N_250_0 ;
    wire \PCH_PWRGD.N_250_0_cascade_ ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \POWERLED.dutycycleZ0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.dutycycle_eena_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.dutycycle_1_0_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_0 ;
    wire \POWERLED.dutycycle_1_0_1 ;
    wire \POWERLED.dutycycleZ1Z_1 ;
    wire \POWERLED.dutycycle_eena_0_cascade_ ;
    wire \POWERLED.dutycycle_1_0_0 ;
    wire \POWERLED.func_state_RNISKPU6Z0Z_0_cascade_ ;
    wire \POWERLED.count_off_1_13 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_off_1_14 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2 ;
    wire \POWERLED.count_off_0_15 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_15_cascade_ ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.dutycycleZ1Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_96_0_a3_0 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_0 ;
    wire \POWERLED.un2_count_clk_17_0_cascade_ ;
    wire bfn_7_7_0_;
    wire \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_cZ0 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI765BZ0Z1 ;
    wire \POWERLED.un1_dutycycle_94_cry_2 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI886BZ0Z1 ;
    wire \POWERLED.un1_dutycycle_94_cry_3 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.dutycycleZ1Z_5 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4AZ0Z1 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNICGABZ0Z1 ;
    wire bfn_7_8_0_;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ;
    wire \POWERLED.un1_dutycycle_94_cry_8_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCBZ0Z1 ;
    wire \POWERLED.un1_dutycycle_94_cry_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_11 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_12 ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_11 ;
    wire \POWERLED.N_115_f0_1 ;
    wire \POWERLED.N_366_cascade_ ;
    wire \POWERLED.dutycycle_RNI2O4A1Z0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI2O4A1_2Z0Z_2 ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m1_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_5 ;
    wire \POWERLED.func_state_RNI_0Z0Z_0_cascade_ ;
    wire \POWERLED.func_state_RNI68EU3Z0Z_1 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ;
    wire \POWERLED.dutycycle_1_0_iv_0_1_5_cascade_ ;
    wire SUSWARN_N_fast;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.m18_e_0 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_c_RNI919HZ0Z1 ;
    wire \POWERLED.dutycycle_1_0_5_cascade_ ;
    wire \POWERLED.func_state_RNIT69J5Z0Z_1 ;
    wire G_155_cascade_;
    wire \POWERLED.N_73 ;
    wire \POWERLED.dutycycle_eena_1 ;
    wire \POWERLED.N_73_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire \POWERLED.N_277 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_2 ;
    wire bfn_7_13_0_;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire bfn_7_14_0_;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7_cascade_ ;
    wire \POWERLED.un85_clk_100khz_1 ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire bfn_7_15_0_;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_2078;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un85_clk_100khz_0 ;
    wire G_9;
    wire bfn_8_1_0_;
    wire \PCH_PWRGD.un2_count_1_axb_2 ;
    wire \PCH_PWRGD.count_rst_12 ;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.un2_count_1_axb_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire bfn_8_2_0_;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.un2_count_1_axb_13 ;
    wire \PCH_PWRGD.count_rst_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.count_rst ;
    wire bfn_8_3_0_;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire bfn_8_4_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_5_0_;
    wire \POWERLED.count_off_RNIBQDB2Z0Z_0_cascade_ ;
    wire \POWERLED.count_offZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_off_0_0 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.count_off_RNIZ0Z_1 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.count_offZ0Z_1_cascade_ ;
    wire \POWERLED.un34_clk_100khz_10 ;
    wire \POWERLED.un34_clk_100khz_8 ;
    wire \POWERLED.un34_clk_100khz_9_cascade_ ;
    wire \POWERLED.un34_clk_100khz_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ;
    wire \POWERLED.N_220_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823 ;
    wire \POWERLED.N_304_cascade_ ;
    wire \POWERLED.N_2216_i_cascade_ ;
    wire \POWERLED.func_state_1_m2s2_i_1_cascade_ ;
    wire \POWERLED.N_160 ;
    wire \POWERLED.N_3_0 ;
    wire slp_s3n_signal_cascade_;
    wire \POWERLED.N_183 ;
    wire \POWERLED.func_state_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.N_162_i ;
    wire \POWERLED.N_335 ;
    wire \POWERLED.func_state_RNI2O4A1Z0Z_1_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.dutycycle_en_9 ;
    wire \POWERLED.func_state_RNI2O4A1_1Z0Z_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.dutycycleZ0Z_11_cascade_ ;
    wire \POWERLED.un1_clk_100khz_42_and_i_0_0 ;
    wire \POWERLED.func_state_RNI2O4A1Z0Z_1 ;
    wire \POWERLED.un1_clk_100khz_47_and_i_0_0_cascade_ ;
    wire \POWERLED.N_399_N ;
    wire \POWERLED.dutycycle_en_11 ;
    wire \POWERLED.m18_e_5 ;
    wire \POWERLED.m18_e_6 ;
    wire \POWERLED.func_m2_0_a2Z0Z_0 ;
    wire \POWERLED.func_m2_0_a2Z0Z_0_cascade_ ;
    wire \POWERLED.count_clk_RNI2O4A1_0Z0Z_10 ;
    wire \POWERLED.func_state_RNI91IA4_0Z0Z_1_cascade_ ;
    wire \POWERLED.func_state_1_m2_0 ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \POWERLED.func_state_1_m2_0_cascade_ ;
    wire \POWERLED.g0_9_1_cascade_ ;
    wire \POWERLED.dutycycle_fb_15_4_0_cascade_ ;
    wire \POWERLED.dutycycle_fb_15_0 ;
    wire \POWERLED.dutycycle_en_14_cascade_ ;
    wire \POWERLED.func_m2_0_a2_isoZ0 ;
    wire \POWERLED.dutycycle_eena_14_0Z0Z_0 ;
    wire \POWERLED.dutycycle_fb_15_1 ;
    wire \POWERLED.g1_0 ;
    wire \POWERLED.g1 ;
    wire \POWERLED.dutycycle_fb_15_2_0 ;
    wire SUSWARN_N_rep1;
    wire \POWERLED.N_340_cascade_ ;
    wire \POWERLED.func_state_RNIRAVV2Z0Z_0 ;
    wire \POWERLED.dutycycle_1_0_5 ;
    wire \POWERLED.dutycycle_fb_15_1_1 ;
    wire \POWERLED.g2_0 ;
    wire \POWERLED.N_398_0 ;
    wire \POWERLED.g0_1_0 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_10 ;
    wire \POWERLED.func_state_1_m2s2_i_a3_0 ;
    wire \POWERLED.dutycycle_0_5 ;
    wire \POWERLED.dutycycle_fb_14_a4_1 ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.count_off_1_sqmuxa ;
    wire \POWERLED.count_off_1_sqmuxa_cascade_ ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_6 ;
    wire \POWERLED.N_325 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_0 ;
    wire \POWERLED.dutycycle_RNINH5P1Z0Z_2 ;
    wire \POWERLED.dutycycle_RNI4G9K2Z0Z_5 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_0_cascade_ ;
    wire \POWERLED.dutycycle_RNO_2Z0Z_5_cascade_ ;
    wire \POWERLED.N_240 ;
    wire \POWERLED.dutycycle_eena_13 ;
    wire \POWERLED.un2_count_clk_17_0_0 ;
    wire \POWERLED.g3 ;
    wire \POWERLED.un1_dutycycle_172_m3_1_0_cascade_ ;
    wire \POWERLED.dutycycle_RNO_3Z0Z_5 ;
    wire \POWERLED.dutycycle_RNIZ0Z_6 ;
    wire \POWERLED.un1_dutycycle_172_m3s4_1 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_6 ;
    wire \POWERLED.N_239 ;
    wire \POWERLED.func_state_RNI_0Z0Z_0 ;
    wire \POWERLED.N_271 ;
    wire \POWERLED.N_366 ;
    wire \POWERLED.N_331 ;
    wire \POWERLED.N_272 ;
    wire \POWERLED.dutycycle_N_3_mux_0_0 ;
    wire \PCH_PWRGD.count_rst_10 ;
    wire \PCH_PWRGD.count_0_4 ;
    wire \PCH_PWRGD.count_rst_11_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.countZ0Z_3_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_8_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.un2_count_1_axb_10 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.countZ0Z_6_cascade_ ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.count_1_i_a2_1_0 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.count_1_i_a2_0_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_2_0 ;
    wire \PCH_PWRGD.count_1_i_a2_11_0_cascade_ ;
    wire \PCH_PWRGD.count_rst_3_cascade_ ;
    wire N_253_cascade_;
    wire \PCH_PWRGD.count_0_0 ;
    wire \PCH_PWRGD.count_RNIM6A821Z0Z_1 ;
    wire \PCH_PWRGD.countZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_2173_i ;
    wire \PCH_PWRGD.count_1_i_a2_11_0 ;
    wire \PCH_PWRGD.N_2173_i_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.m4_0_a2_11_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.m4_0_a2_10 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.m4_0_a2_9 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.m4_0_a2_0 ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire \RSMRST_PWRGD.m4_0_a2_12 ;
    wire \VPP_VDDQ.count_2_1_10_cascade_ ;
    wire \PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0 ;
    wire \PCH_PWRGD.curr_state_0_0 ;
    wire \PCH_PWRGD.m4_0_cascade_ ;
    wire \VPP_VDDQ.count_2_1_8_cascade_ ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.count_2_1_9_cascade_ ;
    wire \VPP_VDDQ.count_2_0_10 ;
    wire v33a_ok;
    wire v5a_ok;
    wire slp_susn;
    wire v1p8a_ok;
    wire rsmrst_pwrgd_signal_cascade_;
    wire \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ;
    wire N_382;
    wire \RSMRST_PWRGD.N_254_i ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire RSMRST_PWRGD_curr_state_0;
    wire \POWERLED.N_301 ;
    wire G_11;
    wire \RSMRST_PWRGD.N_29_2 ;
    wire COUNTER_un4_counter_7_THRU_CO;
    wire \POWERLED.dutycycle_N_3_mux_0 ;
    wire \POWERLED.count_clk_0_7 ;
    wire \POWERLED.count_clk_0_9 ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_1_5 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_off_0_6 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.count_off_0_2 ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.func_state_RNISKPU6Z0Z_0 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_13 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_15 ;
    wire RSMRSTn_rep1;
    wire \POWERLED.N_4_0_3 ;
    wire \POWERLED.func_state_RNIOGRSZ0Z_0 ;
    wire \POWERLED.func_state_1_ss0_i_0_o2_1 ;
    wire \POWERLED.N_76 ;
    wire \POWERLED.func_state_RNI91IA4Z0Z_1_cascade_ ;
    wire \POWERLED.func_state_1_m2_1 ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.func_state_1_m2_1_cascade_ ;
    wire \POWERLED.func_state_enZ0 ;
    wire \POWERLED.un1_N_3_mux_0 ;
    wire N_4_1_cascade_;
    wire G_34_0_a4_0_2_cascade_;
    wire POWERLED_un1_dutycycle_172_m3_0_0;
    wire \POWERLED.N_8_0 ;
    wire \POWERLED.un1_dutycycle_172_m1_ns_1 ;
    wire \POWERLED.dutycycle_RNI_10Z0Z_3 ;
    wire N_11;
    wire \POWERLED.N_319_0 ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.N_297 ;
    wire \POWERLED.un1_func_state25_6_0_a2_1 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_296_N_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_1_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_2 ;
    wire \POWERLED.N_340 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_ ;
    wire \POWERLED.N_284 ;
    wire \POWERLED.func_state_RNIBQDB2Z0Z_0 ;
    wire \POWERLED.N_340_N ;
    wire \POWERLED.func_state_RNI_1Z0Z_0 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_294_N ;
    wire \POWERLED.func_state_1_m2_am_1_1 ;
    wire \POWERLED.func_N_5_mux_0 ;
    wire \POWERLED.func_state_RNIBL3Q3Z0Z_1 ;
    wire \POWERLED.func_state_1_m2s2_i_a2_0_0 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire func_state_RNI_7_1;
    wire N_7;
    wire rsmrstn;
    wire \POWERLED.func_state_RNIZ0Z_1 ;
    wire slp_s3n;
    wire \POWERLED.un1_clk_100khz_51_and_i_a2_6_0_cascade_ ;
    wire \POWERLED.un1_clk_100khz_51_and_i_a2_6_sx_cascade_ ;
    wire \POWERLED.func_state_RNIPUGO_0Z0Z_1_cascade_ ;
    wire \POWERLED.N_309_N ;
    wire \POWERLED.count_clk_RNI2O4A1Z0Z_10 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_o2_4_1_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.N_145_N ;
    wire \POWERLED.un1_clk_100khz_51_and_i_a2_5_0 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_a2_5_0_cascade_ ;
    wire RSMRSTn_fast;
    wire \POWERLED.func_state_RNIPUGOZ0Z_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_1_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire \PCH_PWRGD.count_rst_13 ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \PCH_PWRGD.count_rst_13_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_6_0 ;
    wire \PCH_PWRGD.count_1_i_a2_3_0_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_12_0 ;
    wire \PCH_PWRGD.un2_count_1_axb_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_axb_9_cascade_ ;
    wire \PCH_PWRGD.count_rst_5 ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.countZ0Z_8 ;
    wire \PCH_PWRGD.count_rst_5_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_4_0 ;
    wire \PCH_PWRGD.count_rst_7 ;
    wire \PCH_PWRGD.count_rst_7_cascade_ ;
    wire \PCH_PWRGD.count_1_i_a2_5_0 ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_axb_7 ;
    wire \PCH_PWRGD.count_0_7 ;
    wire \PCH_PWRGD.count_rst_9_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_5_cascade_ ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_11 ;
    wire \PCH_PWRGD.count_0_11 ;
    wire \PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ;
    wire \PCH_PWRGD.N_364 ;
    wire G_1939_cascade_;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire N_218;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire G_1939;
    wire N_218_cascade_;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire \PCH_PWRGD.curr_state_0_1_cascade_ ;
    wire \PCH_PWRGD.N_2190_i ;
    wire \PCH_PWRGD.N_2171_i ;
    wire \PCH_PWRGD.N_2190_i_cascade_ ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire \VPP_VDDQ.N_53_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_0_1 ;
    wire \VPP_VDDQ.N_55_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2_1_3_cascade_ ;
    wire \VPP_VDDQ.count_2_1_2_cascade_ ;
    wire \VPP_VDDQ.count_2_0_2 ;
    wire \VPP_VDDQ.count_2Z0Z_2_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire bfn_11_6_0_;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ;
    wire bfn_11_7_0_;
    wire \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ;
    wire \VPP_VDDQ.count_2_1_7_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.un9_clk_100khz_7_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire \VPP_VDDQ.count_2_1_7 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.count_2_1_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.count_clkZ0Z_14_cascade_ ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.count_clk_0_14 ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ;
    wire \POWERLED.count_clkZ0Z_0_cascade_ ;
    wire \POWERLED.count_clk_RNIZ0Z_0_cascade_ ;
    wire \POWERLED.count_clk_0_4 ;
    wire \POWERLED.count_clk_0_6 ;
    wire \POWERLED.count_clk_0_0 ;
    wire \POWERLED.count_clk_RNIZ0Z_1 ;
    wire \POWERLED.count_clk_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.count_clk_RNI_0Z0Z_1 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_a2_0_0_cascade_ ;
    wire \POWERLED.N_285 ;
    wire \POWERLED.N_177 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_1_cascade_ ;
    wire gpio_fpga_soc_4;
    wire slp_s4n;
    wire \POWERLED.un1_func_state25_4_i_a2_0_cascade_ ;
    wire \POWERLED.func_state_RNIBVNSZ0Z_0 ;
    wire \POWERLED.N_291 ;
    wire \POWERLED.count_clk_en_0_cascade_ ;
    wire \POWERLED.N_396 ;
    wire \POWERLED.func_state_RNI2O4A1_1Z0Z_1 ;
    wire \POWERLED.count_clk_en_2_cascade_ ;
    wire G_155;
    wire \POWERLED.func_state_RNI_2Z0Z_1 ;
    wire \POWERLED.count_off_RNI_0Z0Z_10 ;
    wire \POWERLED.N_176 ;
    wire \POWERLED.N_176_cascade_ ;
    wire \POWERLED.N_2218_i ;
    wire \POWERLED.N_2216_i ;
    wire \POWERLED.N_27 ;
    wire \POWERLED.func_state ;
    wire \POWERLED.N_219 ;
    wire vpp_en;
    wire \VPP_VDDQ.N_64_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire \VPP_VDDQ.curr_state_7_0 ;
    wire \VPP_VDDQ.curr_state_7_0_cascade_ ;
    wire N_246;
    wire N_246_cascade_;
    wire N_381;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire vccst_en;
    wire \VPP_VDDQ.curr_stateZ0Z_0 ;
    wire \VPP_VDDQ.un6_count_10_cascade_ ;
    wire VPP_VDDQ_un6_count;
    wire \VPP_VDDQ.un6_count_8 ;
    wire \VPP_VDDQ.un6_count_11 ;
    wire \VPP_VDDQ.un6_count_9 ;
    wire suswarn_n;
    wire \VPP_VDDQ.N_361_0_cascade_ ;
    wire \VPP_VDDQ.N_62_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_ok_en_cascade_ ;
    wire VPP_VDDQ_delayed_vddq_ok;
    wire vddq_ok;
    wire \VPP_VDDQ.delayed_vddq_ok_en ;
    wire \VPP_VDDQ.delayed_vddq_okZ0 ;
    wire \VPP_VDDQ.N_361_0 ;
    wire N_570_g;
    wire \VPP_VDDQ.N_2192_i ;
    wire \VPP_VDDQ.N_62 ;
    wire \VPP_VDDQ.N_62_i ;
    wire \VPP_VDDQ.count_2_1_14_cascade_ ;
    wire \VPP_VDDQ.count_2_1_4_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ;
    wire \VPP_VDDQ.count_2_0_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ;
    wire \VPP_VDDQ.count_2_0_5 ;
    wire \VPP_VDDQ.count_2_1_5_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.N_174 ;
    wire dsw_pwrok;
    wire vccst_cpu_ok;
    wire v5s_ok;
    wire v33s_ok;
    wire slp_s3n_signal;
    wire \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ;
    wire rsmrst_pwrgd_signal;
    wire vccin_en;
    wire \VPP_VDDQ.un1_count_2_1_axb_6 ;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \VPP_VDDQ.count_2_1_6 ;
    wire \VPP_VDDQ.un9_clk_100khz_9 ;
    wire \VPP_VDDQ.un9_clk_100khz_0_cascade_ ;
    wire \VPP_VDDQ.un9_clk_100khz_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ;
    wire \VPP_VDDQ.N_1_i_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.count_2_1_12 ;
    wire \VPP_VDDQ.count_2_1_13 ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \VPP_VDDQ.count_2Z0Z_13_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.un9_clk_100khz_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ;
    wire \VPP_VDDQ.count_2_0_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ;
    wire \VPP_VDDQ.count_2_0_14 ;
    wire \VPP_VDDQ.un9_clk_100khz_1 ;
    wire \VPP_VDDQ.count_2_1_1 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_1_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1 ;
    wire \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire \VPP_VDDQ.count_2_1_11_cascade_ ;
    wire \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire bfn_12_9_0_;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ;
    wire bfn_12_10_0_;
    wire \POWERLED.un1_count_clk_2_cry_9 ;
    wire \POWERLED.un1_count_clk_2_cry_10 ;
    wire \POWERLED.un1_count_clk_2_cry_11 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_12 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_13 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.count_clkZ0Z_15_cascade_ ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.count_clk_0_10 ;
    wire \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.count_clkZ0Z_10_cascade_ ;
    wire \POWERLED.count_clk_RNIZ0Z_13 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_cascade_ ;
    wire \POWERLED.N_352 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.un2_count_clk_15_0_9_cascade_ ;
    wire \POWERLED.un2_count_clk_15_0_8 ;
    wire \POWERLED.un2_count_clk_15_1 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.un2_count_clk_15_0_10 ;
    wire \POWERLED.count_clk_0_12 ;
    wire \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.count_clkZ0Z_12_cascade_ ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.count_clk_RNIZ0Z_12_cascade_ ;
    wire \POWERLED.un2_count_clk_15_0_7 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.count_clk_RNIZ0Z_12 ;
    wire \POWERLED.count_clkZ0Z_2_cascade_ ;
    wire \POWERLED.count_clk_RNIZ0Z_15 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1 ;
    wire \POWERLED.func_state_RNIH9594_0_1 ;
    wire \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.count_clk_en ;
    wire \VPP_VDDQ.N_66_i ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire bfn_12_14_0_;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire bfn_12_15_0_;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire N_29_g;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_12_16_0_;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire _gnd_net_;
    wire fpga_osc;
    wire \VPP_VDDQ.N_29_0 ;
    wire G_43;

    defparam ipInertedIOPad_VR_READY_VCCINAUX_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__35432),
            .DIN(N__35431),
            .DOUT(N__35430),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__35432),
            .PADOUT(N__35431),
            .PADIN(N__35430),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__35423),
            .DIN(N__35422),
            .DOUT(N__35421),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__35423),
            .PADOUT(N__35422),
            .PADIN(N__35421),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16753),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__35414),
            .DIN(N__35413),
            .DOUT(N__35412),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__35414),
            .PADOUT(N__35413),
            .PADIN(N__35412),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24942),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__35405),
            .DIN(N__35404),
            .DOUT(N__35403),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__35405),
            .PADOUT(N__35404),
            .PADIN(N__35403),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17059),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__35396),
            .DIN(N__35395),
            .DOUT(N__35394),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__35396),
            .PADOUT(N__35395),
            .PADIN(N__35394),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__35387),
            .DIN(N__35386),
            .DOUT(N__35385),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__35387),
            .PADOUT(N__35386),
            .PADIN(N__35385),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__35378),
            .DIN(N__35377),
            .DOUT(N__35376),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__35378),
            .PADOUT(N__35377),
            .PADIN(N__35376),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__35369),
            .DIN(N__35368),
            .DOUT(N__35367),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__35369),
            .PADOUT(N__35368),
            .PADIN(N__35367),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__35360),
            .DIN(N__35359),
            .DOUT(N__35358),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__35360),
            .PADOUT(N__35359),
            .PADIN(N__35358),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16791),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__35351),
            .DIN(N__35350),
            .DOUT(N__35349),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__35351),
            .PADOUT(N__35350),
            .PADIN(N__35349),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__35342),
            .DIN(N__35341),
            .DOUT(N__35340),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__35342),
            .PADOUT(N__35341),
            .PADIN(N__35340),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__35333),
            .DIN(N__35332),
            .DOUT(N__35331),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__35333),
            .PADOUT(N__35332),
            .PADIN(N__35331),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14140),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__35324),
            .DIN(N__35323),
            .DOUT(N__35322),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__35324),
            .PADOUT(N__35323),
            .PADIN(N__35322),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__35315),
            .DIN(N__35314),
            .DOUT(N__35313),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__35315),
            .PADOUT(N__35314),
            .PADIN(N__35313),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__35306),
            .DIN(N__35305),
            .DOUT(N__35304),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__35306),
            .PADOUT(N__35305),
            .PADIN(N__35304),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__35297),
            .DIN(N__35296),
            .DOUT(N__35295),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__35297),
            .PADOUT(N__35296),
            .PADIN(N__35295),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__35288),
            .DIN(N__35287),
            .DOUT(N__35286),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__35288),
            .PADOUT(N__35287),
            .PADIN(N__35286),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30212),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__35279),
            .DIN(N__35278),
            .DOUT(N__35277),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__35279),
            .PADOUT(N__35278),
            .PADIN(N__35277),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__35270),
            .DIN(N__35269),
            .DOUT(N__35268),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__35270),
            .PADOUT(N__35269),
            .PADIN(N__35268),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__35261),
            .DIN(N__35260),
            .DOUT(N__35259),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__35261),
            .PADOUT(N__35260),
            .PADIN(N__35259),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30637),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__35252),
            .DIN(N__35251),
            .DOUT(N__35250),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__35252),
            .PADOUT(N__35251),
            .PADIN(N__35250),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__35243),
            .DIN(N__35242),
            .DOUT(N__35241),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__35243),
            .PADOUT(N__35242),
            .PADIN(N__35241),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__35234),
            .DIN(N__35233),
            .DOUT(N__35232),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__35234),
            .PADOUT(N__35233),
            .PADIN(N__35232),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__35225),
            .DIN(N__35224),
            .DOUT(N__35223),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__35225),
            .PADOUT(N__35224),
            .PADIN(N__35223),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__35216),
            .DIN(N__35215),
            .DOUT(N__35214),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__35216),
            .PADOUT(N__35215),
            .PADIN(N__35214),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26413),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__35207),
            .DIN(N__35206),
            .DOUT(N__35205),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__35207),
            .PADOUT(N__35206),
            .PADIN(N__35205),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__35198),
            .DIN(N__35197),
            .DOUT(N__35196),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__35198),
            .PADOUT(N__35197),
            .PADIN(N__35196),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18721),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__35189),
            .DIN(N__35188),
            .DOUT(N__35187),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__35189),
            .PADOUT(N__35188),
            .PADIN(N__35187),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18781),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__35180),
            .DIN(N__35179),
            .DOUT(N__35178),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__35180),
            .PADOUT(N__35179),
            .PADIN(N__35178),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__35171),
            .DIN(N__35170),
            .DOUT(N__35169),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__35171),
            .PADOUT(N__35170),
            .PADIN(N__35169),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__35162),
            .DIN(N__35161),
            .DOUT(N__35160),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__35162),
            .PADOUT(N__35161),
            .PADIN(N__35160),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__35153),
            .DIN(N__35152),
            .DOUT(N__35151),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__35153),
            .PADOUT(N__35152),
            .PADIN(N__35151),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__35144),
            .DIN(N__35143),
            .DOUT(N__35142),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__35144),
            .PADOUT(N__35143),
            .PADIN(N__35142),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34566),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__35135),
            .DIN(N__35134),
            .DOUT(N__35133),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__35135),
            .PADOUT(N__35134),
            .PADIN(N__35133),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__14665),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__35126),
            .DIN(N__35125),
            .DOUT(N__35124),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__35126),
            .PADOUT(N__35125),
            .PADIN(N__35124),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__35117),
            .DIN(N__35116),
            .DOUT(N__35115),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__35117),
            .PADOUT(N__35116),
            .PADIN(N__35115),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29143),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__35108),
            .DIN(N__35107),
            .DOUT(N__35106),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__35108),
            .PADOUT(N__35107),
            .PADIN(N__35106),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__35099),
            .DIN(N__35098),
            .DOUT(N__35097),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__35099),
            .PADOUT(N__35098),
            .PADIN(N__35097),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__35090),
            .DIN(N__35089),
            .DOUT(N__35088),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__35090),
            .PADOUT(N__35089),
            .PADIN(N__35088),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__35081),
            .DIN(N__35080),
            .DOUT(N__35079),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__35081),
            .PADOUT(N__35080),
            .PADIN(N__35079),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__35072),
            .DIN(N__35071),
            .DOUT(N__35070),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__35072),
            .PADOUT(N__35071),
            .PADIN(N__35070),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24859),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__35063),
            .DIN(N__35062),
            .DOUT(N__35061),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__35063),
            .PADOUT(N__35062),
            .PADIN(N__35061),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__35054),
            .DIN(N__35053),
            .DOUT(N__35052),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__35054),
            .PADOUT(N__35053),
            .PADIN(N__35052),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16795),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__35045),
            .DIN(N__35044),
            .DOUT(N__35043),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__35045),
            .PADOUT(N__35044),
            .PADIN(N__35043),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__35036),
            .DIN(N__35035),
            .DOUT(N__35034),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__35036),
            .PADOUT(N__35035),
            .PADIN(N__35034),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31237),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__35027),
            .DIN(N__35026),
            .DOUT(N__35025),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__35027),
            .PADOUT(N__35026),
            .PADIN(N__35025),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24949),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__35018),
            .DIN(N__35017),
            .DOUT(N__35016),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__35018),
            .PADOUT(N__35017),
            .PADIN(N__35016),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__35009),
            .DIN(N__35008),
            .DOUT(N__35007),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__35009),
            .PADOUT(N__35008),
            .PADIN(N__35007),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__35000),
            .DIN(N__34999),
            .DOUT(N__34998),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__35000),
            .PADOUT(N__34999),
            .PADIN(N__34998),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__34991),
            .DIN(N__34990),
            .DOUT(N__34989),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__34991),
            .PADOUT(N__34990),
            .PADIN(N__34989),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__34982),
            .DIN(N__34981),
            .DOUT(N__34980),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__34982),
            .PADOUT(N__34981),
            .PADIN(N__34980),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30916),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__34973),
            .DIN(N__34972),
            .DOUT(N__34971),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__34973),
            .PADOUT(N__34972),
            .PADIN(N__34971),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__34964),
            .DIN(N__34963),
            .DOUT(N__34962),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__34964),
            .PADOUT(N__34963),
            .PADIN(N__34962),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__34955),
            .DIN(N__34954),
            .DOUT(N__34953),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__34955),
            .PADOUT(N__34954),
            .PADIN(N__34953),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__34946),
            .DIN(N__34945),
            .DOUT(N__34944),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__34946),
            .PADOUT(N__34945),
            .PADIN(N__34944),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__34937),
            .DIN(N__34936),
            .DOUT(N__34935),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__34937),
            .PADOUT(N__34936),
            .PADIN(N__34935),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__34928),
            .DIN(N__34927),
            .DOUT(N__34926),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__34928),
            .PADOUT(N__34927),
            .PADIN(N__34926),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__34919),
            .DIN(N__34918),
            .DOUT(N__34917),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__34919),
            .PADOUT(N__34918),
            .PADIN(N__34917),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18771),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__34910),
            .DIN(N__34909),
            .DOUT(N__34908),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__34910),
            .PADOUT(N__34909),
            .PADIN(N__34908),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__8159 (
            .O(N__34891),
            .I(N__34830));
    InMux I__8158 (
            .O(N__34890),
            .I(N__34830));
    InMux I__8157 (
            .O(N__34889),
            .I(N__34830));
    InMux I__8156 (
            .O(N__34888),
            .I(N__34830));
    InMux I__8155 (
            .O(N__34887),
            .I(N__34821));
    InMux I__8154 (
            .O(N__34886),
            .I(N__34821));
    InMux I__8153 (
            .O(N__34885),
            .I(N__34821));
    InMux I__8152 (
            .O(N__34884),
            .I(N__34821));
    InMux I__8151 (
            .O(N__34883),
            .I(N__34812));
    InMux I__8150 (
            .O(N__34882),
            .I(N__34812));
    InMux I__8149 (
            .O(N__34881),
            .I(N__34812));
    InMux I__8148 (
            .O(N__34880),
            .I(N__34812));
    InMux I__8147 (
            .O(N__34879),
            .I(N__34805));
    InMux I__8146 (
            .O(N__34878),
            .I(N__34805));
    InMux I__8145 (
            .O(N__34877),
            .I(N__34805));
    InMux I__8144 (
            .O(N__34876),
            .I(N__34798));
    InMux I__8143 (
            .O(N__34875),
            .I(N__34798));
    InMux I__8142 (
            .O(N__34874),
            .I(N__34798));
    InMux I__8141 (
            .O(N__34873),
            .I(N__34789));
    InMux I__8140 (
            .O(N__34872),
            .I(N__34789));
    InMux I__8139 (
            .O(N__34871),
            .I(N__34789));
    InMux I__8138 (
            .O(N__34870),
            .I(N__34789));
    InMux I__8137 (
            .O(N__34869),
            .I(N__34780));
    InMux I__8136 (
            .O(N__34868),
            .I(N__34780));
    InMux I__8135 (
            .O(N__34867),
            .I(N__34780));
    InMux I__8134 (
            .O(N__34866),
            .I(N__34780));
    InMux I__8133 (
            .O(N__34865),
            .I(N__34771));
    InMux I__8132 (
            .O(N__34864),
            .I(N__34771));
    InMux I__8131 (
            .O(N__34863),
            .I(N__34771));
    InMux I__8130 (
            .O(N__34862),
            .I(N__34771));
    InMux I__8129 (
            .O(N__34861),
            .I(N__34762));
    InMux I__8128 (
            .O(N__34860),
            .I(N__34762));
    InMux I__8127 (
            .O(N__34859),
            .I(N__34762));
    InMux I__8126 (
            .O(N__34858),
            .I(N__34762));
    InMux I__8125 (
            .O(N__34857),
            .I(N__34759));
    InMux I__8124 (
            .O(N__34856),
            .I(N__34754));
    InMux I__8123 (
            .O(N__34855),
            .I(N__34754));
    InMux I__8122 (
            .O(N__34854),
            .I(N__34745));
    InMux I__8121 (
            .O(N__34853),
            .I(N__34745));
    InMux I__8120 (
            .O(N__34852),
            .I(N__34745));
    InMux I__8119 (
            .O(N__34851),
            .I(N__34745));
    InMux I__8118 (
            .O(N__34850),
            .I(N__34736));
    InMux I__8117 (
            .O(N__34849),
            .I(N__34736));
    InMux I__8116 (
            .O(N__34848),
            .I(N__34736));
    InMux I__8115 (
            .O(N__34847),
            .I(N__34736));
    InMux I__8114 (
            .O(N__34846),
            .I(N__34729));
    InMux I__8113 (
            .O(N__34845),
            .I(N__34729));
    InMux I__8112 (
            .O(N__34844),
            .I(N__34729));
    InMux I__8111 (
            .O(N__34843),
            .I(N__34726));
    InMux I__8110 (
            .O(N__34842),
            .I(N__34721));
    InMux I__8109 (
            .O(N__34841),
            .I(N__34721));
    InMux I__8108 (
            .O(N__34840),
            .I(N__34718));
    InMux I__8107 (
            .O(N__34839),
            .I(N__34715));
    LocalMux I__8106 (
            .O(N__34830),
            .I(N__34707));
    LocalMux I__8105 (
            .O(N__34821),
            .I(N__34703));
    LocalMux I__8104 (
            .O(N__34812),
            .I(N__34700));
    LocalMux I__8103 (
            .O(N__34805),
            .I(N__34697));
    LocalMux I__8102 (
            .O(N__34798),
            .I(N__34693));
    LocalMux I__8101 (
            .O(N__34789),
            .I(N__34690));
    LocalMux I__8100 (
            .O(N__34780),
            .I(N__34684));
    LocalMux I__8099 (
            .O(N__34771),
            .I(N__34681));
    LocalMux I__8098 (
            .O(N__34762),
            .I(N__34678));
    LocalMux I__8097 (
            .O(N__34759),
            .I(N__34675));
    LocalMux I__8096 (
            .O(N__34754),
            .I(N__34672));
    LocalMux I__8095 (
            .O(N__34745),
            .I(N__34669));
    LocalMux I__8094 (
            .O(N__34736),
            .I(N__34666));
    LocalMux I__8093 (
            .O(N__34729),
            .I(N__34663));
    LocalMux I__8092 (
            .O(N__34726),
            .I(N__34660));
    LocalMux I__8091 (
            .O(N__34721),
            .I(N__34657));
    LocalMux I__8090 (
            .O(N__34718),
            .I(N__34654));
    LocalMux I__8089 (
            .O(N__34715),
            .I(N__34651));
    CEMux I__8088 (
            .O(N__34714),
            .I(N__34594));
    CEMux I__8087 (
            .O(N__34713),
            .I(N__34594));
    CEMux I__8086 (
            .O(N__34712),
            .I(N__34594));
    CEMux I__8085 (
            .O(N__34711),
            .I(N__34594));
    CEMux I__8084 (
            .O(N__34710),
            .I(N__34594));
    Glb2LocalMux I__8083 (
            .O(N__34707),
            .I(N__34594));
    CEMux I__8082 (
            .O(N__34706),
            .I(N__34594));
    Glb2LocalMux I__8081 (
            .O(N__34703),
            .I(N__34594));
    Glb2LocalMux I__8080 (
            .O(N__34700),
            .I(N__34594));
    Glb2LocalMux I__8079 (
            .O(N__34697),
            .I(N__34594));
    CEMux I__8078 (
            .O(N__34696),
            .I(N__34594));
    Glb2LocalMux I__8077 (
            .O(N__34693),
            .I(N__34594));
    Glb2LocalMux I__8076 (
            .O(N__34690),
            .I(N__34594));
    CEMux I__8075 (
            .O(N__34689),
            .I(N__34594));
    CEMux I__8074 (
            .O(N__34688),
            .I(N__34594));
    CEMux I__8073 (
            .O(N__34687),
            .I(N__34594));
    Glb2LocalMux I__8072 (
            .O(N__34684),
            .I(N__34594));
    Glb2LocalMux I__8071 (
            .O(N__34681),
            .I(N__34594));
    Glb2LocalMux I__8070 (
            .O(N__34678),
            .I(N__34594));
    Glb2LocalMux I__8069 (
            .O(N__34675),
            .I(N__34594));
    Glb2LocalMux I__8068 (
            .O(N__34672),
            .I(N__34594));
    Glb2LocalMux I__8067 (
            .O(N__34669),
            .I(N__34594));
    Glb2LocalMux I__8066 (
            .O(N__34666),
            .I(N__34594));
    Glb2LocalMux I__8065 (
            .O(N__34663),
            .I(N__34594));
    Glb2LocalMux I__8064 (
            .O(N__34660),
            .I(N__34594));
    Glb2LocalMux I__8063 (
            .O(N__34657),
            .I(N__34594));
    Glb2LocalMux I__8062 (
            .O(N__34654),
            .I(N__34594));
    Glb2LocalMux I__8061 (
            .O(N__34651),
            .I(N__34594));
    GlobalMux I__8060 (
            .O(N__34594),
            .I(N__34591));
    gio2CtrlBuf I__8059 (
            .O(N__34591),
            .I(N_29_g));
    InMux I__8058 (
            .O(N__34588),
            .I(N__34584));
    InMux I__8057 (
            .O(N__34587),
            .I(N__34581));
    LocalMux I__8056 (
            .O(N__34584),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__8055 (
            .O(N__34581),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__8054 (
            .O(N__34576),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    InMux I__8053 (
            .O(N__34573),
            .I(N__34570));
    LocalMux I__8052 (
            .O(N__34570),
            .I(N__34567));
    Span4Mux_s3_v I__8051 (
            .O(N__34567),
            .I(N__34562));
    IoInMux I__8050 (
            .O(N__34566),
            .I(N__34558));
    InMux I__8049 (
            .O(N__34565),
            .I(N__34553));
    Span4Mux_h I__8048 (
            .O(N__34562),
            .I(N__34550));
    InMux I__8047 (
            .O(N__34561),
            .I(N__34547));
    LocalMux I__8046 (
            .O(N__34558),
            .I(N__34544));
    InMux I__8045 (
            .O(N__34557),
            .I(N__34541));
    InMux I__8044 (
            .O(N__34556),
            .I(N__34538));
    LocalMux I__8043 (
            .O(N__34553),
            .I(N__34534));
    Span4Mux_h I__8042 (
            .O(N__34550),
            .I(N__34529));
    LocalMux I__8041 (
            .O(N__34547),
            .I(N__34529));
    Span4Mux_s3_h I__8040 (
            .O(N__34544),
            .I(N__34526));
    LocalMux I__8039 (
            .O(N__34541),
            .I(N__34523));
    LocalMux I__8038 (
            .O(N__34538),
            .I(N__34520));
    InMux I__8037 (
            .O(N__34537),
            .I(N__34517));
    Span4Mux_v I__8036 (
            .O(N__34534),
            .I(N__34514));
    Span4Mux_v I__8035 (
            .O(N__34529),
            .I(N__34511));
    Span4Mux_v I__8034 (
            .O(N__34526),
            .I(N__34506));
    Span4Mux_v I__8033 (
            .O(N__34523),
            .I(N__34506));
    Span4Mux_v I__8032 (
            .O(N__34520),
            .I(N__34501));
    LocalMux I__8031 (
            .O(N__34517),
            .I(N__34501));
    Span4Mux_h I__8030 (
            .O(N__34514),
            .I(N__34497));
    Span4Mux_v I__8029 (
            .O(N__34511),
            .I(N__34494));
    Span4Mux_h I__8028 (
            .O(N__34506),
            .I(N__34489));
    Span4Mux_v I__8027 (
            .O(N__34501),
            .I(N__34489));
    InMux I__8026 (
            .O(N__34500),
            .I(N__34486));
    Odrv4 I__8025 (
            .O(N__34497),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8024 (
            .O(N__34494),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__8023 (
            .O(N__34489),
            .I(CONSTANT_ONE_NET));
    LocalMux I__8022 (
            .O(N__34486),
            .I(CONSTANT_ONE_NET));
    InMux I__8021 (
            .O(N__34477),
            .I(bfn_12_16_0_));
    InMux I__8020 (
            .O(N__34474),
            .I(N__34470));
    InMux I__8019 (
            .O(N__34473),
            .I(N__34467));
    LocalMux I__8018 (
            .O(N__34470),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    LocalMux I__8017 (
            .O(N__34467),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    ClkMux I__8016 (
            .O(N__34462),
            .I(N__34455));
    ClkMux I__8015 (
            .O(N__34461),
            .I(N__34452));
    ClkMux I__8014 (
            .O(N__34460),
            .I(N__34446));
    ClkMux I__8013 (
            .O(N__34459),
            .I(N__34441));
    ClkMux I__8012 (
            .O(N__34458),
            .I(N__34435));
    LocalMux I__8011 (
            .O(N__34455),
            .I(N__34426));
    LocalMux I__8010 (
            .O(N__34452),
            .I(N__34422));
    ClkMux I__8009 (
            .O(N__34451),
            .I(N__34418));
    ClkMux I__8008 (
            .O(N__34450),
            .I(N__34413));
    ClkMux I__8007 (
            .O(N__34449),
            .I(N__34409));
    LocalMux I__8006 (
            .O(N__34446),
            .I(N__34406));
    ClkMux I__8005 (
            .O(N__34445),
            .I(N__34403));
    ClkMux I__8004 (
            .O(N__34444),
            .I(N__34400));
    LocalMux I__8003 (
            .O(N__34441),
            .I(N__34397));
    ClkMux I__8002 (
            .O(N__34440),
            .I(N__34394));
    ClkMux I__8001 (
            .O(N__34439),
            .I(N__34391));
    ClkMux I__8000 (
            .O(N__34438),
            .I(N__34385));
    LocalMux I__7999 (
            .O(N__34435),
            .I(N__34382));
    ClkMux I__7998 (
            .O(N__34434),
            .I(N__34379));
    ClkMux I__7997 (
            .O(N__34433),
            .I(N__34375));
    ClkMux I__7996 (
            .O(N__34432),
            .I(N__34369));
    ClkMux I__7995 (
            .O(N__34431),
            .I(N__34365));
    ClkMux I__7994 (
            .O(N__34430),
            .I(N__34362));
    ClkMux I__7993 (
            .O(N__34429),
            .I(N__34358));
    Span4Mux_s1_h I__7992 (
            .O(N__34426),
            .I(N__34354));
    ClkMux I__7991 (
            .O(N__34425),
            .I(N__34351));
    Span4Mux_s1_h I__7990 (
            .O(N__34422),
            .I(N__34345));
    ClkMux I__7989 (
            .O(N__34421),
            .I(N__34342));
    LocalMux I__7988 (
            .O(N__34418),
            .I(N__34339));
    ClkMux I__7987 (
            .O(N__34417),
            .I(N__34336));
    ClkMux I__7986 (
            .O(N__34416),
            .I(N__34333));
    LocalMux I__7985 (
            .O(N__34413),
            .I(N__34329));
    ClkMux I__7984 (
            .O(N__34412),
            .I(N__34325));
    LocalMux I__7983 (
            .O(N__34409),
            .I(N__34318));
    Span4Mux_v I__7982 (
            .O(N__34406),
            .I(N__34311));
    LocalMux I__7981 (
            .O(N__34403),
            .I(N__34311));
    LocalMux I__7980 (
            .O(N__34400),
            .I(N__34311));
    Span4Mux_v I__7979 (
            .O(N__34397),
            .I(N__34304));
    LocalMux I__7978 (
            .O(N__34394),
            .I(N__34304));
    LocalMux I__7977 (
            .O(N__34391),
            .I(N__34304));
    ClkMux I__7976 (
            .O(N__34390),
            .I(N__34301));
    ClkMux I__7975 (
            .O(N__34389),
            .I(N__34298));
    ClkMux I__7974 (
            .O(N__34388),
            .I(N__34295));
    LocalMux I__7973 (
            .O(N__34385),
            .I(N__34285));
    Span4Mux_h I__7972 (
            .O(N__34382),
            .I(N__34285));
    LocalMux I__7971 (
            .O(N__34379),
            .I(N__34285));
    ClkMux I__7970 (
            .O(N__34378),
            .I(N__34282));
    LocalMux I__7969 (
            .O(N__34375),
            .I(N__34279));
    ClkMux I__7968 (
            .O(N__34374),
            .I(N__34276));
    ClkMux I__7967 (
            .O(N__34373),
            .I(N__34272));
    ClkMux I__7966 (
            .O(N__34372),
            .I(N__34268));
    LocalMux I__7965 (
            .O(N__34369),
            .I(N__34264));
    ClkMux I__7964 (
            .O(N__34368),
            .I(N__34261));
    LocalMux I__7963 (
            .O(N__34365),
            .I(N__34258));
    LocalMux I__7962 (
            .O(N__34362),
            .I(N__34255));
    ClkMux I__7961 (
            .O(N__34361),
            .I(N__34252));
    LocalMux I__7960 (
            .O(N__34358),
            .I(N__34249));
    ClkMux I__7959 (
            .O(N__34357),
            .I(N__34246));
    Span4Mux_v I__7958 (
            .O(N__34354),
            .I(N__34241));
    LocalMux I__7957 (
            .O(N__34351),
            .I(N__34241));
    ClkMux I__7956 (
            .O(N__34350),
            .I(N__34237));
    ClkMux I__7955 (
            .O(N__34349),
            .I(N__34234));
    ClkMux I__7954 (
            .O(N__34348),
            .I(N__34230));
    Span4Mux_v I__7953 (
            .O(N__34345),
            .I(N__34225));
    LocalMux I__7952 (
            .O(N__34342),
            .I(N__34225));
    Span4Mux_s2_h I__7951 (
            .O(N__34339),
            .I(N__34217));
    LocalMux I__7950 (
            .O(N__34336),
            .I(N__34217));
    LocalMux I__7949 (
            .O(N__34333),
            .I(N__34214));
    ClkMux I__7948 (
            .O(N__34332),
            .I(N__34211));
    Span4Mux_s2_h I__7947 (
            .O(N__34329),
            .I(N__34207));
    ClkMux I__7946 (
            .O(N__34328),
            .I(N__34204));
    LocalMux I__7945 (
            .O(N__34325),
            .I(N__34201));
    ClkMux I__7944 (
            .O(N__34324),
            .I(N__34198));
    ClkMux I__7943 (
            .O(N__34323),
            .I(N__34192));
    ClkMux I__7942 (
            .O(N__34322),
            .I(N__34189));
    ClkMux I__7941 (
            .O(N__34321),
            .I(N__34186));
    Span4Mux_h I__7940 (
            .O(N__34318),
            .I(N__34182));
    Span4Mux_v I__7939 (
            .O(N__34311),
            .I(N__34171));
    Span4Mux_v I__7938 (
            .O(N__34304),
            .I(N__34171));
    LocalMux I__7937 (
            .O(N__34301),
            .I(N__34171));
    LocalMux I__7936 (
            .O(N__34298),
            .I(N__34171));
    LocalMux I__7935 (
            .O(N__34295),
            .I(N__34171));
    ClkMux I__7934 (
            .O(N__34294),
            .I(N__34167));
    ClkMux I__7933 (
            .O(N__34293),
            .I(N__34164));
    ClkMux I__7932 (
            .O(N__34292),
            .I(N__34158));
    Span4Mux_v I__7931 (
            .O(N__34285),
            .I(N__34153));
    LocalMux I__7930 (
            .O(N__34282),
            .I(N__34153));
    Span4Mux_s1_h I__7929 (
            .O(N__34279),
            .I(N__34148));
    LocalMux I__7928 (
            .O(N__34276),
            .I(N__34148));
    ClkMux I__7927 (
            .O(N__34275),
            .I(N__34145));
    LocalMux I__7926 (
            .O(N__34272),
            .I(N__34140));
    ClkMux I__7925 (
            .O(N__34271),
            .I(N__34137));
    LocalMux I__7924 (
            .O(N__34268),
            .I(N__34134));
    ClkMux I__7923 (
            .O(N__34267),
            .I(N__34131));
    Span4Mux_h I__7922 (
            .O(N__34264),
            .I(N__34126));
    LocalMux I__7921 (
            .O(N__34261),
            .I(N__34126));
    Span4Mux_v I__7920 (
            .O(N__34258),
            .I(N__34119));
    Span4Mux_s1_h I__7919 (
            .O(N__34255),
            .I(N__34119));
    LocalMux I__7918 (
            .O(N__34252),
            .I(N__34119));
    Span4Mux_s2_h I__7917 (
            .O(N__34249),
            .I(N__34114));
    LocalMux I__7916 (
            .O(N__34246),
            .I(N__34114));
    Span4Mux_h I__7915 (
            .O(N__34241),
            .I(N__34111));
    ClkMux I__7914 (
            .O(N__34240),
            .I(N__34108));
    LocalMux I__7913 (
            .O(N__34237),
            .I(N__34105));
    LocalMux I__7912 (
            .O(N__34234),
            .I(N__34102));
    ClkMux I__7911 (
            .O(N__34233),
            .I(N__34099));
    LocalMux I__7910 (
            .O(N__34230),
            .I(N__34096));
    Span4Mux_s1_h I__7909 (
            .O(N__34225),
            .I(N__34093));
    ClkMux I__7908 (
            .O(N__34224),
            .I(N__34090));
    ClkMux I__7907 (
            .O(N__34223),
            .I(N__34087));
    ClkMux I__7906 (
            .O(N__34222),
            .I(N__34081));
    Span4Mux_v I__7905 (
            .O(N__34217),
            .I(N__34073));
    Span4Mux_s2_h I__7904 (
            .O(N__34214),
            .I(N__34073));
    LocalMux I__7903 (
            .O(N__34211),
            .I(N__34073));
    ClkMux I__7902 (
            .O(N__34210),
            .I(N__34070));
    Span4Mux_v I__7901 (
            .O(N__34207),
            .I(N__34064));
    LocalMux I__7900 (
            .O(N__34204),
            .I(N__34064));
    Span4Mux_s2_h I__7899 (
            .O(N__34201),
            .I(N__34059));
    LocalMux I__7898 (
            .O(N__34198),
            .I(N__34059));
    ClkMux I__7897 (
            .O(N__34197),
            .I(N__34056));
    ClkMux I__7896 (
            .O(N__34196),
            .I(N__34052));
    ClkMux I__7895 (
            .O(N__34195),
            .I(N__34049));
    LocalMux I__7894 (
            .O(N__34192),
            .I(N__34046));
    LocalMux I__7893 (
            .O(N__34189),
            .I(N__34041));
    LocalMux I__7892 (
            .O(N__34186),
            .I(N__34041));
    ClkMux I__7891 (
            .O(N__34185),
            .I(N__34038));
    Span4Mux_v I__7890 (
            .O(N__34182),
            .I(N__34035));
    Span4Mux_v I__7889 (
            .O(N__34171),
            .I(N__34032));
    ClkMux I__7888 (
            .O(N__34170),
            .I(N__34029));
    LocalMux I__7887 (
            .O(N__34167),
            .I(N__34024));
    LocalMux I__7886 (
            .O(N__34164),
            .I(N__34024));
    ClkMux I__7885 (
            .O(N__34163),
            .I(N__34021));
    ClkMux I__7884 (
            .O(N__34162),
            .I(N__34017));
    ClkMux I__7883 (
            .O(N__34161),
            .I(N__34014));
    LocalMux I__7882 (
            .O(N__34158),
            .I(N__34010));
    Span4Mux_v I__7881 (
            .O(N__34153),
            .I(N__34003));
    Span4Mux_v I__7880 (
            .O(N__34148),
            .I(N__34003));
    LocalMux I__7879 (
            .O(N__34145),
            .I(N__34003));
    ClkMux I__7878 (
            .O(N__34144),
            .I(N__34000));
    ClkMux I__7877 (
            .O(N__34143),
            .I(N__33993));
    Span4Mux_s3_h I__7876 (
            .O(N__34140),
            .I(N__33984));
    LocalMux I__7875 (
            .O(N__34137),
            .I(N__33984));
    Span4Mux_s3_h I__7874 (
            .O(N__34134),
            .I(N__33984));
    LocalMux I__7873 (
            .O(N__34131),
            .I(N__33984));
    Span4Mux_v I__7872 (
            .O(N__34126),
            .I(N__33980));
    Span4Mux_h I__7871 (
            .O(N__34119),
            .I(N__33975));
    Span4Mux_h I__7870 (
            .O(N__34114),
            .I(N__33975));
    Span4Mux_h I__7869 (
            .O(N__34111),
            .I(N__33970));
    LocalMux I__7868 (
            .O(N__34108),
            .I(N__33970));
    Span4Mux_s1_h I__7867 (
            .O(N__34105),
            .I(N__33963));
    Span4Mux_h I__7866 (
            .O(N__34102),
            .I(N__33963));
    LocalMux I__7865 (
            .O(N__34099),
            .I(N__33963));
    Span4Mux_s1_h I__7864 (
            .O(N__34096),
            .I(N__33960));
    Span4Mux_h I__7863 (
            .O(N__34093),
            .I(N__33955));
    LocalMux I__7862 (
            .O(N__34090),
            .I(N__33955));
    LocalMux I__7861 (
            .O(N__34087),
            .I(N__33952));
    ClkMux I__7860 (
            .O(N__34086),
            .I(N__33949));
    ClkMux I__7859 (
            .O(N__34085),
            .I(N__33946));
    ClkMux I__7858 (
            .O(N__34084),
            .I(N__33943));
    LocalMux I__7857 (
            .O(N__34081),
            .I(N__33940));
    ClkMux I__7856 (
            .O(N__34080),
            .I(N__33937));
    Span4Mux_v I__7855 (
            .O(N__34073),
            .I(N__33932));
    LocalMux I__7854 (
            .O(N__34070),
            .I(N__33932));
    ClkMux I__7853 (
            .O(N__34069),
            .I(N__33929));
    Span4Mux_v I__7852 (
            .O(N__34064),
            .I(N__33922));
    Span4Mux_h I__7851 (
            .O(N__34059),
            .I(N__33922));
    LocalMux I__7850 (
            .O(N__34056),
            .I(N__33922));
    ClkMux I__7849 (
            .O(N__34055),
            .I(N__33919));
    LocalMux I__7848 (
            .O(N__34052),
            .I(N__33916));
    LocalMux I__7847 (
            .O(N__34049),
            .I(N__33913));
    Span4Mux_v I__7846 (
            .O(N__34046),
            .I(N__33906));
    Span4Mux_h I__7845 (
            .O(N__34041),
            .I(N__33906));
    LocalMux I__7844 (
            .O(N__34038),
            .I(N__33906));
    Span4Mux_h I__7843 (
            .O(N__34035),
            .I(N__33895));
    Span4Mux_h I__7842 (
            .O(N__34032),
            .I(N__33895));
    LocalMux I__7841 (
            .O(N__34029),
            .I(N__33895));
    Span4Mux_h I__7840 (
            .O(N__34024),
            .I(N__33895));
    LocalMux I__7839 (
            .O(N__34021),
            .I(N__33895));
    ClkMux I__7838 (
            .O(N__34020),
            .I(N__33892));
    LocalMux I__7837 (
            .O(N__34017),
            .I(N__33889));
    LocalMux I__7836 (
            .O(N__34014),
            .I(N__33886));
    ClkMux I__7835 (
            .O(N__34013),
            .I(N__33883));
    Span4Mux_s1_h I__7834 (
            .O(N__34010),
            .I(N__33876));
    Span4Mux_s2_v I__7833 (
            .O(N__34003),
            .I(N__33876));
    LocalMux I__7832 (
            .O(N__34000),
            .I(N__33876));
    ClkMux I__7831 (
            .O(N__33999),
            .I(N__33872));
    ClkMux I__7830 (
            .O(N__33998),
            .I(N__33869));
    ClkMux I__7829 (
            .O(N__33997),
            .I(N__33866));
    ClkMux I__7828 (
            .O(N__33996),
            .I(N__33863));
    LocalMux I__7827 (
            .O(N__33993),
            .I(N__33860));
    Span4Mux_v I__7826 (
            .O(N__33984),
            .I(N__33857));
    ClkMux I__7825 (
            .O(N__33983),
            .I(N__33854));
    Span4Mux_v I__7824 (
            .O(N__33980),
            .I(N__33850));
    Span4Mux_v I__7823 (
            .O(N__33975),
            .I(N__33843));
    Span4Mux_v I__7822 (
            .O(N__33970),
            .I(N__33843));
    Span4Mux_h I__7821 (
            .O(N__33963),
            .I(N__33843));
    Span4Mux_h I__7820 (
            .O(N__33960),
            .I(N__33830));
    Span4Mux_v I__7819 (
            .O(N__33955),
            .I(N__33830));
    Span4Mux_h I__7818 (
            .O(N__33952),
            .I(N__33830));
    LocalMux I__7817 (
            .O(N__33949),
            .I(N__33830));
    LocalMux I__7816 (
            .O(N__33946),
            .I(N__33830));
    LocalMux I__7815 (
            .O(N__33943),
            .I(N__33830));
    Span4Mux_s1_h I__7814 (
            .O(N__33940),
            .I(N__33825));
    LocalMux I__7813 (
            .O(N__33937),
            .I(N__33825));
    Span4Mux_v I__7812 (
            .O(N__33932),
            .I(N__33820));
    LocalMux I__7811 (
            .O(N__33929),
            .I(N__33820));
    Span4Mux_v I__7810 (
            .O(N__33922),
            .I(N__33815));
    LocalMux I__7809 (
            .O(N__33919),
            .I(N__33815));
    Span4Mux_v I__7808 (
            .O(N__33916),
            .I(N__33804));
    Span4Mux_h I__7807 (
            .O(N__33913),
            .I(N__33804));
    IoSpan4Mux I__7806 (
            .O(N__33906),
            .I(N__33804));
    Span4Mux_v I__7805 (
            .O(N__33895),
            .I(N__33804));
    LocalMux I__7804 (
            .O(N__33892),
            .I(N__33804));
    Span4Mux_v I__7803 (
            .O(N__33889),
            .I(N__33795));
    Span4Mux_h I__7802 (
            .O(N__33886),
            .I(N__33795));
    LocalMux I__7801 (
            .O(N__33883),
            .I(N__33795));
    Span4Mux_h I__7800 (
            .O(N__33876),
            .I(N__33795));
    ClkMux I__7799 (
            .O(N__33875),
            .I(N__33792));
    LocalMux I__7798 (
            .O(N__33872),
            .I(N__33789));
    LocalMux I__7797 (
            .O(N__33869),
            .I(N__33786));
    LocalMux I__7796 (
            .O(N__33866),
            .I(N__33781));
    LocalMux I__7795 (
            .O(N__33863),
            .I(N__33781));
    Span12Mux_s5_h I__7794 (
            .O(N__33860),
            .I(N__33778));
    Sp12to4 I__7793 (
            .O(N__33857),
            .I(N__33775));
    LocalMux I__7792 (
            .O(N__33854),
            .I(N__33772));
    ClkMux I__7791 (
            .O(N__33853),
            .I(N__33769));
    IoSpan4Mux I__7790 (
            .O(N__33850),
            .I(N__33766));
    Span4Mux_v I__7789 (
            .O(N__33843),
            .I(N__33763));
    Span4Mux_v I__7788 (
            .O(N__33830),
            .I(N__33758));
    Span4Mux_h I__7787 (
            .O(N__33825),
            .I(N__33758));
    IoSpan4Mux I__7786 (
            .O(N__33820),
            .I(N__33751));
    IoSpan4Mux I__7785 (
            .O(N__33815),
            .I(N__33751));
    IoSpan4Mux I__7784 (
            .O(N__33804),
            .I(N__33751));
    Span4Mux_v I__7783 (
            .O(N__33795),
            .I(N__33746));
    LocalMux I__7782 (
            .O(N__33792),
            .I(N__33746));
    Span12Mux_s5_h I__7781 (
            .O(N__33789),
            .I(N__33739));
    Sp12to4 I__7780 (
            .O(N__33786),
            .I(N__33739));
    Sp12to4 I__7779 (
            .O(N__33781),
            .I(N__33739));
    Span12Mux_v I__7778 (
            .O(N__33778),
            .I(N__33730));
    Span12Mux_s6_h I__7777 (
            .O(N__33775),
            .I(N__33730));
    Span12Mux_s5_h I__7776 (
            .O(N__33772),
            .I(N__33730));
    LocalMux I__7775 (
            .O(N__33769),
            .I(N__33730));
    Odrv4 I__7774 (
            .O(N__33766),
            .I(fpga_osc));
    Odrv4 I__7773 (
            .O(N__33763),
            .I(fpga_osc));
    Odrv4 I__7772 (
            .O(N__33758),
            .I(fpga_osc));
    Odrv4 I__7771 (
            .O(N__33751),
            .I(fpga_osc));
    Odrv4 I__7770 (
            .O(N__33746),
            .I(fpga_osc));
    Odrv12 I__7769 (
            .O(N__33739),
            .I(fpga_osc));
    Odrv12 I__7768 (
            .O(N__33730),
            .I(fpga_osc));
    CEMux I__7767 (
            .O(N__33715),
            .I(N__33712));
    LocalMux I__7766 (
            .O(N__33712),
            .I(\VPP_VDDQ.N_29_0 ));
    SRMux I__7765 (
            .O(N__33709),
            .I(N__33706));
    LocalMux I__7764 (
            .O(N__33706),
            .I(N__33700));
    SRMux I__7763 (
            .O(N__33705),
            .I(N__33697));
    SRMux I__7762 (
            .O(N__33704),
            .I(N__33694));
    InMux I__7761 (
            .O(N__33703),
            .I(N__33691));
    Span4Mux_s1_h I__7760 (
            .O(N__33700),
            .I(N__33688));
    LocalMux I__7759 (
            .O(N__33697),
            .I(N__33683));
    LocalMux I__7758 (
            .O(N__33694),
            .I(N__33683));
    LocalMux I__7757 (
            .O(N__33691),
            .I(N__33680));
    Odrv4 I__7756 (
            .O(N__33688),
            .I(G_43));
    Odrv4 I__7755 (
            .O(N__33683),
            .I(G_43));
    Odrv4 I__7754 (
            .O(N__33680),
            .I(G_43));
    InMux I__7753 (
            .O(N__33673),
            .I(N__33669));
    InMux I__7752 (
            .O(N__33672),
            .I(N__33666));
    LocalMux I__7751 (
            .O(N__33669),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__7750 (
            .O(N__33666),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__7749 (
            .O(N__33661),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    InMux I__7748 (
            .O(N__33658),
            .I(N__33654));
    InMux I__7747 (
            .O(N__33657),
            .I(N__33651));
    LocalMux I__7746 (
            .O(N__33654),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__7745 (
            .O(N__33651),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__7744 (
            .O(N__33646),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__7743 (
            .O(N__33643),
            .I(N__33639));
    InMux I__7742 (
            .O(N__33642),
            .I(N__33636));
    LocalMux I__7741 (
            .O(N__33639),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    LocalMux I__7740 (
            .O(N__33636),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__7739 (
            .O(N__33631),
            .I(bfn_12_15_0_));
    InMux I__7738 (
            .O(N__33628),
            .I(N__33624));
    InMux I__7737 (
            .O(N__33627),
            .I(N__33621));
    LocalMux I__7736 (
            .O(N__33624),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__7735 (
            .O(N__33621),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__7734 (
            .O(N__33616),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    CascadeMux I__7733 (
            .O(N__33613),
            .I(N__33609));
    InMux I__7732 (
            .O(N__33612),
            .I(N__33606));
    InMux I__7731 (
            .O(N__33609),
            .I(N__33603));
    LocalMux I__7730 (
            .O(N__33606),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__7729 (
            .O(N__33603),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__7728 (
            .O(N__33598),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    InMux I__7727 (
            .O(N__33595),
            .I(N__33591));
    InMux I__7726 (
            .O(N__33594),
            .I(N__33588));
    LocalMux I__7725 (
            .O(N__33591),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__7724 (
            .O(N__33588),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__7723 (
            .O(N__33583),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    InMux I__7722 (
            .O(N__33580),
            .I(N__33576));
    InMux I__7721 (
            .O(N__33579),
            .I(N__33573));
    LocalMux I__7720 (
            .O(N__33576),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    LocalMux I__7719 (
            .O(N__33573),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__7718 (
            .O(N__33568),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    CascadeMux I__7717 (
            .O(N__33565),
            .I(N__33561));
    InMux I__7716 (
            .O(N__33564),
            .I(N__33558));
    InMux I__7715 (
            .O(N__33561),
            .I(N__33555));
    LocalMux I__7714 (
            .O(N__33558),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__7713 (
            .O(N__33555),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__7712 (
            .O(N__33550),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__7711 (
            .O(N__33547),
            .I(N__33544));
    LocalMux I__7710 (
            .O(N__33544),
            .I(N__33540));
    CascadeMux I__7709 (
            .O(N__33543),
            .I(N__33536));
    Span4Mux_s1_h I__7708 (
            .O(N__33540),
            .I(N__33533));
    InMux I__7707 (
            .O(N__33539),
            .I(N__33530));
    InMux I__7706 (
            .O(N__33536),
            .I(N__33527));
    Odrv4 I__7705 (
            .O(N__33533),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__7704 (
            .O(N__33530),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__7703 (
            .O(N__33527),
            .I(\POWERLED.count_clkZ0Z_4 ));
    InMux I__7702 (
            .O(N__33520),
            .I(N__33517));
    LocalMux I__7701 (
            .O(N__33517),
            .I(\POWERLED.count_clk_RNIZ0Z_12 ));
    CascadeMux I__7700 (
            .O(N__33514),
            .I(\POWERLED.count_clkZ0Z_2_cascade_ ));
    InMux I__7699 (
            .O(N__33511),
            .I(N__33508));
    LocalMux I__7698 (
            .O(N__33508),
            .I(N__33504));
    InMux I__7697 (
            .O(N__33507),
            .I(N__33501));
    Odrv4 I__7696 (
            .O(N__33504),
            .I(\POWERLED.count_clk_RNIZ0Z_15 ));
    LocalMux I__7695 (
            .O(N__33501),
            .I(\POWERLED.count_clk_RNIZ0Z_15 ));
    InMux I__7694 (
            .O(N__33496),
            .I(N__33493));
    LocalMux I__7693 (
            .O(N__33493),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1 ));
    CascadeMux I__7692 (
            .O(N__33490),
            .I(N__33480));
    CascadeMux I__7691 (
            .O(N__33489),
            .I(N__33477));
    CascadeMux I__7690 (
            .O(N__33488),
            .I(N__33472));
    InMux I__7689 (
            .O(N__33487),
            .I(N__33466));
    InMux I__7688 (
            .O(N__33486),
            .I(N__33461));
    InMux I__7687 (
            .O(N__33485),
            .I(N__33461));
    InMux I__7686 (
            .O(N__33484),
            .I(N__33444));
    InMux I__7685 (
            .O(N__33483),
            .I(N__33444));
    InMux I__7684 (
            .O(N__33480),
            .I(N__33444));
    InMux I__7683 (
            .O(N__33477),
            .I(N__33444));
    InMux I__7682 (
            .O(N__33476),
            .I(N__33437));
    InMux I__7681 (
            .O(N__33475),
            .I(N__33437));
    InMux I__7680 (
            .O(N__33472),
            .I(N__33437));
    InMux I__7679 (
            .O(N__33471),
            .I(N__33434));
    InMux I__7678 (
            .O(N__33470),
            .I(N__33429));
    InMux I__7677 (
            .O(N__33469),
            .I(N__33429));
    LocalMux I__7676 (
            .O(N__33466),
            .I(N__33424));
    LocalMux I__7675 (
            .O(N__33461),
            .I(N__33424));
    InMux I__7674 (
            .O(N__33460),
            .I(N__33419));
    InMux I__7673 (
            .O(N__33459),
            .I(N__33419));
    CascadeMux I__7672 (
            .O(N__33458),
            .I(N__33413));
    InMux I__7671 (
            .O(N__33457),
            .I(N__33408));
    InMux I__7670 (
            .O(N__33456),
            .I(N__33403));
    InMux I__7669 (
            .O(N__33455),
            .I(N__33403));
    InMux I__7668 (
            .O(N__33454),
            .I(N__33400));
    InMux I__7667 (
            .O(N__33453),
            .I(N__33397));
    LocalMux I__7666 (
            .O(N__33444),
            .I(N__33392));
    LocalMux I__7665 (
            .O(N__33437),
            .I(N__33392));
    LocalMux I__7664 (
            .O(N__33434),
            .I(N__33383));
    LocalMux I__7663 (
            .O(N__33429),
            .I(N__33383));
    Span4Mux_v I__7662 (
            .O(N__33424),
            .I(N__33383));
    LocalMux I__7661 (
            .O(N__33419),
            .I(N__33383));
    InMux I__7660 (
            .O(N__33418),
            .I(N__33370));
    InMux I__7659 (
            .O(N__33417),
            .I(N__33370));
    InMux I__7658 (
            .O(N__33416),
            .I(N__33370));
    InMux I__7657 (
            .O(N__33413),
            .I(N__33370));
    InMux I__7656 (
            .O(N__33412),
            .I(N__33370));
    InMux I__7655 (
            .O(N__33411),
            .I(N__33370));
    LocalMux I__7654 (
            .O(N__33408),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    LocalMux I__7653 (
            .O(N__33403),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    LocalMux I__7652 (
            .O(N__33400),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    LocalMux I__7651 (
            .O(N__33397),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    Odrv12 I__7650 (
            .O(N__33392),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    Odrv4 I__7649 (
            .O(N__33383),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    LocalMux I__7648 (
            .O(N__33370),
            .I(\POWERLED.func_state_RNIH9594_0_1 ));
    InMux I__7647 (
            .O(N__33355),
            .I(N__33349));
    InMux I__7646 (
            .O(N__33354),
            .I(N__33349));
    LocalMux I__7645 (
            .O(N__33349),
            .I(N__33346));
    Odrv4 I__7644 (
            .O(N__33346),
            .I(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ));
    CascadeMux I__7643 (
            .O(N__33343),
            .I(N__33340));
    InMux I__7642 (
            .O(N__33340),
            .I(N__33337));
    LocalMux I__7641 (
            .O(N__33337),
            .I(\POWERLED.count_clk_0_11 ));
    CEMux I__7640 (
            .O(N__33334),
            .I(N__33328));
    CEMux I__7639 (
            .O(N__33333),
            .I(N__33325));
    CEMux I__7638 (
            .O(N__33332),
            .I(N__33321));
    CEMux I__7637 (
            .O(N__33331),
            .I(N__33313));
    LocalMux I__7636 (
            .O(N__33328),
            .I(N__33310));
    LocalMux I__7635 (
            .O(N__33325),
            .I(N__33307));
    CEMux I__7634 (
            .O(N__33324),
            .I(N__33304));
    LocalMux I__7633 (
            .O(N__33321),
            .I(N__33301));
    CascadeMux I__7632 (
            .O(N__33320),
            .I(N__33298));
    InMux I__7631 (
            .O(N__33319),
            .I(N__33293));
    InMux I__7630 (
            .O(N__33318),
            .I(N__33293));
    CEMux I__7629 (
            .O(N__33317),
            .I(N__33282));
    CEMux I__7628 (
            .O(N__33316),
            .I(N__33279));
    LocalMux I__7627 (
            .O(N__33313),
            .I(N__33276));
    Span4Mux_v I__7626 (
            .O(N__33310),
            .I(N__33271));
    Span4Mux_s0_h I__7625 (
            .O(N__33307),
            .I(N__33271));
    LocalMux I__7624 (
            .O(N__33304),
            .I(N__33268));
    Span4Mux_v I__7623 (
            .O(N__33301),
            .I(N__33264));
    InMux I__7622 (
            .O(N__33298),
            .I(N__33261));
    LocalMux I__7621 (
            .O(N__33293),
            .I(N__33258));
    CascadeMux I__7620 (
            .O(N__33292),
            .I(N__33254));
    InMux I__7619 (
            .O(N__33291),
            .I(N__33247));
    InMux I__7618 (
            .O(N__33290),
            .I(N__33247));
    InMux I__7617 (
            .O(N__33289),
            .I(N__33247));
    InMux I__7616 (
            .O(N__33288),
            .I(N__33238));
    InMux I__7615 (
            .O(N__33287),
            .I(N__33238));
    InMux I__7614 (
            .O(N__33286),
            .I(N__33238));
    InMux I__7613 (
            .O(N__33285),
            .I(N__33238));
    LocalMux I__7612 (
            .O(N__33282),
            .I(N__33232));
    LocalMux I__7611 (
            .O(N__33279),
            .I(N__33229));
    Span4Mux_v I__7610 (
            .O(N__33276),
            .I(N__33224));
    Span4Mux_h I__7609 (
            .O(N__33271),
            .I(N__33224));
    Sp12to4 I__7608 (
            .O(N__33268),
            .I(N__33221));
    InMux I__7607 (
            .O(N__33267),
            .I(N__33218));
    Span4Mux_h I__7606 (
            .O(N__33264),
            .I(N__33211));
    LocalMux I__7605 (
            .O(N__33261),
            .I(N__33211));
    Span4Mux_v I__7604 (
            .O(N__33258),
            .I(N__33211));
    InMux I__7603 (
            .O(N__33257),
            .I(N__33206));
    InMux I__7602 (
            .O(N__33254),
            .I(N__33206));
    LocalMux I__7601 (
            .O(N__33247),
            .I(N__33201));
    LocalMux I__7600 (
            .O(N__33238),
            .I(N__33201));
    InMux I__7599 (
            .O(N__33237),
            .I(N__33194));
    InMux I__7598 (
            .O(N__33236),
            .I(N__33194));
    InMux I__7597 (
            .O(N__33235),
            .I(N__33194));
    Odrv4 I__7596 (
            .O(N__33232),
            .I(\POWERLED.count_clk_en ));
    Odrv12 I__7595 (
            .O(N__33229),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__7594 (
            .O(N__33224),
            .I(\POWERLED.count_clk_en ));
    Odrv12 I__7593 (
            .O(N__33221),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7592 (
            .O(N__33218),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__7591 (
            .O(N__33211),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7590 (
            .O(N__33206),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__7589 (
            .O(N__33201),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__7588 (
            .O(N__33194),
            .I(\POWERLED.count_clk_en ));
    CascadeMux I__7587 (
            .O(N__33175),
            .I(N__33171));
    InMux I__7586 (
            .O(N__33174),
            .I(N__33168));
    InMux I__7585 (
            .O(N__33171),
            .I(N__33165));
    LocalMux I__7584 (
            .O(N__33168),
            .I(\VPP_VDDQ.N_66_i ));
    LocalMux I__7583 (
            .O(N__33165),
            .I(\VPP_VDDQ.N_66_i ));
    CascadeMux I__7582 (
            .O(N__33160),
            .I(N__33156));
    InMux I__7581 (
            .O(N__33159),
            .I(N__33153));
    InMux I__7580 (
            .O(N__33156),
            .I(N__33150));
    LocalMux I__7579 (
            .O(N__33153),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__7578 (
            .O(N__33150),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    InMux I__7577 (
            .O(N__33145),
            .I(N__33141));
    InMux I__7576 (
            .O(N__33144),
            .I(N__33138));
    LocalMux I__7575 (
            .O(N__33141),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__7574 (
            .O(N__33138),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__7573 (
            .O(N__33133),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__7572 (
            .O(N__33130),
            .I(N__33126));
    InMux I__7571 (
            .O(N__33129),
            .I(N__33123));
    LocalMux I__7570 (
            .O(N__33126),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__7569 (
            .O(N__33123),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__7568 (
            .O(N__33118),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    CascadeMux I__7567 (
            .O(N__33115),
            .I(N__33111));
    InMux I__7566 (
            .O(N__33114),
            .I(N__33108));
    InMux I__7565 (
            .O(N__33111),
            .I(N__33105));
    LocalMux I__7564 (
            .O(N__33108),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__7563 (
            .O(N__33105),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__7562 (
            .O(N__33100),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__7561 (
            .O(N__33097),
            .I(N__33093));
    InMux I__7560 (
            .O(N__33096),
            .I(N__33090));
    LocalMux I__7559 (
            .O(N__33093),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__7558 (
            .O(N__33090),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__7557 (
            .O(N__33085),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__7556 (
            .O(N__33082),
            .I(N__33078));
    InMux I__7555 (
            .O(N__33081),
            .I(N__33075));
    LocalMux I__7554 (
            .O(N__33078),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__7553 (
            .O(N__33075),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__7552 (
            .O(N__33070),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__7551 (
            .O(N__33067),
            .I(N__33061));
    InMux I__7550 (
            .O(N__33066),
            .I(N__33061));
    LocalMux I__7549 (
            .O(N__33061),
            .I(N__33057));
    CascadeMux I__7548 (
            .O(N__33060),
            .I(N__33054));
    Span4Mux_v I__7547 (
            .O(N__33057),
            .I(N__33051));
    InMux I__7546 (
            .O(N__33054),
            .I(N__33048));
    Odrv4 I__7545 (
            .O(N__33051),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__7544 (
            .O(N__33048),
            .I(\POWERLED.count_clkZ0Z_3 ));
    CascadeMux I__7543 (
            .O(N__33043),
            .I(N__33040));
    InMux I__7542 (
            .O(N__33040),
            .I(N__33036));
    InMux I__7541 (
            .O(N__33039),
            .I(N__33033));
    LocalMux I__7540 (
            .O(N__33036),
            .I(N__33030));
    LocalMux I__7539 (
            .O(N__33033),
            .I(\POWERLED.count_clkZ0Z_10 ));
    Odrv4 I__7538 (
            .O(N__33030),
            .I(\POWERLED.count_clkZ0Z_10 ));
    CascadeMux I__7537 (
            .O(N__33025),
            .I(N__33021));
    CascadeMux I__7536 (
            .O(N__33024),
            .I(N__33015));
    InMux I__7535 (
            .O(N__33021),
            .I(N__33011));
    CascadeMux I__7534 (
            .O(N__33020),
            .I(N__33008));
    InMux I__7533 (
            .O(N__33019),
            .I(N__33005));
    InMux I__7532 (
            .O(N__33018),
            .I(N__33002));
    InMux I__7531 (
            .O(N__33015),
            .I(N__32997));
    InMux I__7530 (
            .O(N__33014),
            .I(N__32997));
    LocalMux I__7529 (
            .O(N__33011),
            .I(N__32994));
    InMux I__7528 (
            .O(N__33008),
            .I(N__32991));
    LocalMux I__7527 (
            .O(N__33005),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__7526 (
            .O(N__33002),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__7525 (
            .O(N__32997),
            .I(\POWERLED.count_clkZ0Z_1 ));
    Odrv4 I__7524 (
            .O(N__32994),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__7523 (
            .O(N__32991),
            .I(\POWERLED.count_clkZ0Z_1 ));
    CascadeMux I__7522 (
            .O(N__32980),
            .I(\POWERLED.un2_count_clk_15_0_9_cascade_ ));
    InMux I__7521 (
            .O(N__32977),
            .I(N__32974));
    LocalMux I__7520 (
            .O(N__32974),
            .I(\POWERLED.un2_count_clk_15_0_8 ));
    InMux I__7519 (
            .O(N__32971),
            .I(N__32960));
    CascadeMux I__7518 (
            .O(N__32970),
            .I(N__32957));
    InMux I__7517 (
            .O(N__32969),
            .I(N__32953));
    InMux I__7516 (
            .O(N__32968),
            .I(N__32948));
    CascadeMux I__7515 (
            .O(N__32967),
            .I(N__32945));
    InMux I__7514 (
            .O(N__32966),
            .I(N__32939));
    InMux I__7513 (
            .O(N__32965),
            .I(N__32939));
    InMux I__7512 (
            .O(N__32964),
            .I(N__32934));
    InMux I__7511 (
            .O(N__32963),
            .I(N__32934));
    LocalMux I__7510 (
            .O(N__32960),
            .I(N__32931));
    InMux I__7509 (
            .O(N__32957),
            .I(N__32928));
    InMux I__7508 (
            .O(N__32956),
            .I(N__32925));
    LocalMux I__7507 (
            .O(N__32953),
            .I(N__32922));
    InMux I__7506 (
            .O(N__32952),
            .I(N__32919));
    InMux I__7505 (
            .O(N__32951),
            .I(N__32916));
    LocalMux I__7504 (
            .O(N__32948),
            .I(N__32912));
    InMux I__7503 (
            .O(N__32945),
            .I(N__32909));
    InMux I__7502 (
            .O(N__32944),
            .I(N__32906));
    LocalMux I__7501 (
            .O(N__32939),
            .I(N__32901));
    LocalMux I__7500 (
            .O(N__32934),
            .I(N__32901));
    Span4Mux_v I__7499 (
            .O(N__32931),
            .I(N__32898));
    LocalMux I__7498 (
            .O(N__32928),
            .I(N__32893));
    LocalMux I__7497 (
            .O(N__32925),
            .I(N__32893));
    Span4Mux_v I__7496 (
            .O(N__32922),
            .I(N__32886));
    LocalMux I__7495 (
            .O(N__32919),
            .I(N__32886));
    LocalMux I__7494 (
            .O(N__32916),
            .I(N__32886));
    InMux I__7493 (
            .O(N__32915),
            .I(N__32883));
    Span4Mux_v I__7492 (
            .O(N__32912),
            .I(N__32877));
    LocalMux I__7491 (
            .O(N__32909),
            .I(N__32877));
    LocalMux I__7490 (
            .O(N__32906),
            .I(N__32874));
    Span4Mux_v I__7489 (
            .O(N__32901),
            .I(N__32867));
    Span4Mux_v I__7488 (
            .O(N__32898),
            .I(N__32867));
    Span4Mux_v I__7487 (
            .O(N__32893),
            .I(N__32867));
    Span4Mux_v I__7486 (
            .O(N__32886),
            .I(N__32862));
    LocalMux I__7485 (
            .O(N__32883),
            .I(N__32862));
    InMux I__7484 (
            .O(N__32882),
            .I(N__32859));
    Span4Mux_h I__7483 (
            .O(N__32877),
            .I(N__32854));
    Span4Mux_h I__7482 (
            .O(N__32874),
            .I(N__32854));
    Span4Mux_h I__7481 (
            .O(N__32867),
            .I(N__32849));
    Span4Mux_h I__7480 (
            .O(N__32862),
            .I(N__32849));
    LocalMux I__7479 (
            .O(N__32859),
            .I(\POWERLED.un2_count_clk_15_1 ));
    Odrv4 I__7478 (
            .O(N__32854),
            .I(\POWERLED.un2_count_clk_15_1 ));
    Odrv4 I__7477 (
            .O(N__32849),
            .I(\POWERLED.un2_count_clk_15_1 ));
    InMux I__7476 (
            .O(N__32842),
            .I(N__32837));
    InMux I__7475 (
            .O(N__32841),
            .I(N__32832));
    InMux I__7474 (
            .O(N__32840),
            .I(N__32832));
    LocalMux I__7473 (
            .O(N__32837),
            .I(N__32829));
    LocalMux I__7472 (
            .O(N__32832),
            .I(\POWERLED.count_clkZ0Z_8 ));
    Odrv4 I__7471 (
            .O(N__32829),
            .I(\POWERLED.count_clkZ0Z_8 ));
    CascadeMux I__7470 (
            .O(N__32824),
            .I(N__32818));
    InMux I__7469 (
            .O(N__32823),
            .I(N__32813));
    InMux I__7468 (
            .O(N__32822),
            .I(N__32813));
    InMux I__7467 (
            .O(N__32821),
            .I(N__32810));
    InMux I__7466 (
            .O(N__32818),
            .I(N__32807));
    LocalMux I__7465 (
            .O(N__32813),
            .I(N__32804));
    LocalMux I__7464 (
            .O(N__32810),
            .I(N__32801));
    LocalMux I__7463 (
            .O(N__32807),
            .I(N__32798));
    Span4Mux_v I__7462 (
            .O(N__32804),
            .I(N__32795));
    Span4Mux_s2_h I__7461 (
            .O(N__32801),
            .I(N__32792));
    Span4Mux_s2_h I__7460 (
            .O(N__32798),
            .I(N__32789));
    Odrv4 I__7459 (
            .O(N__32795),
            .I(\POWERLED.count_clkZ0Z_9 ));
    Odrv4 I__7458 (
            .O(N__32792),
            .I(\POWERLED.count_clkZ0Z_9 ));
    Odrv4 I__7457 (
            .O(N__32789),
            .I(\POWERLED.count_clkZ0Z_9 ));
    InMux I__7456 (
            .O(N__32782),
            .I(N__32779));
    LocalMux I__7455 (
            .O(N__32779),
            .I(\POWERLED.un2_count_clk_15_0_10 ));
    InMux I__7454 (
            .O(N__32776),
            .I(N__32773));
    LocalMux I__7453 (
            .O(N__32773),
            .I(N__32770));
    Odrv12 I__7452 (
            .O(N__32770),
            .I(\POWERLED.count_clk_0_12 ));
    InMux I__7451 (
            .O(N__32767),
            .I(N__32763));
    InMux I__7450 (
            .O(N__32766),
            .I(N__32760));
    LocalMux I__7449 (
            .O(N__32763),
            .I(N__32757));
    LocalMux I__7448 (
            .O(N__32760),
            .I(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ));
    Odrv4 I__7447 (
            .O(N__32757),
            .I(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ));
    CascadeMux I__7446 (
            .O(N__32752),
            .I(N__32749));
    InMux I__7445 (
            .O(N__32749),
            .I(N__32746));
    LocalMux I__7444 (
            .O(N__32746),
            .I(N__32743));
    Odrv4 I__7443 (
            .O(N__32743),
            .I(\POWERLED.count_clkZ0Z_12 ));
    CascadeMux I__7442 (
            .O(N__32740),
            .I(\POWERLED.count_clkZ0Z_12_cascade_ ));
    CascadeMux I__7441 (
            .O(N__32737),
            .I(N__32732));
    InMux I__7440 (
            .O(N__32736),
            .I(N__32729));
    InMux I__7439 (
            .O(N__32735),
            .I(N__32723));
    InMux I__7438 (
            .O(N__32732),
            .I(N__32723));
    LocalMux I__7437 (
            .O(N__32729),
            .I(N__32720));
    CascadeMux I__7436 (
            .O(N__32728),
            .I(N__32717));
    LocalMux I__7435 (
            .O(N__32723),
            .I(N__32714));
    Span4Mux_s3_h I__7434 (
            .O(N__32720),
            .I(N__32711));
    InMux I__7433 (
            .O(N__32717),
            .I(N__32708));
    Span4Mux_s2_h I__7432 (
            .O(N__32714),
            .I(N__32705));
    Span4Mux_v I__7431 (
            .O(N__32711),
            .I(N__32700));
    LocalMux I__7430 (
            .O(N__32708),
            .I(N__32700));
    Odrv4 I__7429 (
            .O(N__32705),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__7428 (
            .O(N__32700),
            .I(\POWERLED.count_clkZ0Z_7 ));
    CascadeMux I__7427 (
            .O(N__32695),
            .I(\POWERLED.count_clk_RNIZ0Z_12_cascade_ ));
    CascadeMux I__7426 (
            .O(N__32692),
            .I(N__32689));
    InMux I__7425 (
            .O(N__32689),
            .I(N__32686));
    LocalMux I__7424 (
            .O(N__32686),
            .I(\POWERLED.un2_count_clk_15_0_7 ));
    CascadeMux I__7423 (
            .O(N__32683),
            .I(N__32680));
    InMux I__7422 (
            .O(N__32680),
            .I(N__32675));
    InMux I__7421 (
            .O(N__32679),
            .I(N__32672));
    InMux I__7420 (
            .O(N__32678),
            .I(N__32669));
    LocalMux I__7419 (
            .O(N__32675),
            .I(N__32666));
    LocalMux I__7418 (
            .O(N__32672),
            .I(\POWERLED.count_clkZ0Z_11 ));
    LocalMux I__7417 (
            .O(N__32669),
            .I(\POWERLED.count_clkZ0Z_11 ));
    Odrv4 I__7416 (
            .O(N__32666),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__7415 (
            .O(N__32659),
            .I(N__32653));
    InMux I__7414 (
            .O(N__32658),
            .I(N__32653));
    LocalMux I__7413 (
            .O(N__32653),
            .I(N__32650));
    Span4Mux_v I__7412 (
            .O(N__32650),
            .I(N__32647));
    Odrv4 I__7411 (
            .O(N__32647),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    CascadeMux I__7410 (
            .O(N__32644),
            .I(N__32641));
    InMux I__7409 (
            .O(N__32641),
            .I(N__32638));
    LocalMux I__7408 (
            .O(N__32638),
            .I(\POWERLED.count_clk_0_2 ));
    CascadeMux I__7407 (
            .O(N__32635),
            .I(N__32632));
    InMux I__7406 (
            .O(N__32632),
            .I(N__32628));
    InMux I__7405 (
            .O(N__32631),
            .I(N__32625));
    LocalMux I__7404 (
            .O(N__32628),
            .I(N__32622));
    LocalMux I__7403 (
            .O(N__32625),
            .I(\POWERLED.count_clkZ0Z_2 ));
    Odrv12 I__7402 (
            .O(N__32622),
            .I(\POWERLED.count_clkZ0Z_2 ));
    CascadeMux I__7401 (
            .O(N__32617),
            .I(\POWERLED.count_clkZ0Z_15_cascade_ ));
    InMux I__7400 (
            .O(N__32614),
            .I(N__32607));
    InMux I__7399 (
            .O(N__32613),
            .I(N__32602));
    InMux I__7398 (
            .O(N__32612),
            .I(N__32602));
    InMux I__7397 (
            .O(N__32611),
            .I(N__32599));
    InMux I__7396 (
            .O(N__32610),
            .I(N__32596));
    LocalMux I__7395 (
            .O(N__32607),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__7394 (
            .O(N__32602),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__7393 (
            .O(N__32599),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__7392 (
            .O(N__32596),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__7391 (
            .O(N__32587),
            .I(N__32584));
    LocalMux I__7390 (
            .O(N__32584),
            .I(\POWERLED.count_clk_0_1 ));
    InMux I__7389 (
            .O(N__32581),
            .I(N__32575));
    InMux I__7388 (
            .O(N__32580),
            .I(N__32575));
    LocalMux I__7387 (
            .O(N__32575),
            .I(N__32572));
    Odrv4 I__7386 (
            .O(N__32572),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    InMux I__7385 (
            .O(N__32569),
            .I(N__32566));
    LocalMux I__7384 (
            .O(N__32566),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__7383 (
            .O(N__32563),
            .I(N__32560));
    LocalMux I__7382 (
            .O(N__32560),
            .I(\POWERLED.count_clk_0_10 ));
    InMux I__7381 (
            .O(N__32557),
            .I(N__32551));
    InMux I__7380 (
            .O(N__32556),
            .I(N__32551));
    LocalMux I__7379 (
            .O(N__32551),
            .I(N__32548));
    Odrv4 I__7378 (
            .O(N__32548),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    InMux I__7377 (
            .O(N__32545),
            .I(N__32541));
    CascadeMux I__7376 (
            .O(N__32544),
            .I(N__32537));
    LocalMux I__7375 (
            .O(N__32541),
            .I(N__32534));
    InMux I__7374 (
            .O(N__32540),
            .I(N__32531));
    InMux I__7373 (
            .O(N__32537),
            .I(N__32528));
    Odrv4 I__7372 (
            .O(N__32534),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__7371 (
            .O(N__32531),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__7370 (
            .O(N__32528),
            .I(\POWERLED.count_clkZ0Z_6 ));
    CascadeMux I__7369 (
            .O(N__32521),
            .I(\POWERLED.count_clkZ0Z_10_cascade_ ));
    InMux I__7368 (
            .O(N__32518),
            .I(N__32515));
    LocalMux I__7367 (
            .O(N__32515),
            .I(N__32511));
    InMux I__7366 (
            .O(N__32514),
            .I(N__32508));
    Span4Mux_s1_h I__7365 (
            .O(N__32511),
            .I(N__32503));
    LocalMux I__7364 (
            .O(N__32508),
            .I(N__32503));
    Odrv4 I__7363 (
            .O(N__32503),
            .I(\POWERLED.count_clk_RNIZ0Z_13 ));
    CascadeMux I__7362 (
            .O(N__32500),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_cascade_ ));
    InMux I__7361 (
            .O(N__32497),
            .I(N__32485));
    InMux I__7360 (
            .O(N__32496),
            .I(N__32485));
    InMux I__7359 (
            .O(N__32495),
            .I(N__32485));
    InMux I__7358 (
            .O(N__32494),
            .I(N__32485));
    LocalMux I__7357 (
            .O(N__32485),
            .I(N__32481));
    InMux I__7356 (
            .O(N__32484),
            .I(N__32478));
    Odrv4 I__7355 (
            .O(N__32481),
            .I(\POWERLED.N_352 ));
    LocalMux I__7354 (
            .O(N__32478),
            .I(\POWERLED.N_352 ));
    InMux I__7353 (
            .O(N__32473),
            .I(\POWERLED.un1_count_clk_2_cry_11 ));
    CascadeMux I__7352 (
            .O(N__32470),
            .I(N__32466));
    InMux I__7351 (
            .O(N__32469),
            .I(N__32463));
    InMux I__7350 (
            .O(N__32466),
            .I(N__32460));
    LocalMux I__7349 (
            .O(N__32463),
            .I(\POWERLED.count_clkZ0Z_13 ));
    LocalMux I__7348 (
            .O(N__32460),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__7347 (
            .O(N__32455),
            .I(N__32449));
    InMux I__7346 (
            .O(N__32454),
            .I(N__32449));
    LocalMux I__7345 (
            .O(N__32449),
            .I(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ));
    InMux I__7344 (
            .O(N__32446),
            .I(\POWERLED.un1_count_clk_2_cry_12 ));
    CascadeMux I__7343 (
            .O(N__32443),
            .I(N__32440));
    InMux I__7342 (
            .O(N__32440),
            .I(N__32437));
    LocalMux I__7341 (
            .O(N__32437),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__7340 (
            .O(N__32434),
            .I(N__32428));
    InMux I__7339 (
            .O(N__32433),
            .I(N__32428));
    LocalMux I__7338 (
            .O(N__32428),
            .I(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ));
    InMux I__7337 (
            .O(N__32425),
            .I(\POWERLED.un1_count_clk_2_cry_13 ));
    InMux I__7336 (
            .O(N__32422),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    CascadeMux I__7335 (
            .O(N__32419),
            .I(N__32415));
    CascadeMux I__7334 (
            .O(N__32418),
            .I(N__32410));
    InMux I__7333 (
            .O(N__32415),
            .I(N__32407));
    InMux I__7332 (
            .O(N__32414),
            .I(N__32402));
    InMux I__7331 (
            .O(N__32413),
            .I(N__32402));
    InMux I__7330 (
            .O(N__32410),
            .I(N__32399));
    LocalMux I__7329 (
            .O(N__32407),
            .I(N__32396));
    LocalMux I__7328 (
            .O(N__32402),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__7327 (
            .O(N__32399),
            .I(\POWERLED.count_clkZ0Z_5 ));
    Odrv4 I__7326 (
            .O(N__32396),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__7325 (
            .O(N__32389),
            .I(N__32383));
    InMux I__7324 (
            .O(N__32388),
            .I(N__32383));
    LocalMux I__7323 (
            .O(N__32383),
            .I(N__32380));
    Odrv4 I__7322 (
            .O(N__32380),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    InMux I__7321 (
            .O(N__32377),
            .I(N__32374));
    LocalMux I__7320 (
            .O(N__32374),
            .I(\POWERLED.count_clk_0_5 ));
    InMux I__7319 (
            .O(N__32371),
            .I(N__32368));
    LocalMux I__7318 (
            .O(N__32368),
            .I(\POWERLED.count_clk_0_15 ));
    InMux I__7317 (
            .O(N__32365),
            .I(N__32359));
    InMux I__7316 (
            .O(N__32364),
            .I(N__32359));
    LocalMux I__7315 (
            .O(N__32359),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    InMux I__7314 (
            .O(N__32356),
            .I(N__32353));
    LocalMux I__7313 (
            .O(N__32353),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__7312 (
            .O(N__32350),
            .I(N__32346));
    InMux I__7311 (
            .O(N__32349),
            .I(N__32343));
    LocalMux I__7310 (
            .O(N__32346),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    LocalMux I__7309 (
            .O(N__32343),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    InMux I__7308 (
            .O(N__32338),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    InMux I__7307 (
            .O(N__32335),
            .I(N__32331));
    InMux I__7306 (
            .O(N__32334),
            .I(N__32328));
    LocalMux I__7305 (
            .O(N__32331),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    LocalMux I__7304 (
            .O(N__32328),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    InMux I__7303 (
            .O(N__32323),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__7302 (
            .O(N__32320),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__7301 (
            .O(N__32317),
            .I(N__32311));
    InMux I__7300 (
            .O(N__32316),
            .I(N__32311));
    LocalMux I__7299 (
            .O(N__32311),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    InMux I__7298 (
            .O(N__32308),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    CascadeMux I__7297 (
            .O(N__32305),
            .I(N__32301));
    InMux I__7296 (
            .O(N__32304),
            .I(N__32296));
    InMux I__7295 (
            .O(N__32301),
            .I(N__32296));
    LocalMux I__7294 (
            .O(N__32296),
            .I(N__32293));
    Odrv4 I__7293 (
            .O(N__32293),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    InMux I__7292 (
            .O(N__32290),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__7291 (
            .O(N__32287),
            .I(\POWERLED.un1_count_clk_2_cry_7 ));
    CascadeMux I__7290 (
            .O(N__32284),
            .I(N__32280));
    InMux I__7289 (
            .O(N__32283),
            .I(N__32275));
    InMux I__7288 (
            .O(N__32280),
            .I(N__32275));
    LocalMux I__7287 (
            .O(N__32275),
            .I(N__32272));
    Span4Mux_v I__7286 (
            .O(N__32272),
            .I(N__32269));
    Odrv4 I__7285 (
            .O(N__32269),
            .I(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ));
    InMux I__7284 (
            .O(N__32266),
            .I(bfn_12_10_0_));
    InMux I__7283 (
            .O(N__32263),
            .I(\POWERLED.un1_count_clk_2_cry_9 ));
    InMux I__7282 (
            .O(N__32260),
            .I(\POWERLED.un1_count_clk_2_cry_10 ));
    InMux I__7281 (
            .O(N__32257),
            .I(N__32251));
    InMux I__7280 (
            .O(N__32256),
            .I(N__32251));
    LocalMux I__7279 (
            .O(N__32251),
            .I(\VPP_VDDQ.count_2_1_1 ));
    InMux I__7278 (
            .O(N__32248),
            .I(N__32245));
    LocalMux I__7277 (
            .O(N__32245),
            .I(N__32242));
    Odrv4 I__7276 (
            .O(N__32242),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1 ));
    CascadeMux I__7275 (
            .O(N__32239),
            .I(\VPP_VDDQ.un1_count_2_1_axb_1_cascade_ ));
    CascadeMux I__7274 (
            .O(N__32236),
            .I(N__32232));
    CascadeMux I__7273 (
            .O(N__32235),
            .I(N__32229));
    InMux I__7272 (
            .O(N__32232),
            .I(N__32224));
    InMux I__7271 (
            .O(N__32229),
            .I(N__32221));
    InMux I__7270 (
            .O(N__32228),
            .I(N__32216));
    InMux I__7269 (
            .O(N__32227),
            .I(N__32216));
    LocalMux I__7268 (
            .O(N__32224),
            .I(N__32213));
    LocalMux I__7267 (
            .O(N__32221),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__7266 (
            .O(N__32216),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    Odrv12 I__7265 (
            .O(N__32213),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    CascadeMux I__7264 (
            .O(N__32206),
            .I(N__32203));
    InMux I__7263 (
            .O(N__32203),
            .I(N__32200));
    LocalMux I__7262 (
            .O(N__32200),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1 ));
    CascadeMux I__7261 (
            .O(N__32197),
            .I(\VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ));
    CascadeMux I__7260 (
            .O(N__32194),
            .I(N__32191));
    InMux I__7259 (
            .O(N__32191),
            .I(N__32185));
    InMux I__7258 (
            .O(N__32190),
            .I(N__32185));
    LocalMux I__7257 (
            .O(N__32185),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    CascadeMux I__7256 (
            .O(N__32182),
            .I(N__32178));
    CascadeMux I__7255 (
            .O(N__32181),
            .I(N__32174));
    InMux I__7254 (
            .O(N__32178),
            .I(N__32155));
    InMux I__7253 (
            .O(N__32177),
            .I(N__32155));
    InMux I__7252 (
            .O(N__32174),
            .I(N__32155));
    InMux I__7251 (
            .O(N__32173),
            .I(N__32155));
    InMux I__7250 (
            .O(N__32172),
            .I(N__32143));
    InMux I__7249 (
            .O(N__32171),
            .I(N__32130));
    InMux I__7248 (
            .O(N__32170),
            .I(N__32130));
    InMux I__7247 (
            .O(N__32169),
            .I(N__32130));
    InMux I__7246 (
            .O(N__32168),
            .I(N__32130));
    InMux I__7245 (
            .O(N__32167),
            .I(N__32130));
    InMux I__7244 (
            .O(N__32166),
            .I(N__32130));
    InMux I__7243 (
            .O(N__32165),
            .I(N__32127));
    InMux I__7242 (
            .O(N__32164),
            .I(N__32124));
    LocalMux I__7241 (
            .O(N__32155),
            .I(N__32121));
    InMux I__7240 (
            .O(N__32154),
            .I(N__32112));
    InMux I__7239 (
            .O(N__32153),
            .I(N__32112));
    InMux I__7238 (
            .O(N__32152),
            .I(N__32112));
    InMux I__7237 (
            .O(N__32151),
            .I(N__32112));
    CascadeMux I__7236 (
            .O(N__32150),
            .I(N__32108));
    InMux I__7235 (
            .O(N__32149),
            .I(N__32098));
    InMux I__7234 (
            .O(N__32148),
            .I(N__32098));
    InMux I__7233 (
            .O(N__32147),
            .I(N__32098));
    InMux I__7232 (
            .O(N__32146),
            .I(N__32098));
    LocalMux I__7231 (
            .O(N__32143),
            .I(N__32095));
    LocalMux I__7230 (
            .O(N__32130),
            .I(N__32092));
    LocalMux I__7229 (
            .O(N__32127),
            .I(N__32074));
    LocalMux I__7228 (
            .O(N__32124),
            .I(N__32074));
    Span4Mux_h I__7227 (
            .O(N__32121),
            .I(N__32074));
    LocalMux I__7226 (
            .O(N__32112),
            .I(N__32074));
    CascadeMux I__7225 (
            .O(N__32111),
            .I(N__32070));
    InMux I__7224 (
            .O(N__32108),
            .I(N__32065));
    InMux I__7223 (
            .O(N__32107),
            .I(N__32062));
    LocalMux I__7222 (
            .O(N__32098),
            .I(N__32059));
    Span4Mux_v I__7221 (
            .O(N__32095),
            .I(N__32056));
    Span4Mux_h I__7220 (
            .O(N__32092),
            .I(N__32053));
    InMux I__7219 (
            .O(N__32091),
            .I(N__32044));
    InMux I__7218 (
            .O(N__32090),
            .I(N__32044));
    InMux I__7217 (
            .O(N__32089),
            .I(N__32044));
    InMux I__7216 (
            .O(N__32088),
            .I(N__32044));
    InMux I__7215 (
            .O(N__32087),
            .I(N__32033));
    InMux I__7214 (
            .O(N__32086),
            .I(N__32033));
    InMux I__7213 (
            .O(N__32085),
            .I(N__32033));
    InMux I__7212 (
            .O(N__32084),
            .I(N__32033));
    InMux I__7211 (
            .O(N__32083),
            .I(N__32033));
    Span4Mux_v I__7210 (
            .O(N__32074),
            .I(N__32030));
    InMux I__7209 (
            .O(N__32073),
            .I(N__32021));
    InMux I__7208 (
            .O(N__32070),
            .I(N__32021));
    InMux I__7207 (
            .O(N__32069),
            .I(N__32021));
    InMux I__7206 (
            .O(N__32068),
            .I(N__32021));
    LocalMux I__7205 (
            .O(N__32065),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7204 (
            .O(N__32062),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7203 (
            .O(N__32059),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7202 (
            .O(N__32056),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7201 (
            .O(N__32053),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7200 (
            .O(N__32044),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7199 (
            .O(N__32033),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7198 (
            .O(N__32030),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7197 (
            .O(N__32021),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    CascadeMux I__7196 (
            .O(N__32002),
            .I(N__31998));
    InMux I__7195 (
            .O(N__32001),
            .I(N__31993));
    InMux I__7194 (
            .O(N__31998),
            .I(N__31993));
    LocalMux I__7193 (
            .O(N__31993),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ));
    CascadeMux I__7192 (
            .O(N__31990),
            .I(N__31985));
    CascadeMux I__7191 (
            .O(N__31989),
            .I(N__31976));
    InMux I__7190 (
            .O(N__31988),
            .I(N__31968));
    InMux I__7189 (
            .O(N__31985),
            .I(N__31957));
    InMux I__7188 (
            .O(N__31984),
            .I(N__31957));
    InMux I__7187 (
            .O(N__31983),
            .I(N__31957));
    InMux I__7186 (
            .O(N__31982),
            .I(N__31957));
    InMux I__7185 (
            .O(N__31981),
            .I(N__31957));
    InMux I__7184 (
            .O(N__31980),
            .I(N__31954));
    CascadeMux I__7183 (
            .O(N__31979),
            .I(N__31944));
    InMux I__7182 (
            .O(N__31976),
            .I(N__31936));
    InMux I__7181 (
            .O(N__31975),
            .I(N__31936));
    InMux I__7180 (
            .O(N__31974),
            .I(N__31931));
    InMux I__7179 (
            .O(N__31973),
            .I(N__31931));
    CascadeMux I__7178 (
            .O(N__31972),
            .I(N__31928));
    InMux I__7177 (
            .O(N__31971),
            .I(N__31922));
    LocalMux I__7176 (
            .O(N__31968),
            .I(N__31915));
    LocalMux I__7175 (
            .O(N__31957),
            .I(N__31915));
    LocalMux I__7174 (
            .O(N__31954),
            .I(N__31915));
    CascadeMux I__7173 (
            .O(N__31953),
            .I(N__31903));
    InMux I__7172 (
            .O(N__31952),
            .I(N__31898));
    InMux I__7171 (
            .O(N__31951),
            .I(N__31889));
    InMux I__7170 (
            .O(N__31950),
            .I(N__31889));
    InMux I__7169 (
            .O(N__31949),
            .I(N__31889));
    InMux I__7168 (
            .O(N__31948),
            .I(N__31889));
    InMux I__7167 (
            .O(N__31947),
            .I(N__31884));
    InMux I__7166 (
            .O(N__31944),
            .I(N__31884));
    InMux I__7165 (
            .O(N__31943),
            .I(N__31881));
    InMux I__7164 (
            .O(N__31942),
            .I(N__31876));
    InMux I__7163 (
            .O(N__31941),
            .I(N__31876));
    LocalMux I__7162 (
            .O(N__31936),
            .I(N__31871));
    LocalMux I__7161 (
            .O(N__31931),
            .I(N__31871));
    InMux I__7160 (
            .O(N__31928),
            .I(N__31866));
    InMux I__7159 (
            .O(N__31927),
            .I(N__31866));
    InMux I__7158 (
            .O(N__31926),
            .I(N__31861));
    InMux I__7157 (
            .O(N__31925),
            .I(N__31861));
    LocalMux I__7156 (
            .O(N__31922),
            .I(N__31856));
    Span4Mux_v I__7155 (
            .O(N__31915),
            .I(N__31856));
    InMux I__7154 (
            .O(N__31914),
            .I(N__31845));
    InMux I__7153 (
            .O(N__31913),
            .I(N__31845));
    InMux I__7152 (
            .O(N__31912),
            .I(N__31845));
    InMux I__7151 (
            .O(N__31911),
            .I(N__31845));
    InMux I__7150 (
            .O(N__31910),
            .I(N__31845));
    InMux I__7149 (
            .O(N__31909),
            .I(N__31836));
    InMux I__7148 (
            .O(N__31908),
            .I(N__31836));
    InMux I__7147 (
            .O(N__31907),
            .I(N__31836));
    InMux I__7146 (
            .O(N__31906),
            .I(N__31836));
    InMux I__7145 (
            .O(N__31903),
            .I(N__31829));
    InMux I__7144 (
            .O(N__31902),
            .I(N__31829));
    InMux I__7143 (
            .O(N__31901),
            .I(N__31829));
    LocalMux I__7142 (
            .O(N__31898),
            .I(N__31824));
    LocalMux I__7141 (
            .O(N__31889),
            .I(N__31824));
    LocalMux I__7140 (
            .O(N__31884),
            .I(N__31815));
    LocalMux I__7139 (
            .O(N__31881),
            .I(N__31815));
    LocalMux I__7138 (
            .O(N__31876),
            .I(N__31815));
    Span4Mux_v I__7137 (
            .O(N__31871),
            .I(N__31815));
    LocalMux I__7136 (
            .O(N__31866),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7135 (
            .O(N__31861),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__7134 (
            .O(N__31856),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7133 (
            .O(N__31845),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7132 (
            .O(N__31836),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    LocalMux I__7131 (
            .O(N__31829),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv12 I__7130 (
            .O(N__31824),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__7129 (
            .O(N__31815),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    InMux I__7128 (
            .O(N__31798),
            .I(N__31787));
    CascadeMux I__7127 (
            .O(N__31797),
            .I(N__31771));
    CascadeMux I__7126 (
            .O(N__31796),
            .I(N__31767));
    InMux I__7125 (
            .O(N__31795),
            .I(N__31749));
    InMux I__7124 (
            .O(N__31794),
            .I(N__31749));
    InMux I__7123 (
            .O(N__31793),
            .I(N__31749));
    InMux I__7122 (
            .O(N__31792),
            .I(N__31749));
    InMux I__7121 (
            .O(N__31791),
            .I(N__31749));
    InMux I__7120 (
            .O(N__31790),
            .I(N__31749));
    LocalMux I__7119 (
            .O(N__31787),
            .I(N__31739));
    InMux I__7118 (
            .O(N__31786),
            .I(N__31730));
    InMux I__7117 (
            .O(N__31785),
            .I(N__31730));
    InMux I__7116 (
            .O(N__31784),
            .I(N__31730));
    InMux I__7115 (
            .O(N__31783),
            .I(N__31730));
    InMux I__7114 (
            .O(N__31782),
            .I(N__31721));
    InMux I__7113 (
            .O(N__31781),
            .I(N__31721));
    InMux I__7112 (
            .O(N__31780),
            .I(N__31721));
    InMux I__7111 (
            .O(N__31779),
            .I(N__31721));
    InMux I__7110 (
            .O(N__31778),
            .I(N__31710));
    InMux I__7109 (
            .O(N__31777),
            .I(N__31710));
    InMux I__7108 (
            .O(N__31776),
            .I(N__31710));
    InMux I__7107 (
            .O(N__31775),
            .I(N__31710));
    InMux I__7106 (
            .O(N__31774),
            .I(N__31710));
    InMux I__7105 (
            .O(N__31771),
            .I(N__31707));
    InMux I__7104 (
            .O(N__31770),
            .I(N__31702));
    InMux I__7103 (
            .O(N__31767),
            .I(N__31702));
    InMux I__7102 (
            .O(N__31766),
            .I(N__31699));
    InMux I__7101 (
            .O(N__31765),
            .I(N__31690));
    InMux I__7100 (
            .O(N__31764),
            .I(N__31690));
    InMux I__7099 (
            .O(N__31763),
            .I(N__31690));
    InMux I__7098 (
            .O(N__31762),
            .I(N__31690));
    LocalMux I__7097 (
            .O(N__31749),
            .I(N__31687));
    InMux I__7096 (
            .O(N__31748),
            .I(N__31680));
    InMux I__7095 (
            .O(N__31747),
            .I(N__31680));
    InMux I__7094 (
            .O(N__31746),
            .I(N__31680));
    InMux I__7093 (
            .O(N__31745),
            .I(N__31671));
    InMux I__7092 (
            .O(N__31744),
            .I(N__31671));
    InMux I__7091 (
            .O(N__31743),
            .I(N__31671));
    InMux I__7090 (
            .O(N__31742),
            .I(N__31671));
    Span4Mux_h I__7089 (
            .O(N__31739),
            .I(N__31664));
    LocalMux I__7088 (
            .O(N__31730),
            .I(N__31664));
    LocalMux I__7087 (
            .O(N__31721),
            .I(N__31664));
    LocalMux I__7086 (
            .O(N__31710),
            .I(N__31661));
    LocalMux I__7085 (
            .O(N__31707),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7084 (
            .O(N__31702),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7083 (
            .O(N__31699),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7082 (
            .O(N__31690),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7081 (
            .O(N__31687),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7080 (
            .O(N__31680),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7079 (
            .O(N__31671),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7078 (
            .O(N__31664),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7077 (
            .O(N__31661),
            .I(\VPP_VDDQ.N_1_i ));
    InMux I__7076 (
            .O(N__31642),
            .I(N__31639));
    LocalMux I__7075 (
            .O(N__31639),
            .I(\VPP_VDDQ.count_2_0_11 ));
    CascadeMux I__7074 (
            .O(N__31636),
            .I(\VPP_VDDQ.count_2_1_11_cascade_ ));
    CEMux I__7073 (
            .O(N__31633),
            .I(N__31628));
    CEMux I__7072 (
            .O(N__31632),
            .I(N__31623));
    CEMux I__7071 (
            .O(N__31631),
            .I(N__31615));
    LocalMux I__7070 (
            .O(N__31628),
            .I(N__31612));
    InMux I__7069 (
            .O(N__31627),
            .I(N__31607));
    InMux I__7068 (
            .O(N__31626),
            .I(N__31607));
    LocalMux I__7067 (
            .O(N__31623),
            .I(N__31601));
    CEMux I__7066 (
            .O(N__31622),
            .I(N__31598));
    CEMux I__7065 (
            .O(N__31621),
            .I(N__31595));
    InMux I__7064 (
            .O(N__31620),
            .I(N__31591));
    InMux I__7063 (
            .O(N__31619),
            .I(N__31584));
    InMux I__7062 (
            .O(N__31618),
            .I(N__31584));
    LocalMux I__7061 (
            .O(N__31615),
            .I(N__31577));
    Span4Mux_v I__7060 (
            .O(N__31612),
            .I(N__31577));
    LocalMux I__7059 (
            .O(N__31607),
            .I(N__31577));
    InMux I__7058 (
            .O(N__31606),
            .I(N__31570));
    InMux I__7057 (
            .O(N__31605),
            .I(N__31570));
    InMux I__7056 (
            .O(N__31604),
            .I(N__31570));
    Span4Mux_h I__7055 (
            .O(N__31601),
            .I(N__31559));
    LocalMux I__7054 (
            .O(N__31598),
            .I(N__31559));
    LocalMux I__7053 (
            .O(N__31595),
            .I(N__31559));
    CEMux I__7052 (
            .O(N__31594),
            .I(N__31556));
    LocalMux I__7051 (
            .O(N__31591),
            .I(N__31553));
    InMux I__7050 (
            .O(N__31590),
            .I(N__31542));
    InMux I__7049 (
            .O(N__31589),
            .I(N__31542));
    LocalMux I__7048 (
            .O(N__31584),
            .I(N__31535));
    Span4Mux_h I__7047 (
            .O(N__31577),
            .I(N__31535));
    LocalMux I__7046 (
            .O(N__31570),
            .I(N__31535));
    CEMux I__7045 (
            .O(N__31569),
            .I(N__31526));
    InMux I__7044 (
            .O(N__31568),
            .I(N__31526));
    InMux I__7043 (
            .O(N__31567),
            .I(N__31526));
    InMux I__7042 (
            .O(N__31566),
            .I(N__31526));
    Span4Mux_v I__7041 (
            .O(N__31559),
            .I(N__31523));
    LocalMux I__7040 (
            .O(N__31556),
            .I(N__31520));
    Span4Mux_v I__7039 (
            .O(N__31553),
            .I(N__31517));
    InMux I__7038 (
            .O(N__31552),
            .I(N__31510));
    InMux I__7037 (
            .O(N__31551),
            .I(N__31510));
    InMux I__7036 (
            .O(N__31550),
            .I(N__31510));
    InMux I__7035 (
            .O(N__31549),
            .I(N__31507));
    InMux I__7034 (
            .O(N__31548),
            .I(N__31502));
    InMux I__7033 (
            .O(N__31547),
            .I(N__31502));
    LocalMux I__7032 (
            .O(N__31542),
            .I(N__31495));
    Sp12to4 I__7031 (
            .O(N__31535),
            .I(N__31495));
    LocalMux I__7030 (
            .O(N__31526),
            .I(N__31495));
    Odrv4 I__7029 (
            .O(N__31523),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    Odrv4 I__7028 (
            .O(N__31520),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    Odrv4 I__7027 (
            .O(N__31517),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    LocalMux I__7026 (
            .O(N__31510),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    LocalMux I__7025 (
            .O(N__31507),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    LocalMux I__7024 (
            .O(N__31502),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    Odrv12 I__7023 (
            .O(N__31495),
            .I(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ));
    InMux I__7022 (
            .O(N__31480),
            .I(N__31476));
    InMux I__7021 (
            .O(N__31479),
            .I(N__31473));
    LocalMux I__7020 (
            .O(N__31476),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    LocalMux I__7019 (
            .O(N__31473),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    InMux I__7018 (
            .O(N__31468),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    InMux I__7017 (
            .O(N__31465),
            .I(N__31462));
    LocalMux I__7016 (
            .O(N__31462),
            .I(\VPP_VDDQ.count_2_1_12 ));
    InMux I__7015 (
            .O(N__31459),
            .I(N__31456));
    LocalMux I__7014 (
            .O(N__31456),
            .I(\VPP_VDDQ.count_2_1_13 ));
    InMux I__7013 (
            .O(N__31453),
            .I(N__31450));
    LocalMux I__7012 (
            .O(N__31450),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    InMux I__7011 (
            .O(N__31447),
            .I(N__31443));
    InMux I__7010 (
            .O(N__31446),
            .I(N__31440));
    LocalMux I__7009 (
            .O(N__31443),
            .I(N__31437));
    LocalMux I__7008 (
            .O(N__31440),
            .I(N__31434));
    Odrv4 I__7007 (
            .O(N__31437),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    Odrv4 I__7006 (
            .O(N__31434),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    InMux I__7005 (
            .O(N__31429),
            .I(N__31425));
    InMux I__7004 (
            .O(N__31428),
            .I(N__31422));
    LocalMux I__7003 (
            .O(N__31425),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    LocalMux I__7002 (
            .O(N__31422),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    CascadeMux I__7001 (
            .O(N__31417),
            .I(\VPP_VDDQ.count_2Z0Z_13_cascade_ ));
    InMux I__7000 (
            .O(N__31414),
            .I(N__31411));
    LocalMux I__6999 (
            .O(N__31411),
            .I(N__31407));
    InMux I__6998 (
            .O(N__31410),
            .I(N__31404));
    Sp12to4 I__6997 (
            .O(N__31407),
            .I(N__31401));
    LocalMux I__6996 (
            .O(N__31404),
            .I(N__31398));
    Odrv12 I__6995 (
            .O(N__31401),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    Odrv4 I__6994 (
            .O(N__31398),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    InMux I__6993 (
            .O(N__31393),
            .I(N__31390));
    LocalMux I__6992 (
            .O(N__31390),
            .I(\VPP_VDDQ.un9_clk_100khz_10 ));
    CascadeMux I__6991 (
            .O(N__31387),
            .I(N__31383));
    CascadeMux I__6990 (
            .O(N__31386),
            .I(N__31380));
    InMux I__6989 (
            .O(N__31383),
            .I(N__31375));
    InMux I__6988 (
            .O(N__31380),
            .I(N__31375));
    LocalMux I__6987 (
            .O(N__31375),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ));
    InMux I__6986 (
            .O(N__31372),
            .I(N__31369));
    LocalMux I__6985 (
            .O(N__31369),
            .I(\VPP_VDDQ.count_2_0_12 ));
    CascadeMux I__6984 (
            .O(N__31366),
            .I(N__31362));
    CascadeMux I__6983 (
            .O(N__31365),
            .I(N__31359));
    InMux I__6982 (
            .O(N__31362),
            .I(N__31356));
    InMux I__6981 (
            .O(N__31359),
            .I(N__31353));
    LocalMux I__6980 (
            .O(N__31356),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    LocalMux I__6979 (
            .O(N__31353),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    InMux I__6978 (
            .O(N__31348),
            .I(N__31345));
    LocalMux I__6977 (
            .O(N__31345),
            .I(\VPP_VDDQ.count_2_0_13 ));
    InMux I__6976 (
            .O(N__31342),
            .I(N__31339));
    LocalMux I__6975 (
            .O(N__31339),
            .I(N__31335));
    InMux I__6974 (
            .O(N__31338),
            .I(N__31332));
    Span4Mux_s1_h I__6973 (
            .O(N__31335),
            .I(N__31329));
    LocalMux I__6972 (
            .O(N__31332),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    Odrv4 I__6971 (
            .O(N__31329),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ));
    InMux I__6970 (
            .O(N__31324),
            .I(N__31321));
    LocalMux I__6969 (
            .O(N__31321),
            .I(N__31318));
    Odrv4 I__6968 (
            .O(N__31318),
            .I(\VPP_VDDQ.count_2_0_14 ));
    InMux I__6967 (
            .O(N__31315),
            .I(N__31312));
    LocalMux I__6966 (
            .O(N__31312),
            .I(N__31309));
    Odrv4 I__6965 (
            .O(N__31309),
            .I(\VPP_VDDQ.un9_clk_100khz_1 ));
    InMux I__6964 (
            .O(N__31306),
            .I(N__31303));
    LocalMux I__6963 (
            .O(N__31303),
            .I(\VPP_VDDQ.count_2_0_5 ));
    CascadeMux I__6962 (
            .O(N__31300),
            .I(\VPP_VDDQ.count_2_1_5_cascade_ ));
    InMux I__6961 (
            .O(N__31297),
            .I(N__31293));
    InMux I__6960 (
            .O(N__31296),
            .I(N__31290));
    LocalMux I__6959 (
            .O(N__31293),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    LocalMux I__6958 (
            .O(N__31290),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    InMux I__6957 (
            .O(N__31285),
            .I(N__31282));
    LocalMux I__6956 (
            .O(N__31282),
            .I(N__31279));
    Span4Mux_v I__6955 (
            .O(N__31279),
            .I(N__31276));
    Span4Mux_h I__6954 (
            .O(N__31276),
            .I(N__31273));
    Span4Mux_h I__6953 (
            .O(N__31273),
            .I(N__31270));
    Odrv4 I__6952 (
            .O(N__31270),
            .I(vr_ready_vccin));
    CascadeMux I__6951 (
            .O(N__31267),
            .I(N__31264));
    InMux I__6950 (
            .O(N__31264),
            .I(N__31258));
    InMux I__6949 (
            .O(N__31263),
            .I(N__31258));
    LocalMux I__6948 (
            .O(N__31258),
            .I(N__31255));
    Span4Mux_v I__6947 (
            .O(N__31255),
            .I(N__31250));
    InMux I__6946 (
            .O(N__31254),
            .I(N__31245));
    InMux I__6945 (
            .O(N__31253),
            .I(N__31245));
    Span4Mux_h I__6944 (
            .O(N__31250),
            .I(N__31240));
    LocalMux I__6943 (
            .O(N__31245),
            .I(N__31240));
    Odrv4 I__6942 (
            .O(N__31240),
            .I(\PCH_PWRGD.N_174 ));
    IoInMux I__6941 (
            .O(N__31237),
            .I(N__31233));
    InMux I__6940 (
            .O(N__31236),
            .I(N__31230));
    LocalMux I__6939 (
            .O(N__31233),
            .I(N__31227));
    LocalMux I__6938 (
            .O(N__31230),
            .I(N__31224));
    Span4Mux_s0_h I__6937 (
            .O(N__31227),
            .I(N__31221));
    Span12Mux_s3_h I__6936 (
            .O(N__31224),
            .I(N__31218));
    Span4Mux_v I__6935 (
            .O(N__31221),
            .I(N__31215));
    Odrv12 I__6934 (
            .O(N__31218),
            .I(dsw_pwrok));
    Odrv4 I__6933 (
            .O(N__31215),
            .I(dsw_pwrok));
    InMux I__6932 (
            .O(N__31210),
            .I(N__31207));
    LocalMux I__6931 (
            .O(N__31207),
            .I(N__31204));
    Span4Mux_v I__6930 (
            .O(N__31204),
            .I(N__31201));
    Odrv4 I__6929 (
            .O(N__31201),
            .I(vccst_cpu_ok));
    CascadeMux I__6928 (
            .O(N__31198),
            .I(N__31195));
    InMux I__6927 (
            .O(N__31195),
            .I(N__31192));
    LocalMux I__6926 (
            .O(N__31192),
            .I(v5s_ok));
    InMux I__6925 (
            .O(N__31189),
            .I(N__31186));
    LocalMux I__6924 (
            .O(N__31186),
            .I(N__31183));
    Span12Mux_v I__6923 (
            .O(N__31183),
            .I(N__31180));
    Odrv12 I__6922 (
            .O(N__31180),
            .I(v33s_ok));
    CascadeMux I__6921 (
            .O(N__31177),
            .I(N__31173));
    InMux I__6920 (
            .O(N__31176),
            .I(N__31168));
    InMux I__6919 (
            .O(N__31173),
            .I(N__31168));
    LocalMux I__6918 (
            .O(N__31168),
            .I(N__31160));
    CascadeMux I__6917 (
            .O(N__31167),
            .I(N__31155));
    InMux I__6916 (
            .O(N__31166),
            .I(N__31150));
    CascadeMux I__6915 (
            .O(N__31165),
            .I(N__31142));
    InMux I__6914 (
            .O(N__31164),
            .I(N__31134));
    InMux I__6913 (
            .O(N__31163),
            .I(N__31134));
    Span4Mux_s3_v I__6912 (
            .O(N__31160),
            .I(N__31129));
    InMux I__6911 (
            .O(N__31159),
            .I(N__31124));
    InMux I__6910 (
            .O(N__31158),
            .I(N__31124));
    InMux I__6909 (
            .O(N__31155),
            .I(N__31121));
    CascadeMux I__6908 (
            .O(N__31154),
            .I(N__31117));
    CascadeMux I__6907 (
            .O(N__31153),
            .I(N__31111));
    LocalMux I__6906 (
            .O(N__31150),
            .I(N__31105));
    InMux I__6905 (
            .O(N__31149),
            .I(N__31102));
    InMux I__6904 (
            .O(N__31148),
            .I(N__31099));
    InMux I__6903 (
            .O(N__31147),
            .I(N__31090));
    InMux I__6902 (
            .O(N__31146),
            .I(N__31090));
    InMux I__6901 (
            .O(N__31145),
            .I(N__31090));
    InMux I__6900 (
            .O(N__31142),
            .I(N__31090));
    InMux I__6899 (
            .O(N__31141),
            .I(N__31085));
    InMux I__6898 (
            .O(N__31140),
            .I(N__31085));
    InMux I__6897 (
            .O(N__31139),
            .I(N__31082));
    LocalMux I__6896 (
            .O(N__31134),
            .I(N__31079));
    InMux I__6895 (
            .O(N__31133),
            .I(N__31076));
    InMux I__6894 (
            .O(N__31132),
            .I(N__31073));
    Span4Mux_h I__6893 (
            .O(N__31129),
            .I(N__31068));
    LocalMux I__6892 (
            .O(N__31124),
            .I(N__31068));
    LocalMux I__6891 (
            .O(N__31121),
            .I(N__31065));
    InMux I__6890 (
            .O(N__31120),
            .I(N__31060));
    InMux I__6889 (
            .O(N__31117),
            .I(N__31060));
    InMux I__6888 (
            .O(N__31116),
            .I(N__31055));
    InMux I__6887 (
            .O(N__31115),
            .I(N__31055));
    InMux I__6886 (
            .O(N__31114),
            .I(N__31050));
    InMux I__6885 (
            .O(N__31111),
            .I(N__31050));
    InMux I__6884 (
            .O(N__31110),
            .I(N__31045));
    InMux I__6883 (
            .O(N__31109),
            .I(N__31045));
    CascadeMux I__6882 (
            .O(N__31108),
            .I(N__31042));
    Span4Mux_v I__6881 (
            .O(N__31105),
            .I(N__31039));
    LocalMux I__6880 (
            .O(N__31102),
            .I(N__31032));
    LocalMux I__6879 (
            .O(N__31099),
            .I(N__31032));
    LocalMux I__6878 (
            .O(N__31090),
            .I(N__31032));
    LocalMux I__6877 (
            .O(N__31085),
            .I(N__31029));
    LocalMux I__6876 (
            .O(N__31082),
            .I(N__31019));
    Span4Mux_h I__6875 (
            .O(N__31079),
            .I(N__31019));
    LocalMux I__6874 (
            .O(N__31076),
            .I(N__31019));
    LocalMux I__6873 (
            .O(N__31073),
            .I(N__31016));
    Span4Mux_h I__6872 (
            .O(N__31068),
            .I(N__31013));
    Span4Mux_h I__6871 (
            .O(N__31065),
            .I(N__31006));
    LocalMux I__6870 (
            .O(N__31060),
            .I(N__31006));
    LocalMux I__6869 (
            .O(N__31055),
            .I(N__31006));
    LocalMux I__6868 (
            .O(N__31050),
            .I(N__31001));
    LocalMux I__6867 (
            .O(N__31045),
            .I(N__31001));
    InMux I__6866 (
            .O(N__31042),
            .I(N__30998));
    Span4Mux_h I__6865 (
            .O(N__31039),
            .I(N__30991));
    Span4Mux_v I__6864 (
            .O(N__31032),
            .I(N__30991));
    Span4Mux_s3_h I__6863 (
            .O(N__31029),
            .I(N__30991));
    InMux I__6862 (
            .O(N__31028),
            .I(N__30984));
    InMux I__6861 (
            .O(N__31027),
            .I(N__30984));
    InMux I__6860 (
            .O(N__31026),
            .I(N__30984));
    Span4Mux_v I__6859 (
            .O(N__31019),
            .I(N__30981));
    Span4Mux_v I__6858 (
            .O(N__31016),
            .I(N__30972));
    Span4Mux_v I__6857 (
            .O(N__31013),
            .I(N__30972));
    Span4Mux_v I__6856 (
            .O(N__31006),
            .I(N__30972));
    Span4Mux_v I__6855 (
            .O(N__31001),
            .I(N__30972));
    LocalMux I__6854 (
            .O(N__30998),
            .I(slp_s3n_signal));
    Odrv4 I__6853 (
            .O(N__30991),
            .I(slp_s3n_signal));
    LocalMux I__6852 (
            .O(N__30984),
            .I(slp_s3n_signal));
    Odrv4 I__6851 (
            .O(N__30981),
            .I(slp_s3n_signal));
    Odrv4 I__6850 (
            .O(N__30972),
            .I(slp_s3n_signal));
    CascadeMux I__6849 (
            .O(N__30961),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ));
    InMux I__6848 (
            .O(N__30958),
            .I(N__30955));
    LocalMux I__6847 (
            .O(N__30955),
            .I(N__30952));
    Span4Mux_v I__6846 (
            .O(N__30952),
            .I(N__30947));
    InMux I__6845 (
            .O(N__30951),
            .I(N__30942));
    InMux I__6844 (
            .O(N__30950),
            .I(N__30942));
    Span4Mux_s0_h I__6843 (
            .O(N__30947),
            .I(N__30935));
    LocalMux I__6842 (
            .O(N__30942),
            .I(N__30932));
    InMux I__6841 (
            .O(N__30941),
            .I(N__30923));
    InMux I__6840 (
            .O(N__30940),
            .I(N__30923));
    InMux I__6839 (
            .O(N__30939),
            .I(N__30923));
    InMux I__6838 (
            .O(N__30938),
            .I(N__30923));
    Odrv4 I__6837 (
            .O(N__30935),
            .I(rsmrst_pwrgd_signal));
    Odrv12 I__6836 (
            .O(N__30932),
            .I(rsmrst_pwrgd_signal));
    LocalMux I__6835 (
            .O(N__30923),
            .I(rsmrst_pwrgd_signal));
    IoInMux I__6834 (
            .O(N__30916),
            .I(N__30913));
    LocalMux I__6833 (
            .O(N__30913),
            .I(N__30910));
    IoSpan4Mux I__6832 (
            .O(N__30910),
            .I(N__30907));
    Span4Mux_s3_v I__6831 (
            .O(N__30907),
            .I(N__30904));
    Span4Mux_v I__6830 (
            .O(N__30904),
            .I(N__30901));
    Odrv4 I__6829 (
            .O(N__30901),
            .I(vccin_en));
    InMux I__6828 (
            .O(N__30898),
            .I(N__30895));
    LocalMux I__6827 (
            .O(N__30895),
            .I(\VPP_VDDQ.un1_count_2_1_axb_6 ));
    InMux I__6826 (
            .O(N__30892),
            .I(N__30888));
    InMux I__6825 (
            .O(N__30891),
            .I(N__30885));
    LocalMux I__6824 (
            .O(N__30888),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    LocalMux I__6823 (
            .O(N__30885),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    InMux I__6822 (
            .O(N__30880),
            .I(N__30874));
    InMux I__6821 (
            .O(N__30879),
            .I(N__30874));
    LocalMux I__6820 (
            .O(N__30874),
            .I(N__30871));
    Odrv4 I__6819 (
            .O(N__30871),
            .I(\VPP_VDDQ.count_2_1_6 ));
    InMux I__6818 (
            .O(N__30868),
            .I(N__30865));
    LocalMux I__6817 (
            .O(N__30865),
            .I(\VPP_VDDQ.un9_clk_100khz_9 ));
    CascadeMux I__6816 (
            .O(N__30862),
            .I(\VPP_VDDQ.un9_clk_100khz_0_cascade_ ));
    InMux I__6815 (
            .O(N__30859),
            .I(N__30856));
    LocalMux I__6814 (
            .O(N__30856),
            .I(N__30853));
    Odrv4 I__6813 (
            .O(N__30853),
            .I(\VPP_VDDQ.un9_clk_100khz_13 ));
    CascadeMux I__6812 (
            .O(N__30850),
            .I(N__30847));
    InMux I__6811 (
            .O(N__30847),
            .I(N__30843));
    InMux I__6810 (
            .O(N__30846),
            .I(N__30840));
    LocalMux I__6809 (
            .O(N__30843),
            .I(N__30837));
    LocalMux I__6808 (
            .O(N__30840),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ));
    Odrv12 I__6807 (
            .O(N__30837),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ));
    CascadeMux I__6806 (
            .O(N__30832),
            .I(\VPP_VDDQ.N_1_i_cascade_ ));
    CascadeMux I__6805 (
            .O(N__30829),
            .I(N__30826));
    InMux I__6804 (
            .O(N__30826),
            .I(N__30820));
    InMux I__6803 (
            .O(N__30825),
            .I(N__30820));
    LocalMux I__6802 (
            .O(N__30820),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    InMux I__6801 (
            .O(N__30817),
            .I(N__30814));
    LocalMux I__6800 (
            .O(N__30814),
            .I(\VPP_VDDQ.N_361_0 ));
    CascadeMux I__6799 (
            .O(N__30811),
            .I(N__30804));
    InMux I__6798 (
            .O(N__30810),
            .I(N__30800));
    InMux I__6797 (
            .O(N__30809),
            .I(N__30797));
    InMux I__6796 (
            .O(N__30808),
            .I(N__30794));
    InMux I__6795 (
            .O(N__30807),
            .I(N__30789));
    InMux I__6794 (
            .O(N__30804),
            .I(N__30789));
    InMux I__6793 (
            .O(N__30803),
            .I(N__30786));
    LocalMux I__6792 (
            .O(N__30800),
            .I(N__30775));
    LocalMux I__6791 (
            .O(N__30797),
            .I(N__30772));
    LocalMux I__6790 (
            .O(N__30794),
            .I(N__30769));
    LocalMux I__6789 (
            .O(N__30789),
            .I(N__30766));
    LocalMux I__6788 (
            .O(N__30786),
            .I(N__30763));
    CEMux I__6787 (
            .O(N__30785),
            .I(N__30736));
    CEMux I__6786 (
            .O(N__30784),
            .I(N__30736));
    CEMux I__6785 (
            .O(N__30783),
            .I(N__30736));
    CEMux I__6784 (
            .O(N__30782),
            .I(N__30736));
    CEMux I__6783 (
            .O(N__30781),
            .I(N__30736));
    CEMux I__6782 (
            .O(N__30780),
            .I(N__30736));
    CEMux I__6781 (
            .O(N__30779),
            .I(N__30736));
    CEMux I__6780 (
            .O(N__30778),
            .I(N__30736));
    Glb2LocalMux I__6779 (
            .O(N__30775),
            .I(N__30736));
    Glb2LocalMux I__6778 (
            .O(N__30772),
            .I(N__30736));
    Glb2LocalMux I__6777 (
            .O(N__30769),
            .I(N__30736));
    Glb2LocalMux I__6776 (
            .O(N__30766),
            .I(N__30736));
    Glb2LocalMux I__6775 (
            .O(N__30763),
            .I(N__30736));
    GlobalMux I__6774 (
            .O(N__30736),
            .I(N__30733));
    gio2CtrlBuf I__6773 (
            .O(N__30733),
            .I(N_570_g));
    CascadeMux I__6772 (
            .O(N__30730),
            .I(N__30727));
    InMux I__6771 (
            .O(N__30727),
            .I(N__30721));
    InMux I__6770 (
            .O(N__30726),
            .I(N__30721));
    LocalMux I__6769 (
            .O(N__30721),
            .I(\VPP_VDDQ.N_2192_i ));
    InMux I__6768 (
            .O(N__30718),
            .I(N__30713));
    InMux I__6767 (
            .O(N__30717),
            .I(N__30708));
    InMux I__6766 (
            .O(N__30716),
            .I(N__30708));
    LocalMux I__6765 (
            .O(N__30713),
            .I(\VPP_VDDQ.N_62 ));
    LocalMux I__6764 (
            .O(N__30708),
            .I(\VPP_VDDQ.N_62 ));
    SRMux I__6763 (
            .O(N__30703),
            .I(N__30700));
    LocalMux I__6762 (
            .O(N__30700),
            .I(N__30697));
    Odrv4 I__6761 (
            .O(N__30697),
            .I(\VPP_VDDQ.N_62_i ));
    CascadeMux I__6760 (
            .O(N__30694),
            .I(\VPP_VDDQ.count_2_1_14_cascade_ ));
    CascadeMux I__6759 (
            .O(N__30691),
            .I(\VPP_VDDQ.count_2_1_4_cascade_ ));
    CascadeMux I__6758 (
            .O(N__30688),
            .I(N__30684));
    CascadeMux I__6757 (
            .O(N__30687),
            .I(N__30681));
    InMux I__6756 (
            .O(N__30684),
            .I(N__30676));
    InMux I__6755 (
            .O(N__30681),
            .I(N__30676));
    LocalMux I__6754 (
            .O(N__30676),
            .I(N__30673));
    Span4Mux_s0_h I__6753 (
            .O(N__30673),
            .I(N__30670));
    Odrv4 I__6752 (
            .O(N__30670),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ));
    InMux I__6751 (
            .O(N__30667),
            .I(N__30664));
    LocalMux I__6750 (
            .O(N__30664),
            .I(\VPP_VDDQ.count_2_0_4 ));
    CascadeMux I__6749 (
            .O(N__30661),
            .I(N__30657));
    InMux I__6748 (
            .O(N__30660),
            .I(N__30652));
    InMux I__6747 (
            .O(N__30657),
            .I(N__30652));
    LocalMux I__6746 (
            .O(N__30652),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ));
    InMux I__6745 (
            .O(N__30649),
            .I(N__30646));
    LocalMux I__6744 (
            .O(N__30646),
            .I(\VPP_VDDQ.un6_count_11 ));
    InMux I__6743 (
            .O(N__30643),
            .I(N__30640));
    LocalMux I__6742 (
            .O(N__30640),
            .I(\VPP_VDDQ.un6_count_9 ));
    IoInMux I__6741 (
            .O(N__30637),
            .I(N__30633));
    CascadeMux I__6740 (
            .O(N__30636),
            .I(N__30627));
    LocalMux I__6739 (
            .O(N__30633),
            .I(N__30624));
    CascadeMux I__6738 (
            .O(N__30632),
            .I(N__30621));
    CascadeMux I__6737 (
            .O(N__30631),
            .I(N__30617));
    InMux I__6736 (
            .O(N__30630),
            .I(N__30607));
    InMux I__6735 (
            .O(N__30627),
            .I(N__30607));
    Span4Mux_s0_h I__6734 (
            .O(N__30624),
            .I(N__30596));
    InMux I__6733 (
            .O(N__30621),
            .I(N__30589));
    InMux I__6732 (
            .O(N__30620),
            .I(N__30589));
    InMux I__6731 (
            .O(N__30617),
            .I(N__30589));
    InMux I__6730 (
            .O(N__30616),
            .I(N__30580));
    InMux I__6729 (
            .O(N__30615),
            .I(N__30580));
    InMux I__6728 (
            .O(N__30614),
            .I(N__30580));
    InMux I__6727 (
            .O(N__30613),
            .I(N__30580));
    InMux I__6726 (
            .O(N__30612),
            .I(N__30571));
    LocalMux I__6725 (
            .O(N__30607),
            .I(N__30568));
    InMux I__6724 (
            .O(N__30606),
            .I(N__30565));
    InMux I__6723 (
            .O(N__30605),
            .I(N__30558));
    InMux I__6722 (
            .O(N__30604),
            .I(N__30558));
    InMux I__6721 (
            .O(N__30603),
            .I(N__30558));
    InMux I__6720 (
            .O(N__30602),
            .I(N__30549));
    InMux I__6719 (
            .O(N__30601),
            .I(N__30549));
    InMux I__6718 (
            .O(N__30600),
            .I(N__30549));
    InMux I__6717 (
            .O(N__30599),
            .I(N__30549));
    Span4Mux_v I__6716 (
            .O(N__30596),
            .I(N__30539));
    LocalMux I__6715 (
            .O(N__30589),
            .I(N__30539));
    LocalMux I__6714 (
            .O(N__30580),
            .I(N__30539));
    InMux I__6713 (
            .O(N__30579),
            .I(N__30532));
    InMux I__6712 (
            .O(N__30578),
            .I(N__30532));
    InMux I__6711 (
            .O(N__30577),
            .I(N__30532));
    InMux I__6710 (
            .O(N__30576),
            .I(N__30526));
    InMux I__6709 (
            .O(N__30575),
            .I(N__30526));
    InMux I__6708 (
            .O(N__30574),
            .I(N__30523));
    LocalMux I__6707 (
            .O(N__30571),
            .I(N__30520));
    Span4Mux_s2_h I__6706 (
            .O(N__30568),
            .I(N__30511));
    LocalMux I__6705 (
            .O(N__30565),
            .I(N__30511));
    LocalMux I__6704 (
            .O(N__30558),
            .I(N__30511));
    LocalMux I__6703 (
            .O(N__30549),
            .I(N__30511));
    InMux I__6702 (
            .O(N__30548),
            .I(N__30508));
    InMux I__6701 (
            .O(N__30547),
            .I(N__30503));
    InMux I__6700 (
            .O(N__30546),
            .I(N__30503));
    Span4Mux_v I__6699 (
            .O(N__30539),
            .I(N__30498));
    LocalMux I__6698 (
            .O(N__30532),
            .I(N__30498));
    InMux I__6697 (
            .O(N__30531),
            .I(N__30495));
    LocalMux I__6696 (
            .O(N__30526),
            .I(N__30492));
    LocalMux I__6695 (
            .O(N__30523),
            .I(N__30485));
    Span4Mux_v I__6694 (
            .O(N__30520),
            .I(N__30485));
    Span4Mux_v I__6693 (
            .O(N__30511),
            .I(N__30482));
    LocalMux I__6692 (
            .O(N__30508),
            .I(N__30477));
    LocalMux I__6691 (
            .O(N__30503),
            .I(N__30477));
    Span4Mux_h I__6690 (
            .O(N__30498),
            .I(N__30474));
    LocalMux I__6689 (
            .O(N__30495),
            .I(N__30469));
    Span4Mux_s3_h I__6688 (
            .O(N__30492),
            .I(N__30469));
    InMux I__6687 (
            .O(N__30491),
            .I(N__30466));
    InMux I__6686 (
            .O(N__30490),
            .I(N__30462));
    Span4Mux_v I__6685 (
            .O(N__30485),
            .I(N__30457));
    Span4Mux_h I__6684 (
            .O(N__30482),
            .I(N__30457));
    Span4Mux_s2_h I__6683 (
            .O(N__30477),
            .I(N__30454));
    Span4Mux_h I__6682 (
            .O(N__30474),
            .I(N__30447));
    Span4Mux_v I__6681 (
            .O(N__30469),
            .I(N__30447));
    LocalMux I__6680 (
            .O(N__30466),
            .I(N__30447));
    InMux I__6679 (
            .O(N__30465),
            .I(N__30444));
    LocalMux I__6678 (
            .O(N__30462),
            .I(suswarn_n));
    Odrv4 I__6677 (
            .O(N__30457),
            .I(suswarn_n));
    Odrv4 I__6676 (
            .O(N__30454),
            .I(suswarn_n));
    Odrv4 I__6675 (
            .O(N__30447),
            .I(suswarn_n));
    LocalMux I__6674 (
            .O(N__30444),
            .I(suswarn_n));
    CascadeMux I__6673 (
            .O(N__30433),
            .I(\VPP_VDDQ.N_361_0_cascade_ ));
    CascadeMux I__6672 (
            .O(N__30430),
            .I(\VPP_VDDQ.N_62_cascade_ ));
    CascadeMux I__6671 (
            .O(N__30427),
            .I(\VPP_VDDQ.delayed_vddq_ok_en_cascade_ ));
    InMux I__6670 (
            .O(N__30424),
            .I(N__30421));
    LocalMux I__6669 (
            .O(N__30421),
            .I(N__30418));
    Span12Mux_s11_h I__6668 (
            .O(N__30418),
            .I(N__30415));
    Odrv12 I__6667 (
            .O(N__30415),
            .I(VPP_VDDQ_delayed_vddq_ok));
    CascadeMux I__6666 (
            .O(N__30412),
            .I(N__30407));
    CascadeMux I__6665 (
            .O(N__30411),
            .I(N__30403));
    InMux I__6664 (
            .O(N__30410),
            .I(N__30396));
    InMux I__6663 (
            .O(N__30407),
            .I(N__30389));
    InMux I__6662 (
            .O(N__30406),
            .I(N__30389));
    InMux I__6661 (
            .O(N__30403),
            .I(N__30389));
    InMux I__6660 (
            .O(N__30402),
            .I(N__30380));
    InMux I__6659 (
            .O(N__30401),
            .I(N__30380));
    InMux I__6658 (
            .O(N__30400),
            .I(N__30380));
    InMux I__6657 (
            .O(N__30399),
            .I(N__30380));
    LocalMux I__6656 (
            .O(N__30396),
            .I(N__30375));
    LocalMux I__6655 (
            .O(N__30389),
            .I(N__30375));
    LocalMux I__6654 (
            .O(N__30380),
            .I(N__30372));
    Span4Mux_v I__6653 (
            .O(N__30375),
            .I(N__30365));
    Span4Mux_v I__6652 (
            .O(N__30372),
            .I(N__30365));
    InMux I__6651 (
            .O(N__30371),
            .I(N__30360));
    InMux I__6650 (
            .O(N__30370),
            .I(N__30360));
    Span4Mux_v I__6649 (
            .O(N__30365),
            .I(N__30353));
    LocalMux I__6648 (
            .O(N__30360),
            .I(N__30353));
    InMux I__6647 (
            .O(N__30359),
            .I(N__30348));
    InMux I__6646 (
            .O(N__30358),
            .I(N__30348));
    Span4Mux_v I__6645 (
            .O(N__30353),
            .I(N__30345));
    LocalMux I__6644 (
            .O(N__30348),
            .I(N__30342));
    Odrv4 I__6643 (
            .O(N__30345),
            .I(vddq_ok));
    Odrv12 I__6642 (
            .O(N__30342),
            .I(vddq_ok));
    CascadeMux I__6641 (
            .O(N__30337),
            .I(N__30334));
    InMux I__6640 (
            .O(N__30334),
            .I(N__30331));
    LocalMux I__6639 (
            .O(N__30331),
            .I(\VPP_VDDQ.delayed_vddq_ok_en ));
    InMux I__6638 (
            .O(N__30328),
            .I(N__30322));
    InMux I__6637 (
            .O(N__30327),
            .I(N__30322));
    LocalMux I__6636 (
            .O(N__30322),
            .I(\VPP_VDDQ.delayed_vddq_okZ0 ));
    InMux I__6635 (
            .O(N__30319),
            .I(N__30316));
    LocalMux I__6634 (
            .O(N__30316),
            .I(\VPP_VDDQ.curr_state_7_0 ));
    CascadeMux I__6633 (
            .O(N__30313),
            .I(\VPP_VDDQ.curr_state_7_0_cascade_ ));
    InMux I__6632 (
            .O(N__30310),
            .I(N__30307));
    LocalMux I__6631 (
            .O(N__30307),
            .I(N__30304));
    Span4Mux_s2_v I__6630 (
            .O(N__30304),
            .I(N__30300));
    InMux I__6629 (
            .O(N__30303),
            .I(N__30297));
    Odrv4 I__6628 (
            .O(N__30300),
            .I(N_246));
    LocalMux I__6627 (
            .O(N__30297),
            .I(N_246));
    CascadeMux I__6626 (
            .O(N__30292),
            .I(N_246_cascade_));
    InMux I__6625 (
            .O(N__30289),
            .I(N__30285));
    InMux I__6624 (
            .O(N__30288),
            .I(N__30282));
    LocalMux I__6623 (
            .O(N__30285),
            .I(N_381));
    LocalMux I__6622 (
            .O(N__30282),
            .I(N_381));
    InMux I__6621 (
            .O(N__30277),
            .I(N__30266));
    InMux I__6620 (
            .O(N__30276),
            .I(N__30266));
    InMux I__6619 (
            .O(N__30275),
            .I(N__30266));
    InMux I__6618 (
            .O(N__30274),
            .I(N__30261));
    InMux I__6617 (
            .O(N__30273),
            .I(N__30261));
    LocalMux I__6616 (
            .O(N__30266),
            .I(N__30257));
    LocalMux I__6615 (
            .O(N__30261),
            .I(N__30254));
    InMux I__6614 (
            .O(N__30260),
            .I(N__30251));
    Span4Mux_s2_h I__6613 (
            .O(N__30257),
            .I(N__30248));
    Span12Mux_s3_h I__6612 (
            .O(N__30254),
            .I(N__30245));
    LocalMux I__6611 (
            .O(N__30251),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    Odrv4 I__6610 (
            .O(N__30248),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    Odrv12 I__6609 (
            .O(N__30245),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    InMux I__6608 (
            .O(N__30238),
            .I(N__30234));
    CascadeMux I__6607 (
            .O(N__30237),
            .I(N__30230));
    LocalMux I__6606 (
            .O(N__30234),
            .I(N__30225));
    InMux I__6605 (
            .O(N__30233),
            .I(N__30222));
    InMux I__6604 (
            .O(N__30230),
            .I(N__30219));
    CascadeMux I__6603 (
            .O(N__30229),
            .I(N__30215));
    InMux I__6602 (
            .O(N__30228),
            .I(N__30209));
    Span4Mux_h I__6601 (
            .O(N__30225),
            .I(N__30206));
    LocalMux I__6600 (
            .O(N__30222),
            .I(N__30201));
    LocalMux I__6599 (
            .O(N__30219),
            .I(N__30201));
    InMux I__6598 (
            .O(N__30218),
            .I(N__30194));
    InMux I__6597 (
            .O(N__30215),
            .I(N__30194));
    InMux I__6596 (
            .O(N__30214),
            .I(N__30194));
    InMux I__6595 (
            .O(N__30213),
            .I(N__30191));
    IoInMux I__6594 (
            .O(N__30212),
            .I(N__30185));
    LocalMux I__6593 (
            .O(N__30209),
            .I(N__30178));
    Span4Mux_h I__6592 (
            .O(N__30206),
            .I(N__30178));
    Span4Mux_v I__6591 (
            .O(N__30201),
            .I(N__30178));
    LocalMux I__6590 (
            .O(N__30194),
            .I(N__30175));
    LocalMux I__6589 (
            .O(N__30191),
            .I(N__30172));
    InMux I__6588 (
            .O(N__30190),
            .I(N__30169));
    InMux I__6587 (
            .O(N__30189),
            .I(N__30166));
    CascadeMux I__6586 (
            .O(N__30188),
            .I(N__30161));
    LocalMux I__6585 (
            .O(N__30185),
            .I(N__30156));
    Span4Mux_v I__6584 (
            .O(N__30178),
            .I(N__30153));
    Span4Mux_s2_h I__6583 (
            .O(N__30175),
            .I(N__30150));
    Span4Mux_v I__6582 (
            .O(N__30172),
            .I(N__30144));
    LocalMux I__6581 (
            .O(N__30169),
            .I(N__30144));
    LocalMux I__6580 (
            .O(N__30166),
            .I(N__30141));
    InMux I__6579 (
            .O(N__30165),
            .I(N__30136));
    InMux I__6578 (
            .O(N__30164),
            .I(N__30136));
    InMux I__6577 (
            .O(N__30161),
            .I(N__30129));
    InMux I__6576 (
            .O(N__30160),
            .I(N__30129));
    InMux I__6575 (
            .O(N__30159),
            .I(N__30129));
    Span12Mux_s8_h I__6574 (
            .O(N__30156),
            .I(N__30126));
    Span4Mux_s0_h I__6573 (
            .O(N__30153),
            .I(N__30123));
    Span4Mux_v I__6572 (
            .O(N__30150),
            .I(N__30120));
    InMux I__6571 (
            .O(N__30149),
            .I(N__30117));
    Span4Mux_h I__6570 (
            .O(N__30144),
            .I(N__30108));
    Span4Mux_v I__6569 (
            .O(N__30141),
            .I(N__30108));
    LocalMux I__6568 (
            .O(N__30136),
            .I(N__30108));
    LocalMux I__6567 (
            .O(N__30129),
            .I(N__30108));
    Odrv12 I__6566 (
            .O(N__30126),
            .I(vccst_en));
    Odrv4 I__6565 (
            .O(N__30123),
            .I(vccst_en));
    Odrv4 I__6564 (
            .O(N__30120),
            .I(vccst_en));
    LocalMux I__6563 (
            .O(N__30117),
            .I(vccst_en));
    Odrv4 I__6562 (
            .O(N__30108),
            .I(vccst_en));
    InMux I__6561 (
            .O(N__30097),
            .I(N__30089));
    InMux I__6560 (
            .O(N__30096),
            .I(N__30089));
    InMux I__6559 (
            .O(N__30095),
            .I(N__30084));
    InMux I__6558 (
            .O(N__30094),
            .I(N__30084));
    LocalMux I__6557 (
            .O(N__30089),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__6556 (
            .O(N__30084),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    CascadeMux I__6555 (
            .O(N__30079),
            .I(\VPP_VDDQ.un6_count_10_cascade_ ));
    InMux I__6554 (
            .O(N__30076),
            .I(N__30073));
    LocalMux I__6553 (
            .O(N__30073),
            .I(N__30069));
    InMux I__6552 (
            .O(N__30072),
            .I(N__30066));
    Odrv4 I__6551 (
            .O(N__30069),
            .I(VPP_VDDQ_un6_count));
    LocalMux I__6550 (
            .O(N__30066),
            .I(VPP_VDDQ_un6_count));
    InMux I__6549 (
            .O(N__30061),
            .I(N__30058));
    LocalMux I__6548 (
            .O(N__30058),
            .I(\VPP_VDDQ.un6_count_8 ));
    InMux I__6547 (
            .O(N__30055),
            .I(N__30052));
    LocalMux I__6546 (
            .O(N__30052),
            .I(N__30045));
    InMux I__6545 (
            .O(N__30051),
            .I(N__30042));
    InMux I__6544 (
            .O(N__30050),
            .I(N__30039));
    InMux I__6543 (
            .O(N__30049),
            .I(N__30032));
    InMux I__6542 (
            .O(N__30048),
            .I(N__30032));
    Span4Mux_v I__6541 (
            .O(N__30045),
            .I(N__30027));
    LocalMux I__6540 (
            .O(N__30042),
            .I(N__30027));
    LocalMux I__6539 (
            .O(N__30039),
            .I(N__30024));
    InMux I__6538 (
            .O(N__30038),
            .I(N__30021));
    InMux I__6537 (
            .O(N__30037),
            .I(N__30018));
    LocalMux I__6536 (
            .O(N__30032),
            .I(N__30013));
    Span4Mux_h I__6535 (
            .O(N__30027),
            .I(N__30013));
    Odrv4 I__6534 (
            .O(N__30024),
            .I(\POWERLED.N_396 ));
    LocalMux I__6533 (
            .O(N__30021),
            .I(\POWERLED.N_396 ));
    LocalMux I__6532 (
            .O(N__30018),
            .I(\POWERLED.N_396 ));
    Odrv4 I__6531 (
            .O(N__30013),
            .I(\POWERLED.N_396 ));
    InMux I__6530 (
            .O(N__30004),
            .I(N__29999));
    InMux I__6529 (
            .O(N__30003),
            .I(N__29996));
    InMux I__6528 (
            .O(N__30002),
            .I(N__29978));
    LocalMux I__6527 (
            .O(N__29999),
            .I(N__29973));
    LocalMux I__6526 (
            .O(N__29996),
            .I(N__29973));
    InMux I__6525 (
            .O(N__29995),
            .I(N__29970));
    InMux I__6524 (
            .O(N__29994),
            .I(N__29967));
    InMux I__6523 (
            .O(N__29993),
            .I(N__29958));
    InMux I__6522 (
            .O(N__29992),
            .I(N__29958));
    InMux I__6521 (
            .O(N__29991),
            .I(N__29958));
    InMux I__6520 (
            .O(N__29990),
            .I(N__29958));
    InMux I__6519 (
            .O(N__29989),
            .I(N__29953));
    InMux I__6518 (
            .O(N__29988),
            .I(N__29953));
    InMux I__6517 (
            .O(N__29987),
            .I(N__29948));
    InMux I__6516 (
            .O(N__29986),
            .I(N__29948));
    InMux I__6515 (
            .O(N__29985),
            .I(N__29945));
    InMux I__6514 (
            .O(N__29984),
            .I(N__29940));
    InMux I__6513 (
            .O(N__29983),
            .I(N__29936));
    InMux I__6512 (
            .O(N__29982),
            .I(N__29931));
    InMux I__6511 (
            .O(N__29981),
            .I(N__29931));
    LocalMux I__6510 (
            .O(N__29978),
            .I(N__29928));
    Span4Mux_h I__6509 (
            .O(N__29973),
            .I(N__29923));
    LocalMux I__6508 (
            .O(N__29970),
            .I(N__29923));
    LocalMux I__6507 (
            .O(N__29967),
            .I(N__29918));
    LocalMux I__6506 (
            .O(N__29958),
            .I(N__29918));
    LocalMux I__6505 (
            .O(N__29953),
            .I(N__29908));
    LocalMux I__6504 (
            .O(N__29948),
            .I(N__29908));
    LocalMux I__6503 (
            .O(N__29945),
            .I(N__29905));
    InMux I__6502 (
            .O(N__29944),
            .I(N__29900));
    InMux I__6501 (
            .O(N__29943),
            .I(N__29900));
    LocalMux I__6500 (
            .O(N__29940),
            .I(N__29897));
    InMux I__6499 (
            .O(N__29939),
            .I(N__29893));
    LocalMux I__6498 (
            .O(N__29936),
            .I(N__29890));
    LocalMux I__6497 (
            .O(N__29931),
            .I(N__29887));
    Span4Mux_v I__6496 (
            .O(N__29928),
            .I(N__29880));
    Span4Mux_v I__6495 (
            .O(N__29923),
            .I(N__29880));
    Span4Mux_v I__6494 (
            .O(N__29918),
            .I(N__29880));
    InMux I__6493 (
            .O(N__29917),
            .I(N__29875));
    InMux I__6492 (
            .O(N__29916),
            .I(N__29875));
    InMux I__6491 (
            .O(N__29915),
            .I(N__29872));
    InMux I__6490 (
            .O(N__29914),
            .I(N__29867));
    InMux I__6489 (
            .O(N__29913),
            .I(N__29867));
    Span4Mux_h I__6488 (
            .O(N__29908),
            .I(N__29864));
    Span4Mux_v I__6487 (
            .O(N__29905),
            .I(N__29857));
    LocalMux I__6486 (
            .O(N__29900),
            .I(N__29857));
    Span4Mux_h I__6485 (
            .O(N__29897),
            .I(N__29857));
    InMux I__6484 (
            .O(N__29896),
            .I(N__29854));
    LocalMux I__6483 (
            .O(N__29893),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    Odrv4 I__6482 (
            .O(N__29890),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    Odrv12 I__6481 (
            .O(N__29887),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    Odrv4 I__6480 (
            .O(N__29880),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    LocalMux I__6479 (
            .O(N__29875),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    LocalMux I__6478 (
            .O(N__29872),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    LocalMux I__6477 (
            .O(N__29867),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    Odrv4 I__6476 (
            .O(N__29864),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    Odrv4 I__6475 (
            .O(N__29857),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    LocalMux I__6474 (
            .O(N__29854),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ));
    CascadeMux I__6473 (
            .O(N__29833),
            .I(\POWERLED.count_clk_en_2_cascade_ ));
    CascadeMux I__6472 (
            .O(N__29830),
            .I(N__29822));
    CascadeMux I__6471 (
            .O(N__29829),
            .I(N__29817));
    CascadeMux I__6470 (
            .O(N__29828),
            .I(N__29813));
    InMux I__6469 (
            .O(N__29827),
            .I(N__29803));
    IoInMux I__6468 (
            .O(N__29826),
            .I(N__29800));
    InMux I__6467 (
            .O(N__29825),
            .I(N__29797));
    InMux I__6466 (
            .O(N__29822),
            .I(N__29790));
    InMux I__6465 (
            .O(N__29821),
            .I(N__29790));
    InMux I__6464 (
            .O(N__29820),
            .I(N__29790));
    InMux I__6463 (
            .O(N__29817),
            .I(N__29781));
    InMux I__6462 (
            .O(N__29816),
            .I(N__29781));
    InMux I__6461 (
            .O(N__29813),
            .I(N__29781));
    InMux I__6460 (
            .O(N__29812),
            .I(N__29781));
    CascadeMux I__6459 (
            .O(N__29811),
            .I(N__29775));
    InMux I__6458 (
            .O(N__29810),
            .I(N__29763));
    InMux I__6457 (
            .O(N__29809),
            .I(N__29763));
    InMux I__6456 (
            .O(N__29808),
            .I(N__29763));
    InMux I__6455 (
            .O(N__29807),
            .I(N__29763));
    CascadeMux I__6454 (
            .O(N__29806),
            .I(N__29760));
    LocalMux I__6453 (
            .O(N__29803),
            .I(N__29755));
    LocalMux I__6452 (
            .O(N__29800),
            .I(N__29752));
    LocalMux I__6451 (
            .O(N__29797),
            .I(N__29745));
    LocalMux I__6450 (
            .O(N__29790),
            .I(N__29745));
    LocalMux I__6449 (
            .O(N__29781),
            .I(N__29745));
    InMux I__6448 (
            .O(N__29780),
            .I(N__29738));
    InMux I__6447 (
            .O(N__29779),
            .I(N__29738));
    InMux I__6446 (
            .O(N__29778),
            .I(N__29735));
    InMux I__6445 (
            .O(N__29775),
            .I(N__29728));
    InMux I__6444 (
            .O(N__29774),
            .I(N__29728));
    InMux I__6443 (
            .O(N__29773),
            .I(N__29728));
    InMux I__6442 (
            .O(N__29772),
            .I(N__29725));
    LocalMux I__6441 (
            .O(N__29763),
            .I(N__29722));
    InMux I__6440 (
            .O(N__29760),
            .I(N__29717));
    InMux I__6439 (
            .O(N__29759),
            .I(N__29717));
    InMux I__6438 (
            .O(N__29758),
            .I(N__29714));
    Span4Mux_v I__6437 (
            .O(N__29755),
            .I(N__29708));
    Span4Mux_s3_h I__6436 (
            .O(N__29752),
            .I(N__29705));
    Span4Mux_v I__6435 (
            .O(N__29745),
            .I(N__29702));
    InMux I__6434 (
            .O(N__29744),
            .I(N__29697));
    InMux I__6433 (
            .O(N__29743),
            .I(N__29697));
    LocalMux I__6432 (
            .O(N__29738),
            .I(N__29694));
    LocalMux I__6431 (
            .O(N__29735),
            .I(N__29689));
    LocalMux I__6430 (
            .O(N__29728),
            .I(N__29689));
    LocalMux I__6429 (
            .O(N__29725),
            .I(N__29682));
    Span4Mux_h I__6428 (
            .O(N__29722),
            .I(N__29682));
    LocalMux I__6427 (
            .O(N__29717),
            .I(N__29682));
    LocalMux I__6426 (
            .O(N__29714),
            .I(N__29679));
    InMux I__6425 (
            .O(N__29713),
            .I(N__29675));
    InMux I__6424 (
            .O(N__29712),
            .I(N__29672));
    InMux I__6423 (
            .O(N__29711),
            .I(N__29669));
    Span4Mux_v I__6422 (
            .O(N__29708),
            .I(N__29664));
    Span4Mux_h I__6421 (
            .O(N__29705),
            .I(N__29664));
    Span4Mux_v I__6420 (
            .O(N__29702),
            .I(N__29661));
    LocalMux I__6419 (
            .O(N__29697),
            .I(N__29658));
    Span4Mux_v I__6418 (
            .O(N__29694),
            .I(N__29649));
    Span4Mux_h I__6417 (
            .O(N__29689),
            .I(N__29649));
    Span4Mux_v I__6416 (
            .O(N__29682),
            .I(N__29649));
    Span4Mux_h I__6415 (
            .O(N__29679),
            .I(N__29649));
    InMux I__6414 (
            .O(N__29678),
            .I(N__29646));
    LocalMux I__6413 (
            .O(N__29675),
            .I(N__29643));
    LocalMux I__6412 (
            .O(N__29672),
            .I(G_155));
    LocalMux I__6411 (
            .O(N__29669),
            .I(G_155));
    Odrv4 I__6410 (
            .O(N__29664),
            .I(G_155));
    Odrv4 I__6409 (
            .O(N__29661),
            .I(G_155));
    Odrv4 I__6408 (
            .O(N__29658),
            .I(G_155));
    Odrv4 I__6407 (
            .O(N__29649),
            .I(G_155));
    LocalMux I__6406 (
            .O(N__29646),
            .I(G_155));
    Odrv12 I__6405 (
            .O(N__29643),
            .I(G_155));
    InMux I__6404 (
            .O(N__29626),
            .I(N__29622));
    InMux I__6403 (
            .O(N__29625),
            .I(N__29617));
    LocalMux I__6402 (
            .O(N__29622),
            .I(N__29614));
    InMux I__6401 (
            .O(N__29621),
            .I(N__29611));
    InMux I__6400 (
            .O(N__29620),
            .I(N__29608));
    LocalMux I__6399 (
            .O(N__29617),
            .I(N__29605));
    Span4Mux_h I__6398 (
            .O(N__29614),
            .I(N__29602));
    LocalMux I__6397 (
            .O(N__29611),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    LocalMux I__6396 (
            .O(N__29608),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    Odrv4 I__6395 (
            .O(N__29605),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    Odrv4 I__6394 (
            .O(N__29602),
            .I(\POWERLED.func_state_RNI_2Z0Z_1 ));
    CascadeMux I__6393 (
            .O(N__29593),
            .I(N__29584));
    InMux I__6392 (
            .O(N__29592),
            .I(N__29575));
    InMux I__6391 (
            .O(N__29591),
            .I(N__29575));
    InMux I__6390 (
            .O(N__29590),
            .I(N__29575));
    InMux I__6389 (
            .O(N__29589),
            .I(N__29570));
    InMux I__6388 (
            .O(N__29588),
            .I(N__29567));
    InMux I__6387 (
            .O(N__29587),
            .I(N__29564));
    InMux I__6386 (
            .O(N__29584),
            .I(N__29557));
    InMux I__6385 (
            .O(N__29583),
            .I(N__29557));
    InMux I__6384 (
            .O(N__29582),
            .I(N__29557));
    LocalMux I__6383 (
            .O(N__29575),
            .I(N__29554));
    CascadeMux I__6382 (
            .O(N__29574),
            .I(N__29551));
    CascadeMux I__6381 (
            .O(N__29573),
            .I(N__29548));
    LocalMux I__6380 (
            .O(N__29570),
            .I(N__29545));
    LocalMux I__6379 (
            .O(N__29567),
            .I(N__29536));
    LocalMux I__6378 (
            .O(N__29564),
            .I(N__29536));
    LocalMux I__6377 (
            .O(N__29557),
            .I(N__29536));
    Span4Mux_s3_h I__6376 (
            .O(N__29554),
            .I(N__29536));
    InMux I__6375 (
            .O(N__29551),
            .I(N__29533));
    InMux I__6374 (
            .O(N__29548),
            .I(N__29530));
    Span4Mux_v I__6373 (
            .O(N__29545),
            .I(N__29525));
    Span4Mux_v I__6372 (
            .O(N__29536),
            .I(N__29525));
    LocalMux I__6371 (
            .O(N__29533),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    LocalMux I__6370 (
            .O(N__29530),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__6369 (
            .O(N__29525),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    InMux I__6368 (
            .O(N__29518),
            .I(N__29515));
    LocalMux I__6367 (
            .O(N__29515),
            .I(\POWERLED.N_176 ));
    CascadeMux I__6366 (
            .O(N__29512),
            .I(\POWERLED.N_176_cascade_ ));
    InMux I__6365 (
            .O(N__29509),
            .I(N__29506));
    LocalMux I__6364 (
            .O(N__29506),
            .I(N__29501));
    InMux I__6363 (
            .O(N__29505),
            .I(N__29496));
    InMux I__6362 (
            .O(N__29504),
            .I(N__29496));
    Span4Mux_v I__6361 (
            .O(N__29501),
            .I(N__29491));
    LocalMux I__6360 (
            .O(N__29496),
            .I(N__29491));
    Odrv4 I__6359 (
            .O(N__29491),
            .I(\POWERLED.N_2218_i ));
    InMux I__6358 (
            .O(N__29488),
            .I(N__29485));
    LocalMux I__6357 (
            .O(N__29485),
            .I(N__29482));
    Span4Mux_v I__6356 (
            .O(N__29482),
            .I(N__29475));
    CascadeMux I__6355 (
            .O(N__29481),
            .I(N__29470));
    InMux I__6354 (
            .O(N__29480),
            .I(N__29466));
    InMux I__6353 (
            .O(N__29479),
            .I(N__29461));
    InMux I__6352 (
            .O(N__29478),
            .I(N__29461));
    IoSpan4Mux I__6351 (
            .O(N__29475),
            .I(N__29455));
    InMux I__6350 (
            .O(N__29474),
            .I(N__29452));
    CascadeMux I__6349 (
            .O(N__29473),
            .I(N__29448));
    InMux I__6348 (
            .O(N__29470),
            .I(N__29442));
    InMux I__6347 (
            .O(N__29469),
            .I(N__29442));
    LocalMux I__6346 (
            .O(N__29466),
            .I(N__29439));
    LocalMux I__6345 (
            .O(N__29461),
            .I(N__29436));
    InMux I__6344 (
            .O(N__29460),
            .I(N__29433));
    InMux I__6343 (
            .O(N__29459),
            .I(N__29430));
    InMux I__6342 (
            .O(N__29458),
            .I(N__29427));
    Span4Mux_s3_h I__6341 (
            .O(N__29455),
            .I(N__29419));
    LocalMux I__6340 (
            .O(N__29452),
            .I(N__29419));
    InMux I__6339 (
            .O(N__29451),
            .I(N__29412));
    InMux I__6338 (
            .O(N__29448),
            .I(N__29412));
    InMux I__6337 (
            .O(N__29447),
            .I(N__29412));
    LocalMux I__6336 (
            .O(N__29442),
            .I(N__29409));
    Span4Mux_h I__6335 (
            .O(N__29439),
            .I(N__29398));
    Span4Mux_s3_v I__6334 (
            .O(N__29436),
            .I(N__29398));
    LocalMux I__6333 (
            .O(N__29433),
            .I(N__29398));
    LocalMux I__6332 (
            .O(N__29430),
            .I(N__29398));
    LocalMux I__6331 (
            .O(N__29427),
            .I(N__29398));
    InMux I__6330 (
            .O(N__29426),
            .I(N__29393));
    InMux I__6329 (
            .O(N__29425),
            .I(N__29393));
    InMux I__6328 (
            .O(N__29424),
            .I(N__29389));
    Span4Mux_h I__6327 (
            .O(N__29419),
            .I(N__29384));
    LocalMux I__6326 (
            .O(N__29412),
            .I(N__29384));
    Span4Mux_v I__6325 (
            .O(N__29409),
            .I(N__29375));
    Span4Mux_v I__6324 (
            .O(N__29398),
            .I(N__29375));
    LocalMux I__6323 (
            .O(N__29393),
            .I(N__29375));
    CascadeMux I__6322 (
            .O(N__29392),
            .I(N__29372));
    LocalMux I__6321 (
            .O(N__29389),
            .I(N__29366));
    Span4Mux_v I__6320 (
            .O(N__29384),
            .I(N__29366));
    InMux I__6319 (
            .O(N__29383),
            .I(N__29361));
    InMux I__6318 (
            .O(N__29382),
            .I(N__29361));
    Sp12to4 I__6317 (
            .O(N__29375),
            .I(N__29358));
    InMux I__6316 (
            .O(N__29372),
            .I(N__29353));
    InMux I__6315 (
            .O(N__29371),
            .I(N__29353));
    Odrv4 I__6314 (
            .O(N__29366),
            .I(\POWERLED.N_2216_i ));
    LocalMux I__6313 (
            .O(N__29361),
            .I(\POWERLED.N_2216_i ));
    Odrv12 I__6312 (
            .O(N__29358),
            .I(\POWERLED.N_2216_i ));
    LocalMux I__6311 (
            .O(N__29353),
            .I(\POWERLED.N_2216_i ));
    InMux I__6310 (
            .O(N__29344),
            .I(N__29341));
    LocalMux I__6309 (
            .O(N__29341),
            .I(N__29338));
    Odrv4 I__6308 (
            .O(N__29338),
            .I(\POWERLED.N_27 ));
    CascadeMux I__6307 (
            .O(N__29335),
            .I(N__29326));
    CascadeMux I__6306 (
            .O(N__29334),
            .I(N__29323));
    InMux I__6305 (
            .O(N__29333),
            .I(N__29319));
    InMux I__6304 (
            .O(N__29332),
            .I(N__29308));
    InMux I__6303 (
            .O(N__29331),
            .I(N__29308));
    CascadeMux I__6302 (
            .O(N__29330),
            .I(N__29298));
    CascadeMux I__6301 (
            .O(N__29329),
            .I(N__29295));
    InMux I__6300 (
            .O(N__29326),
            .I(N__29291));
    InMux I__6299 (
            .O(N__29323),
            .I(N__29288));
    InMux I__6298 (
            .O(N__29322),
            .I(N__29285));
    LocalMux I__6297 (
            .O(N__29319),
            .I(N__29282));
    InMux I__6296 (
            .O(N__29318),
            .I(N__29279));
    InMux I__6295 (
            .O(N__29317),
            .I(N__29272));
    InMux I__6294 (
            .O(N__29316),
            .I(N__29272));
    InMux I__6293 (
            .O(N__29315),
            .I(N__29272));
    InMux I__6292 (
            .O(N__29314),
            .I(N__29269));
    InMux I__6291 (
            .O(N__29313),
            .I(N__29266));
    LocalMux I__6290 (
            .O(N__29308),
            .I(N__29263));
    InMux I__6289 (
            .O(N__29307),
            .I(N__29256));
    InMux I__6288 (
            .O(N__29306),
            .I(N__29256));
    InMux I__6287 (
            .O(N__29305),
            .I(N__29256));
    InMux I__6286 (
            .O(N__29304),
            .I(N__29253));
    InMux I__6285 (
            .O(N__29303),
            .I(N__29250));
    InMux I__6284 (
            .O(N__29302),
            .I(N__29247));
    InMux I__6283 (
            .O(N__29301),
            .I(N__29241));
    InMux I__6282 (
            .O(N__29298),
            .I(N__29241));
    InMux I__6281 (
            .O(N__29295),
            .I(N__29236));
    InMux I__6280 (
            .O(N__29294),
            .I(N__29236));
    LocalMux I__6279 (
            .O(N__29291),
            .I(N__29229));
    LocalMux I__6278 (
            .O(N__29288),
            .I(N__29229));
    LocalMux I__6277 (
            .O(N__29285),
            .I(N__29229));
    Span4Mux_v I__6276 (
            .O(N__29282),
            .I(N__29224));
    LocalMux I__6275 (
            .O(N__29279),
            .I(N__29224));
    LocalMux I__6274 (
            .O(N__29272),
            .I(N__29220));
    LocalMux I__6273 (
            .O(N__29269),
            .I(N__29215));
    LocalMux I__6272 (
            .O(N__29266),
            .I(N__29215));
    Span4Mux_h I__6271 (
            .O(N__29263),
            .I(N__29210));
    LocalMux I__6270 (
            .O(N__29256),
            .I(N__29210));
    LocalMux I__6269 (
            .O(N__29253),
            .I(N__29203));
    LocalMux I__6268 (
            .O(N__29250),
            .I(N__29203));
    LocalMux I__6267 (
            .O(N__29247),
            .I(N__29203));
    InMux I__6266 (
            .O(N__29246),
            .I(N__29199));
    LocalMux I__6265 (
            .O(N__29241),
            .I(N__29196));
    LocalMux I__6264 (
            .O(N__29236),
            .I(N__29193));
    Span4Mux_v I__6263 (
            .O(N__29229),
            .I(N__29188));
    Span4Mux_h I__6262 (
            .O(N__29224),
            .I(N__29188));
    InMux I__6261 (
            .O(N__29223),
            .I(N__29185));
    Span4Mux_h I__6260 (
            .O(N__29220),
            .I(N__29176));
    Span4Mux_v I__6259 (
            .O(N__29215),
            .I(N__29176));
    Span4Mux_v I__6258 (
            .O(N__29210),
            .I(N__29176));
    Span4Mux_v I__6257 (
            .O(N__29203),
            .I(N__29176));
    InMux I__6256 (
            .O(N__29202),
            .I(N__29173));
    LocalMux I__6255 (
            .O(N__29199),
            .I(N__29166));
    Span4Mux_h I__6254 (
            .O(N__29196),
            .I(N__29166));
    Span4Mux_s2_h I__6253 (
            .O(N__29193),
            .I(N__29166));
    Odrv4 I__6252 (
            .O(N__29188),
            .I(\POWERLED.func_state ));
    LocalMux I__6251 (
            .O(N__29185),
            .I(\POWERLED.func_state ));
    Odrv4 I__6250 (
            .O(N__29176),
            .I(\POWERLED.func_state ));
    LocalMux I__6249 (
            .O(N__29173),
            .I(\POWERLED.func_state ));
    Odrv4 I__6248 (
            .O(N__29166),
            .I(\POWERLED.func_state ));
    InMux I__6247 (
            .O(N__29155),
            .I(N__29152));
    LocalMux I__6246 (
            .O(N__29152),
            .I(N__29149));
    Span4Mux_s1_h I__6245 (
            .O(N__29149),
            .I(N__29146));
    Odrv4 I__6244 (
            .O(N__29146),
            .I(\POWERLED.N_219 ));
    IoInMux I__6243 (
            .O(N__29143),
            .I(N__29140));
    LocalMux I__6242 (
            .O(N__29140),
            .I(N__29137));
    Odrv4 I__6241 (
            .O(N__29137),
            .I(vpp_en));
    CascadeMux I__6240 (
            .O(N__29134),
            .I(\VPP_VDDQ.N_64_cascade_ ));
    CascadeMux I__6239 (
            .O(N__29131),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ));
    InMux I__6238 (
            .O(N__29128),
            .I(N__29122));
    InMux I__6237 (
            .O(N__29127),
            .I(N__29122));
    LocalMux I__6236 (
            .O(N__29122),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    CascadeMux I__6235 (
            .O(N__29119),
            .I(\POWERLED.count_clk_RNIZ0Z_1_cascade_ ));
    InMux I__6234 (
            .O(N__29116),
            .I(N__29110));
    InMux I__6233 (
            .O(N__29115),
            .I(N__29110));
    LocalMux I__6232 (
            .O(N__29110),
            .I(N__29106));
    InMux I__6231 (
            .O(N__29109),
            .I(N__29103));
    Span4Mux_h I__6230 (
            .O(N__29106),
            .I(N__29100));
    LocalMux I__6229 (
            .O(N__29103),
            .I(\POWERLED.count_clk_RNI_0Z0Z_1 ));
    Odrv4 I__6228 (
            .O(N__29100),
            .I(\POWERLED.count_clk_RNI_0Z0Z_1 ));
    CascadeMux I__6227 (
            .O(N__29095),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_a2_0_0_cascade_ ));
    InMux I__6226 (
            .O(N__29092),
            .I(N__29089));
    LocalMux I__6225 (
            .O(N__29089),
            .I(N__29086));
    Span4Mux_s1_h I__6224 (
            .O(N__29086),
            .I(N__29083));
    Span4Mux_v I__6223 (
            .O(N__29083),
            .I(N__29080));
    Odrv4 I__6222 (
            .O(N__29080),
            .I(\POWERLED.N_285 ));
    InMux I__6221 (
            .O(N__29077),
            .I(N__29074));
    LocalMux I__6220 (
            .O(N__29074),
            .I(\POWERLED.N_177 ));
    CascadeMux I__6219 (
            .O(N__29071),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_1_cascade_ ));
    CascadeMux I__6218 (
            .O(N__29068),
            .I(N__29063));
    InMux I__6217 (
            .O(N__29067),
            .I(N__29055));
    InMux I__6216 (
            .O(N__29066),
            .I(N__29055));
    InMux I__6215 (
            .O(N__29063),
            .I(N__29052));
    InMux I__6214 (
            .O(N__29062),
            .I(N__29044));
    InMux I__6213 (
            .O(N__29061),
            .I(N__29044));
    InMux I__6212 (
            .O(N__29060),
            .I(N__29041));
    LocalMux I__6211 (
            .O(N__29055),
            .I(N__29037));
    LocalMux I__6210 (
            .O(N__29052),
            .I(N__29034));
    InMux I__6209 (
            .O(N__29051),
            .I(N__29031));
    InMux I__6208 (
            .O(N__29050),
            .I(N__29026));
    InMux I__6207 (
            .O(N__29049),
            .I(N__29026));
    LocalMux I__6206 (
            .O(N__29044),
            .I(N__29021));
    LocalMux I__6205 (
            .O(N__29041),
            .I(N__29021));
    InMux I__6204 (
            .O(N__29040),
            .I(N__29018));
    Span4Mux_v I__6203 (
            .O(N__29037),
            .I(N__29011));
    Span4Mux_h I__6202 (
            .O(N__29034),
            .I(N__29011));
    LocalMux I__6201 (
            .O(N__29031),
            .I(N__29011));
    LocalMux I__6200 (
            .O(N__29026),
            .I(N__29008));
    Span4Mux_v I__6199 (
            .O(N__29021),
            .I(N__29003));
    LocalMux I__6198 (
            .O(N__29018),
            .I(N__29003));
    Span4Mux_v I__6197 (
            .O(N__29011),
            .I(N__29000));
    Span4Mux_v I__6196 (
            .O(N__29008),
            .I(N__28995));
    Span4Mux_h I__6195 (
            .O(N__29003),
            .I(N__28995));
    Span4Mux_v I__6194 (
            .O(N__29000),
            .I(N__28992));
    Span4Mux_v I__6193 (
            .O(N__28995),
            .I(N__28989));
    Odrv4 I__6192 (
            .O(N__28992),
            .I(gpio_fpga_soc_4));
    Odrv4 I__6191 (
            .O(N__28989),
            .I(gpio_fpga_soc_4));
    InMux I__6190 (
            .O(N__28984),
            .I(N__28974));
    InMux I__6189 (
            .O(N__28983),
            .I(N__28974));
    InMux I__6188 (
            .O(N__28982),
            .I(N__28971));
    InMux I__6187 (
            .O(N__28981),
            .I(N__28966));
    InMux I__6186 (
            .O(N__28980),
            .I(N__28966));
    InMux I__6185 (
            .O(N__28979),
            .I(N__28963));
    LocalMux I__6184 (
            .O(N__28974),
            .I(N__28950));
    LocalMux I__6183 (
            .O(N__28971),
            .I(N__28950));
    LocalMux I__6182 (
            .O(N__28966),
            .I(N__28945));
    LocalMux I__6181 (
            .O(N__28963),
            .I(N__28945));
    InMux I__6180 (
            .O(N__28962),
            .I(N__28942));
    InMux I__6179 (
            .O(N__28961),
            .I(N__28932));
    InMux I__6178 (
            .O(N__28960),
            .I(N__28932));
    InMux I__6177 (
            .O(N__28959),
            .I(N__28932));
    InMux I__6176 (
            .O(N__28958),
            .I(N__28932));
    InMux I__6175 (
            .O(N__28957),
            .I(N__28927));
    InMux I__6174 (
            .O(N__28956),
            .I(N__28927));
    InMux I__6173 (
            .O(N__28955),
            .I(N__28924));
    Span4Mux_v I__6172 (
            .O(N__28950),
            .I(N__28917));
    Span4Mux_h I__6171 (
            .O(N__28945),
            .I(N__28917));
    LocalMux I__6170 (
            .O(N__28942),
            .I(N__28917));
    InMux I__6169 (
            .O(N__28941),
            .I(N__28914));
    LocalMux I__6168 (
            .O(N__28932),
            .I(N__28905));
    LocalMux I__6167 (
            .O(N__28927),
            .I(N__28902));
    LocalMux I__6166 (
            .O(N__28924),
            .I(N__28898));
    Span4Mux_h I__6165 (
            .O(N__28917),
            .I(N__28893));
    LocalMux I__6164 (
            .O(N__28914),
            .I(N__28893));
    InMux I__6163 (
            .O(N__28913),
            .I(N__28886));
    InMux I__6162 (
            .O(N__28912),
            .I(N__28886));
    InMux I__6161 (
            .O(N__28911),
            .I(N__28886));
    InMux I__6160 (
            .O(N__28910),
            .I(N__28882));
    InMux I__6159 (
            .O(N__28909),
            .I(N__28879));
    InMux I__6158 (
            .O(N__28908),
            .I(N__28876));
    Span4Mux_v I__6157 (
            .O(N__28905),
            .I(N__28871));
    Span4Mux_v I__6156 (
            .O(N__28902),
            .I(N__28871));
    InMux I__6155 (
            .O(N__28901),
            .I(N__28868));
    Span4Mux_v I__6154 (
            .O(N__28898),
            .I(N__28861));
    Span4Mux_v I__6153 (
            .O(N__28893),
            .I(N__28861));
    LocalMux I__6152 (
            .O(N__28886),
            .I(N__28861));
    InMux I__6151 (
            .O(N__28885),
            .I(N__28858));
    LocalMux I__6150 (
            .O(N__28882),
            .I(N__28847));
    LocalMux I__6149 (
            .O(N__28879),
            .I(N__28847));
    LocalMux I__6148 (
            .O(N__28876),
            .I(N__28847));
    Sp12to4 I__6147 (
            .O(N__28871),
            .I(N__28847));
    LocalMux I__6146 (
            .O(N__28868),
            .I(N__28847));
    Span4Mux_h I__6145 (
            .O(N__28861),
            .I(N__28842));
    LocalMux I__6144 (
            .O(N__28858),
            .I(N__28842));
    Span12Mux_s8_h I__6143 (
            .O(N__28847),
            .I(N__28839));
    IoSpan4Mux I__6142 (
            .O(N__28842),
            .I(N__28836));
    Odrv12 I__6141 (
            .O(N__28839),
            .I(slp_s4n));
    Odrv4 I__6140 (
            .O(N__28836),
            .I(slp_s4n));
    CascadeMux I__6139 (
            .O(N__28831),
            .I(\POWERLED.un1_func_state25_4_i_a2_0_cascade_ ));
    InMux I__6138 (
            .O(N__28828),
            .I(N__28824));
    CascadeMux I__6137 (
            .O(N__28827),
            .I(N__28821));
    LocalMux I__6136 (
            .O(N__28824),
            .I(N__28817));
    InMux I__6135 (
            .O(N__28821),
            .I(N__28814));
    CascadeMux I__6134 (
            .O(N__28820),
            .I(N__28811));
    Span4Mux_s3_h I__6133 (
            .O(N__28817),
            .I(N__28808));
    LocalMux I__6132 (
            .O(N__28814),
            .I(N__28805));
    InMux I__6131 (
            .O(N__28811),
            .I(N__28802));
    Odrv4 I__6130 (
            .O(N__28808),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0 ));
    Odrv4 I__6129 (
            .O(N__28805),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0 ));
    LocalMux I__6128 (
            .O(N__28802),
            .I(\POWERLED.func_state_RNIBVNSZ0Z_0 ));
    InMux I__6127 (
            .O(N__28795),
            .I(N__28792));
    LocalMux I__6126 (
            .O(N__28792),
            .I(\POWERLED.N_291 ));
    CascadeMux I__6125 (
            .O(N__28789),
            .I(\POWERLED.count_clk_en_0_cascade_ ));
    CascadeMux I__6124 (
            .O(N__28786),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ));
    CascadeMux I__6123 (
            .O(N__28783),
            .I(\POWERLED.count_clkZ0Z_0_cascade_ ));
    CascadeMux I__6122 (
            .O(N__28780),
            .I(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ));
    InMux I__6121 (
            .O(N__28777),
            .I(N__28774));
    LocalMux I__6120 (
            .O(N__28774),
            .I(\POWERLED.count_clk_0_4 ));
    CascadeMux I__6119 (
            .O(N__28771),
            .I(N__28768));
    InMux I__6118 (
            .O(N__28768),
            .I(N__28765));
    LocalMux I__6117 (
            .O(N__28765),
            .I(\POWERLED.count_clk_0_6 ));
    InMux I__6116 (
            .O(N__28762),
            .I(N__28759));
    LocalMux I__6115 (
            .O(N__28759),
            .I(\POWERLED.count_clk_0_0 ));
    InMux I__6114 (
            .O(N__28756),
            .I(N__28750));
    InMux I__6113 (
            .O(N__28755),
            .I(N__28750));
    LocalMux I__6112 (
            .O(N__28750),
            .I(N__28747));
    Span4Mux_h I__6111 (
            .O(N__28747),
            .I(N__28744));
    Odrv4 I__6110 (
            .O(N__28744),
            .I(\POWERLED.count_clk_RNIZ0Z_1 ));
    InMux I__6109 (
            .O(N__28741),
            .I(N__28738));
    LocalMux I__6108 (
            .O(N__28738),
            .I(\POWERLED.count_clk_0_3 ));
    CascadeMux I__6107 (
            .O(N__28735),
            .I(\POWERLED.count_clkZ0Z_14_cascade_ ));
    InMux I__6106 (
            .O(N__28732),
            .I(N__28729));
    LocalMux I__6105 (
            .O(N__28729),
            .I(\POWERLED.count_clk_0_13 ));
    InMux I__6104 (
            .O(N__28726),
            .I(N__28723));
    LocalMux I__6103 (
            .O(N__28723),
            .I(\POWERLED.count_clk_0_14 ));
    CascadeMux I__6102 (
            .O(N__28720),
            .I(\VPP_VDDQ.count_2_1_7_cascade_ ));
    InMux I__6101 (
            .O(N__28717),
            .I(N__28713));
    InMux I__6100 (
            .O(N__28716),
            .I(N__28710));
    LocalMux I__6099 (
            .O(N__28713),
            .I(N__28707));
    LocalMux I__6098 (
            .O(N__28710),
            .I(N__28704));
    Span4Mux_v I__6097 (
            .O(N__28707),
            .I(N__28701));
    Span4Mux_s2_h I__6096 (
            .O(N__28704),
            .I(N__28698));
    Odrv4 I__6095 (
            .O(N__28701),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    Odrv4 I__6094 (
            .O(N__28698),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    CascadeMux I__6093 (
            .O(N__28693),
            .I(\VPP_VDDQ.un9_clk_100khz_7_cascade_ ));
    InMux I__6092 (
            .O(N__28690),
            .I(N__28686));
    InMux I__6091 (
            .O(N__28689),
            .I(N__28683));
    LocalMux I__6090 (
            .O(N__28686),
            .I(N__28678));
    LocalMux I__6089 (
            .O(N__28683),
            .I(N__28678));
    Span4Mux_v I__6088 (
            .O(N__28678),
            .I(N__28675));
    Odrv4 I__6087 (
            .O(N__28675),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    InMux I__6086 (
            .O(N__28672),
            .I(N__28669));
    LocalMux I__6085 (
            .O(N__28669),
            .I(\VPP_VDDQ.count_2_1_7 ));
    InMux I__6084 (
            .O(N__28666),
            .I(N__28663));
    LocalMux I__6083 (
            .O(N__28663),
            .I(N__28660));
    Odrv4 I__6082 (
            .O(N__28660),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    InMux I__6081 (
            .O(N__28657),
            .I(N__28651));
    InMux I__6080 (
            .O(N__28656),
            .I(N__28651));
    LocalMux I__6079 (
            .O(N__28651),
            .I(N__28648));
    Odrv4 I__6078 (
            .O(N__28648),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ));
    InMux I__6077 (
            .O(N__28645),
            .I(N__28639));
    InMux I__6076 (
            .O(N__28644),
            .I(N__28639));
    LocalMux I__6075 (
            .O(N__28639),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    CascadeMux I__6074 (
            .O(N__28636),
            .I(\VPP_VDDQ.count_2_1_0_cascade_ ));
    CascadeMux I__6073 (
            .O(N__28633),
            .I(\VPP_VDDQ.count_2Z0Z_0_cascade_ ));
    InMux I__6072 (
            .O(N__28630),
            .I(N__28627));
    LocalMux I__6071 (
            .O(N__28627),
            .I(\VPP_VDDQ.count_2_0_0 ));
    InMux I__6070 (
            .O(N__28624),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__6069 (
            .O(N__28621),
            .I(N__28618));
    LocalMux I__6068 (
            .O(N__28618),
            .I(N__28614));
    InMux I__6067 (
            .O(N__28617),
            .I(N__28611));
    Span4Mux_s3_h I__6066 (
            .O(N__28614),
            .I(N__28608));
    LocalMux I__6065 (
            .O(N__28611),
            .I(N__28605));
    Odrv4 I__6064 (
            .O(N__28608),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    Odrv12 I__6063 (
            .O(N__28605),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    CascadeMux I__6062 (
            .O(N__28600),
            .I(N__28596));
    CascadeMux I__6061 (
            .O(N__28599),
            .I(N__28593));
    InMux I__6060 (
            .O(N__28596),
            .I(N__28588));
    InMux I__6059 (
            .O(N__28593),
            .I(N__28588));
    LocalMux I__6058 (
            .O(N__28588),
            .I(N__28585));
    Odrv4 I__6057 (
            .O(N__28585),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ));
    InMux I__6056 (
            .O(N__28582),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    CascadeMux I__6055 (
            .O(N__28579),
            .I(N__28575));
    InMux I__6054 (
            .O(N__28578),
            .I(N__28570));
    InMux I__6053 (
            .O(N__28575),
            .I(N__28570));
    LocalMux I__6052 (
            .O(N__28570),
            .I(N__28567));
    Span4Mux_v I__6051 (
            .O(N__28567),
            .I(N__28564));
    Odrv4 I__6050 (
            .O(N__28564),
            .I(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ));
    InMux I__6049 (
            .O(N__28561),
            .I(bfn_11_7_0_));
    CascadeMux I__6048 (
            .O(N__28558),
            .I(N__28554));
    CascadeMux I__6047 (
            .O(N__28557),
            .I(N__28551));
    InMux I__6046 (
            .O(N__28554),
            .I(N__28548));
    InMux I__6045 (
            .O(N__28551),
            .I(N__28545));
    LocalMux I__6044 (
            .O(N__28548),
            .I(N__28542));
    LocalMux I__6043 (
            .O(N__28545),
            .I(N__28539));
    Span4Mux_v I__6042 (
            .O(N__28542),
            .I(N__28536));
    Span4Mux_h I__6041 (
            .O(N__28539),
            .I(N__28533));
    Odrv4 I__6040 (
            .O(N__28536),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ));
    Odrv4 I__6039 (
            .O(N__28533),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ));
    InMux I__6038 (
            .O(N__28528),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__6037 (
            .O(N__28525),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__6036 (
            .O(N__28522),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    InMux I__6035 (
            .O(N__28519),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    InMux I__6034 (
            .O(N__28516),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__6033 (
            .O(N__28513),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    CascadeMux I__6032 (
            .O(N__28510),
            .I(N__28506));
    InMux I__6031 (
            .O(N__28509),
            .I(N__28501));
    InMux I__6030 (
            .O(N__28506),
            .I(N__28501));
    LocalMux I__6029 (
            .O(N__28501),
            .I(N__28498));
    Odrv4 I__6028 (
            .O(N__28498),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ));
    CascadeMux I__6027 (
            .O(N__28495),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ));
    InMux I__6026 (
            .O(N__28492),
            .I(N__28489));
    LocalMux I__6025 (
            .O(N__28489),
            .I(\VPP_VDDQ.count_2_0_15 ));
    InMux I__6024 (
            .O(N__28486),
            .I(N__28483));
    LocalMux I__6023 (
            .O(N__28483),
            .I(\VPP_VDDQ.count_2_0_3 ));
    InMux I__6022 (
            .O(N__28480),
            .I(N__28477));
    LocalMux I__6021 (
            .O(N__28477),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    CascadeMux I__6020 (
            .O(N__28474),
            .I(N__28470));
    InMux I__6019 (
            .O(N__28473),
            .I(N__28465));
    InMux I__6018 (
            .O(N__28470),
            .I(N__28465));
    LocalMux I__6017 (
            .O(N__28465),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ));
    InMux I__6016 (
            .O(N__28462),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    InMux I__6015 (
            .O(N__28459),
            .I(N__28455));
    InMux I__6014 (
            .O(N__28458),
            .I(N__28452));
    LocalMux I__6013 (
            .O(N__28455),
            .I(N__28449));
    LocalMux I__6012 (
            .O(N__28452),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    Odrv4 I__6011 (
            .O(N__28449),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    InMux I__6010 (
            .O(N__28444),
            .I(N__28440));
    InMux I__6009 (
            .O(N__28443),
            .I(N__28437));
    LocalMux I__6008 (
            .O(N__28440),
            .I(N__28434));
    LocalMux I__6007 (
            .O(N__28437),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    Odrv4 I__6006 (
            .O(N__28434),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ));
    InMux I__6005 (
            .O(N__28429),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__6004 (
            .O(N__28426),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    InMux I__6003 (
            .O(N__28423),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    InMux I__6002 (
            .O(N__28420),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    CascadeMux I__6001 (
            .O(N__28417),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    InMux I__6000 (
            .O(N__28414),
            .I(N__28411));
    LocalMux I__5999 (
            .O(N__28411),
            .I(\VPP_VDDQ.curr_state_2_0_1 ));
    CascadeMux I__5998 (
            .O(N__28408),
            .I(\VPP_VDDQ.N_55_cascade_ ));
    CascadeMux I__5997 (
            .O(N__28405),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ));
    CascadeMux I__5996 (
            .O(N__28402),
            .I(\VPP_VDDQ.count_2_1_3_cascade_ ));
    CascadeMux I__5995 (
            .O(N__28399),
            .I(\VPP_VDDQ.count_2_1_2_cascade_ ));
    InMux I__5994 (
            .O(N__28396),
            .I(N__28393));
    LocalMux I__5993 (
            .O(N__28393),
            .I(\VPP_VDDQ.count_2_0_2 ));
    CascadeMux I__5992 (
            .O(N__28390),
            .I(\VPP_VDDQ.count_2Z0Z_2_cascade_ ));
    CascadeMux I__5991 (
            .O(N__28387),
            .I(G_1939_cascade_));
    InMux I__5990 (
            .O(N__28384),
            .I(N__28380));
    InMux I__5989 (
            .O(N__28383),
            .I(N__28377));
    LocalMux I__5988 (
            .O(N__28380),
            .I(N__28373));
    LocalMux I__5987 (
            .O(N__28377),
            .I(N__28370));
    InMux I__5986 (
            .O(N__28376),
            .I(N__28367));
    Span4Mux_h I__5985 (
            .O(N__28373),
            .I(N__28362));
    Span4Mux_s2_h I__5984 (
            .O(N__28370),
            .I(N__28362));
    LocalMux I__5983 (
            .O(N__28367),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__5982 (
            .O(N__28362),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__5981 (
            .O(N__28357),
            .I(N__28354));
    LocalMux I__5980 (
            .O(N__28354),
            .I(N__28350));
    InMux I__5979 (
            .O(N__28353),
            .I(N__28347));
    Span4Mux_s2_v I__5978 (
            .O(N__28350),
            .I(N__28344));
    LocalMux I__5977 (
            .O(N__28347),
            .I(N_218));
    Odrv4 I__5976 (
            .O(N__28344),
            .I(N_218));
    InMux I__5975 (
            .O(N__28339),
            .I(N__28336));
    LocalMux I__5974 (
            .O(N__28336),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    InMux I__5973 (
            .O(N__28333),
            .I(N__28327));
    InMux I__5972 (
            .O(N__28332),
            .I(N__28327));
    LocalMux I__5971 (
            .O(N__28327),
            .I(N__28323));
    InMux I__5970 (
            .O(N__28326),
            .I(N__28320));
    Span4Mux_h I__5969 (
            .O(N__28323),
            .I(N__28317));
    LocalMux I__5968 (
            .O(N__28320),
            .I(G_1939));
    Odrv4 I__5967 (
            .O(N__28317),
            .I(G_1939));
    CascadeMux I__5966 (
            .O(N__28312),
            .I(N_218_cascade_));
    InMux I__5965 (
            .O(N__28309),
            .I(N__28306));
    LocalMux I__5964 (
            .O(N__28306),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    CascadeMux I__5963 (
            .O(N__28303),
            .I(\PCH_PWRGD.curr_state_0_1_cascade_ ));
    InMux I__5962 (
            .O(N__28300),
            .I(N__28294));
    InMux I__5961 (
            .O(N__28299),
            .I(N__28294));
    LocalMux I__5960 (
            .O(N__28294),
            .I(N__28291));
    Span4Mux_s2_v I__5959 (
            .O(N__28291),
            .I(N__28287));
    InMux I__5958 (
            .O(N__28290),
            .I(N__28284));
    Odrv4 I__5957 (
            .O(N__28287),
            .I(\PCH_PWRGD.N_2190_i ));
    LocalMux I__5956 (
            .O(N__28284),
            .I(\PCH_PWRGD.N_2190_i ));
    InMux I__5955 (
            .O(N__28279),
            .I(N__28275));
    InMux I__5954 (
            .O(N__28278),
            .I(N__28272));
    LocalMux I__5953 (
            .O(N__28275),
            .I(N__28267));
    LocalMux I__5952 (
            .O(N__28272),
            .I(N__28264));
    InMux I__5951 (
            .O(N__28271),
            .I(N__28261));
    InMux I__5950 (
            .O(N__28270),
            .I(N__28258));
    Span4Mux_s3_v I__5949 (
            .O(N__28267),
            .I(N__28253));
    Span4Mux_s3_v I__5948 (
            .O(N__28264),
            .I(N__28253));
    LocalMux I__5947 (
            .O(N__28261),
            .I(\PCH_PWRGD.N_2171_i ));
    LocalMux I__5946 (
            .O(N__28258),
            .I(\PCH_PWRGD.N_2171_i ));
    Odrv4 I__5945 (
            .O(N__28253),
            .I(\PCH_PWRGD.N_2171_i ));
    CascadeMux I__5944 (
            .O(N__28246),
            .I(\PCH_PWRGD.N_2190_i_cascade_ ));
    SRMux I__5943 (
            .O(N__28243),
            .I(N__28236));
    InMux I__5942 (
            .O(N__28242),
            .I(N__28229));
    SRMux I__5941 (
            .O(N__28241),
            .I(N__28229));
    CascadeMux I__5940 (
            .O(N__28240),
            .I(N__28219));
    CascadeMux I__5939 (
            .O(N__28239),
            .I(N__28213));
    LocalMux I__5938 (
            .O(N__28236),
            .I(N__28200));
    CascadeMux I__5937 (
            .O(N__28235),
            .I(N__28197));
    CascadeMux I__5936 (
            .O(N__28234),
            .I(N__28194));
    LocalMux I__5935 (
            .O(N__28229),
            .I(N__28190));
    SRMux I__5934 (
            .O(N__28228),
            .I(N__28187));
    InMux I__5933 (
            .O(N__28227),
            .I(N__28182));
    SRMux I__5932 (
            .O(N__28226),
            .I(N__28182));
    InMux I__5931 (
            .O(N__28225),
            .I(N__28179));
    InMux I__5930 (
            .O(N__28224),
            .I(N__28174));
    InMux I__5929 (
            .O(N__28223),
            .I(N__28174));
    InMux I__5928 (
            .O(N__28222),
            .I(N__28171));
    InMux I__5927 (
            .O(N__28219),
            .I(N__28163));
    InMux I__5926 (
            .O(N__28218),
            .I(N__28160));
    SRMux I__5925 (
            .O(N__28217),
            .I(N__28151));
    InMux I__5924 (
            .O(N__28216),
            .I(N__28151));
    InMux I__5923 (
            .O(N__28213),
            .I(N__28151));
    InMux I__5922 (
            .O(N__28212),
            .I(N__28151));
    InMux I__5921 (
            .O(N__28211),
            .I(N__28140));
    InMux I__5920 (
            .O(N__28210),
            .I(N__28140));
    InMux I__5919 (
            .O(N__28209),
            .I(N__28140));
    InMux I__5918 (
            .O(N__28208),
            .I(N__28140));
    InMux I__5917 (
            .O(N__28207),
            .I(N__28140));
    InMux I__5916 (
            .O(N__28206),
            .I(N__28131));
    InMux I__5915 (
            .O(N__28205),
            .I(N__28131));
    InMux I__5914 (
            .O(N__28204),
            .I(N__28131));
    InMux I__5913 (
            .O(N__28203),
            .I(N__28131));
    Span4Mux_s3_v I__5912 (
            .O(N__28200),
            .I(N__28128));
    InMux I__5911 (
            .O(N__28197),
            .I(N__28121));
    InMux I__5910 (
            .O(N__28194),
            .I(N__28121));
    InMux I__5909 (
            .O(N__28193),
            .I(N__28121));
    Span4Mux_v I__5908 (
            .O(N__28190),
            .I(N__28114));
    LocalMux I__5907 (
            .O(N__28187),
            .I(N__28114));
    LocalMux I__5906 (
            .O(N__28182),
            .I(N__28114));
    LocalMux I__5905 (
            .O(N__28179),
            .I(N__28107));
    LocalMux I__5904 (
            .O(N__28174),
            .I(N__28107));
    LocalMux I__5903 (
            .O(N__28171),
            .I(N__28107));
    SRMux I__5902 (
            .O(N__28170),
            .I(N__28098));
    InMux I__5901 (
            .O(N__28169),
            .I(N__28098));
    InMux I__5900 (
            .O(N__28168),
            .I(N__28098));
    InMux I__5899 (
            .O(N__28167),
            .I(N__28098));
    InMux I__5898 (
            .O(N__28166),
            .I(N__28095));
    LocalMux I__5897 (
            .O(N__28163),
            .I(N__28084));
    LocalMux I__5896 (
            .O(N__28160),
            .I(N__28084));
    LocalMux I__5895 (
            .O(N__28151),
            .I(N__28084));
    LocalMux I__5894 (
            .O(N__28140),
            .I(N__28084));
    LocalMux I__5893 (
            .O(N__28131),
            .I(N__28084));
    Span4Mux_h I__5892 (
            .O(N__28128),
            .I(N__28080));
    LocalMux I__5891 (
            .O(N__28121),
            .I(N__28075));
    Span4Mux_h I__5890 (
            .O(N__28114),
            .I(N__28075));
    Span4Mux_s2_v I__5889 (
            .O(N__28107),
            .I(N__28072));
    LocalMux I__5888 (
            .O(N__28098),
            .I(N__28069));
    LocalMux I__5887 (
            .O(N__28095),
            .I(N__28064));
    Span4Mux_s2_v I__5886 (
            .O(N__28084),
            .I(N__28064));
    InMux I__5885 (
            .O(N__28083),
            .I(N__28061));
    Odrv4 I__5884 (
            .O(N__28080),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__5883 (
            .O(N__28075),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__5882 (
            .O(N__28072),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__5881 (
            .O(N__28069),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__5880 (
            .O(N__28064),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__5879 (
            .O(N__28061),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    InMux I__5878 (
            .O(N__28048),
            .I(N__28045));
    LocalMux I__5877 (
            .O(N__28045),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    CascadeMux I__5876 (
            .O(N__28042),
            .I(\VPP_VDDQ.N_53_cascade_ ));
    InMux I__5875 (
            .O(N__28039),
            .I(N__28036));
    LocalMux I__5874 (
            .O(N__28036),
            .I(\PCH_PWRGD.count_rst_7 ));
    CascadeMux I__5873 (
            .O(N__28033),
            .I(\PCH_PWRGD.count_rst_7_cascade_ ));
    InMux I__5872 (
            .O(N__28030),
            .I(N__28027));
    LocalMux I__5871 (
            .O(N__28027),
            .I(\PCH_PWRGD.count_1_i_a2_5_0 ));
    InMux I__5870 (
            .O(N__28024),
            .I(N__28018));
    InMux I__5869 (
            .O(N__28023),
            .I(N__28018));
    LocalMux I__5868 (
            .O(N__28018),
            .I(N__28015));
    Span4Mux_s3_h I__5867 (
            .O(N__28015),
            .I(N__28012));
    Odrv4 I__5866 (
            .O(N__28012),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    CascadeMux I__5865 (
            .O(N__28009),
            .I(N__28006));
    InMux I__5864 (
            .O(N__28006),
            .I(N__28003));
    LocalMux I__5863 (
            .O(N__28003),
            .I(N__27998));
    InMux I__5862 (
            .O(N__28002),
            .I(N__27993));
    InMux I__5861 (
            .O(N__28001),
            .I(N__27993));
    Span4Mux_s1_v I__5860 (
            .O(N__27998),
            .I(N__27990));
    LocalMux I__5859 (
            .O(N__27993),
            .I(\PCH_PWRGD.un2_count_1_axb_7 ));
    Odrv4 I__5858 (
            .O(N__27990),
            .I(\PCH_PWRGD.un2_count_1_axb_7 ));
    InMux I__5857 (
            .O(N__27985),
            .I(N__27979));
    InMux I__5856 (
            .O(N__27984),
            .I(N__27979));
    LocalMux I__5855 (
            .O(N__27979),
            .I(\PCH_PWRGD.count_0_7 ));
    CascadeMux I__5854 (
            .O(N__27976),
            .I(\PCH_PWRGD.count_rst_9_cascade_ ));
    InMux I__5853 (
            .O(N__27973),
            .I(N__27970));
    LocalMux I__5852 (
            .O(N__27970),
            .I(N__27967));
    Span4Mux_s1_v I__5851 (
            .O(N__27967),
            .I(N__27962));
    InMux I__5850 (
            .O(N__27966),
            .I(N__27957));
    InMux I__5849 (
            .O(N__27965),
            .I(N__27957));
    Odrv4 I__5848 (
            .O(N__27962),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__5847 (
            .O(N__27957),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    CascadeMux I__5846 (
            .O(N__27952),
            .I(N__27949));
    InMux I__5845 (
            .O(N__27949),
            .I(N__27943));
    InMux I__5844 (
            .O(N__27948),
            .I(N__27943));
    LocalMux I__5843 (
            .O(N__27943),
            .I(N__27940));
    Span4Mux_v I__5842 (
            .O(N__27940),
            .I(N__27937));
    Odrv4 I__5841 (
            .O(N__27937),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__5840 (
            .O(N__27934),
            .I(\PCH_PWRGD.countZ0Z_5_cascade_ ));
    InMux I__5839 (
            .O(N__27931),
            .I(N__27928));
    LocalMux I__5838 (
            .O(N__27928),
            .I(\PCH_PWRGD.count_0_5 ));
    InMux I__5837 (
            .O(N__27925),
            .I(N__27922));
    LocalMux I__5836 (
            .O(N__27922),
            .I(N__27918));
    InMux I__5835 (
            .O(N__27921),
            .I(N__27915));
    Odrv4 I__5834 (
            .O(N__27918),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    LocalMux I__5833 (
            .O(N__27915),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    CascadeMux I__5832 (
            .O(N__27910),
            .I(N__27906));
    InMux I__5831 (
            .O(N__27909),
            .I(N__27902));
    InMux I__5830 (
            .O(N__27906),
            .I(N__27899));
    CascadeMux I__5829 (
            .O(N__27905),
            .I(N__27895));
    LocalMux I__5828 (
            .O(N__27902),
            .I(N__27890));
    LocalMux I__5827 (
            .O(N__27899),
            .I(N__27890));
    CascadeMux I__5826 (
            .O(N__27898),
            .I(N__27887));
    InMux I__5825 (
            .O(N__27895),
            .I(N__27884));
    Span4Mux_s2_v I__5824 (
            .O(N__27890),
            .I(N__27881));
    InMux I__5823 (
            .O(N__27887),
            .I(N__27878));
    LocalMux I__5822 (
            .O(N__27884),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    Odrv4 I__5821 (
            .O(N__27881),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    LocalMux I__5820 (
            .O(N__27878),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    InMux I__5819 (
            .O(N__27871),
            .I(N__27868));
    LocalMux I__5818 (
            .O(N__27868),
            .I(N__27865));
    Span4Mux_h I__5817 (
            .O(N__27865),
            .I(N__27862));
    Odrv4 I__5816 (
            .O(N__27862),
            .I(\PCH_PWRGD.count_0_11 ));
    CEMux I__5815 (
            .O(N__27859),
            .I(N__27853));
    CascadeMux I__5814 (
            .O(N__27858),
            .I(N__27846));
    InMux I__5813 (
            .O(N__27857),
            .I(N__27839));
    CEMux I__5812 (
            .O(N__27856),
            .I(N__27839));
    LocalMux I__5811 (
            .O(N__27853),
            .I(N__27835));
    InMux I__5810 (
            .O(N__27852),
            .I(N__27822));
    InMux I__5809 (
            .O(N__27851),
            .I(N__27822));
    InMux I__5808 (
            .O(N__27850),
            .I(N__27822));
    InMux I__5807 (
            .O(N__27849),
            .I(N__27822));
    InMux I__5806 (
            .O(N__27846),
            .I(N__27815));
    CEMux I__5805 (
            .O(N__27845),
            .I(N__27815));
    CEMux I__5804 (
            .O(N__27844),
            .I(N__27812));
    LocalMux I__5803 (
            .O(N__27839),
            .I(N__27799));
    CEMux I__5802 (
            .O(N__27838),
            .I(N__27796));
    Span4Mux_s1_v I__5801 (
            .O(N__27835),
            .I(N__27793));
    CEMux I__5800 (
            .O(N__27834),
            .I(N__27784));
    InMux I__5799 (
            .O(N__27833),
            .I(N__27784));
    InMux I__5798 (
            .O(N__27832),
            .I(N__27784));
    InMux I__5797 (
            .O(N__27831),
            .I(N__27784));
    LocalMux I__5796 (
            .O(N__27822),
            .I(N__27781));
    InMux I__5795 (
            .O(N__27821),
            .I(N__27776));
    InMux I__5794 (
            .O(N__27820),
            .I(N__27773));
    LocalMux I__5793 (
            .O(N__27815),
            .I(N__27770));
    LocalMux I__5792 (
            .O(N__27812),
            .I(N__27767));
    InMux I__5791 (
            .O(N__27811),
            .I(N__27764));
    InMux I__5790 (
            .O(N__27810),
            .I(N__27755));
    InMux I__5789 (
            .O(N__27809),
            .I(N__27755));
    InMux I__5788 (
            .O(N__27808),
            .I(N__27755));
    InMux I__5787 (
            .O(N__27807),
            .I(N__27755));
    InMux I__5786 (
            .O(N__27806),
            .I(N__27750));
    InMux I__5785 (
            .O(N__27805),
            .I(N__27750));
    InMux I__5784 (
            .O(N__27804),
            .I(N__27743));
    InMux I__5783 (
            .O(N__27803),
            .I(N__27743));
    InMux I__5782 (
            .O(N__27802),
            .I(N__27743));
    Span4Mux_s1_h I__5781 (
            .O(N__27799),
            .I(N__27732));
    LocalMux I__5780 (
            .O(N__27796),
            .I(N__27732));
    Span4Mux_s1_h I__5779 (
            .O(N__27793),
            .I(N__27732));
    LocalMux I__5778 (
            .O(N__27784),
            .I(N__27732));
    Span4Mux_s1_v I__5777 (
            .O(N__27781),
            .I(N__27732));
    InMux I__5776 (
            .O(N__27780),
            .I(N__27727));
    InMux I__5775 (
            .O(N__27779),
            .I(N__27727));
    LocalMux I__5774 (
            .O(N__27776),
            .I(N__27722));
    LocalMux I__5773 (
            .O(N__27773),
            .I(N__27722));
    Odrv4 I__5772 (
            .O(N__27770),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    Odrv4 I__5771 (
            .O(N__27767),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    LocalMux I__5770 (
            .O(N__27764),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    LocalMux I__5769 (
            .O(N__27755),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    LocalMux I__5768 (
            .O(N__27750),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    LocalMux I__5767 (
            .O(N__27743),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    Odrv4 I__5766 (
            .O(N__27732),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    LocalMux I__5765 (
            .O(N__27727),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    Odrv12 I__5764 (
            .O(N__27722),
            .I(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ));
    InMux I__5763 (
            .O(N__27703),
            .I(N__27686));
    InMux I__5762 (
            .O(N__27702),
            .I(N__27686));
    InMux I__5761 (
            .O(N__27701),
            .I(N__27674));
    InMux I__5760 (
            .O(N__27700),
            .I(N__27674));
    InMux I__5759 (
            .O(N__27699),
            .I(N__27674));
    InMux I__5758 (
            .O(N__27698),
            .I(N__27674));
    InMux I__5757 (
            .O(N__27697),
            .I(N__27674));
    InMux I__5756 (
            .O(N__27696),
            .I(N__27671));
    InMux I__5755 (
            .O(N__27695),
            .I(N__27659));
    InMux I__5754 (
            .O(N__27694),
            .I(N__27659));
    InMux I__5753 (
            .O(N__27693),
            .I(N__27659));
    InMux I__5752 (
            .O(N__27692),
            .I(N__27659));
    InMux I__5751 (
            .O(N__27691),
            .I(N__27659));
    LocalMux I__5750 (
            .O(N__27686),
            .I(N__27656));
    InMux I__5749 (
            .O(N__27685),
            .I(N__27653));
    LocalMux I__5748 (
            .O(N__27674),
            .I(N__27648));
    LocalMux I__5747 (
            .O(N__27671),
            .I(N__27648));
    InMux I__5746 (
            .O(N__27670),
            .I(N__27645));
    LocalMux I__5745 (
            .O(N__27659),
            .I(N__27642));
    Span4Mux_s2_v I__5744 (
            .O(N__27656),
            .I(N__27633));
    LocalMux I__5743 (
            .O(N__27653),
            .I(N__27633));
    Span4Mux_s2_v I__5742 (
            .O(N__27648),
            .I(N__27633));
    LocalMux I__5741 (
            .O(N__27645),
            .I(N__27633));
    Odrv4 I__5740 (
            .O(N__27642),
            .I(\PCH_PWRGD.N_364 ));
    Odrv4 I__5739 (
            .O(N__27633),
            .I(\PCH_PWRGD.N_364 ));
    CascadeMux I__5738 (
            .O(N__27628),
            .I(N__27625));
    InMux I__5737 (
            .O(N__27625),
            .I(N__27621));
    InMux I__5736 (
            .O(N__27624),
            .I(N__27618));
    LocalMux I__5735 (
            .O(N__27621),
            .I(N__27615));
    LocalMux I__5734 (
            .O(N__27618),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    Odrv12 I__5733 (
            .O(N__27615),
            .I(\PCH_PWRGD.un2_count_1_axb_1 ));
    CascadeMux I__5732 (
            .O(N__27610),
            .I(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ));
    InMux I__5731 (
            .O(N__27607),
            .I(N__27600));
    InMux I__5730 (
            .O(N__27606),
            .I(N__27600));
    InMux I__5729 (
            .O(N__27605),
            .I(N__27597));
    LocalMux I__5728 (
            .O(N__27600),
            .I(N__27594));
    LocalMux I__5727 (
            .O(N__27597),
            .I(N__27591));
    Span4Mux_s2_h I__5726 (
            .O(N__27594),
            .I(N__27588));
    Odrv4 I__5725 (
            .O(N__27591),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    Odrv4 I__5724 (
            .O(N__27588),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    InMux I__5723 (
            .O(N__27583),
            .I(N__27580));
    LocalMux I__5722 (
            .O(N__27580),
            .I(\PCH_PWRGD.count_rst_13 ));
    InMux I__5721 (
            .O(N__27577),
            .I(N__27571));
    InMux I__5720 (
            .O(N__27576),
            .I(N__27571));
    LocalMux I__5719 (
            .O(N__27571),
            .I(\PCH_PWRGD.count_0_1 ));
    CascadeMux I__5718 (
            .O(N__27568),
            .I(\PCH_PWRGD.count_rst_13_cascade_ ));
    InMux I__5717 (
            .O(N__27565),
            .I(N__27562));
    LocalMux I__5716 (
            .O(N__27562),
            .I(N__27559));
    Odrv4 I__5715 (
            .O(N__27559),
            .I(\PCH_PWRGD.count_1_i_a2_6_0 ));
    CascadeMux I__5714 (
            .O(N__27556),
            .I(\PCH_PWRGD.count_1_i_a2_3_0_cascade_ ));
    InMux I__5713 (
            .O(N__27553),
            .I(N__27546));
    InMux I__5712 (
            .O(N__27552),
            .I(N__27546));
    InMux I__5711 (
            .O(N__27551),
            .I(N__27543));
    LocalMux I__5710 (
            .O(N__27546),
            .I(N__27540));
    LocalMux I__5709 (
            .O(N__27543),
            .I(N__27537));
    Span4Mux_v I__5708 (
            .O(N__27540),
            .I(N__27534));
    Span4Mux_h I__5707 (
            .O(N__27537),
            .I(N__27531));
    Odrv4 I__5706 (
            .O(N__27534),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    Odrv4 I__5705 (
            .O(N__27531),
            .I(\PCH_PWRGD.count_1_i_a2_12_0 ));
    CascadeMux I__5704 (
            .O(N__27526),
            .I(N__27522));
    InMux I__5703 (
            .O(N__27525),
            .I(N__27519));
    InMux I__5702 (
            .O(N__27522),
            .I(N__27516));
    LocalMux I__5701 (
            .O(N__27519),
            .I(N__27513));
    LocalMux I__5700 (
            .O(N__27516),
            .I(N__27508));
    Span4Mux_v I__5699 (
            .O(N__27513),
            .I(N__27508));
    Odrv4 I__5698 (
            .O(N__27508),
            .I(\PCH_PWRGD.un2_count_1_axb_9 ));
    InMux I__5697 (
            .O(N__27505),
            .I(N__27502));
    LocalMux I__5696 (
            .O(N__27502),
            .I(N__27498));
    InMux I__5695 (
            .O(N__27501),
            .I(N__27495));
    Span4Mux_s1_v I__5694 (
            .O(N__27498),
            .I(N__27492));
    LocalMux I__5693 (
            .O(N__27495),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    Odrv4 I__5692 (
            .O(N__27492),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__5691 (
            .O(N__27487),
            .I(\PCH_PWRGD.un2_count_1_axb_9_cascade_ ));
    InMux I__5690 (
            .O(N__27484),
            .I(N__27481));
    LocalMux I__5689 (
            .O(N__27481),
            .I(\PCH_PWRGD.count_rst_5 ));
    InMux I__5688 (
            .O(N__27478),
            .I(N__27472));
    InMux I__5687 (
            .O(N__27477),
            .I(N__27472));
    LocalMux I__5686 (
            .O(N__27472),
            .I(N__27469));
    Odrv4 I__5685 (
            .O(N__27469),
            .I(\PCH_PWRGD.count_0_9 ));
    InMux I__5684 (
            .O(N__27466),
            .I(N__27461));
    CascadeMux I__5683 (
            .O(N__27465),
            .I(N__27458));
    CascadeMux I__5682 (
            .O(N__27464),
            .I(N__27455));
    LocalMux I__5681 (
            .O(N__27461),
            .I(N__27452));
    InMux I__5680 (
            .O(N__27458),
            .I(N__27449));
    InMux I__5679 (
            .O(N__27455),
            .I(N__27446));
    Odrv12 I__5678 (
            .O(N__27452),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__5677 (
            .O(N__27449),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__5676 (
            .O(N__27446),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    CascadeMux I__5675 (
            .O(N__27439),
            .I(\PCH_PWRGD.count_rst_5_cascade_ ));
    InMux I__5674 (
            .O(N__27436),
            .I(N__27433));
    LocalMux I__5673 (
            .O(N__27433),
            .I(\PCH_PWRGD.count_1_i_a2_4_0 ));
    InMux I__5672 (
            .O(N__27430),
            .I(N__27425));
    InMux I__5671 (
            .O(N__27429),
            .I(N__27416));
    InMux I__5670 (
            .O(N__27428),
            .I(N__27413));
    LocalMux I__5669 (
            .O(N__27425),
            .I(N__27408));
    InMux I__5668 (
            .O(N__27424),
            .I(N__27403));
    InMux I__5667 (
            .O(N__27423),
            .I(N__27403));
    InMux I__5666 (
            .O(N__27422),
            .I(N__27400));
    InMux I__5665 (
            .O(N__27421),
            .I(N__27397));
    InMux I__5664 (
            .O(N__27420),
            .I(N__27392));
    InMux I__5663 (
            .O(N__27419),
            .I(N__27392));
    LocalMux I__5662 (
            .O(N__27416),
            .I(N__27387));
    LocalMux I__5661 (
            .O(N__27413),
            .I(N__27387));
    InMux I__5660 (
            .O(N__27412),
            .I(N__27384));
    CascadeMux I__5659 (
            .O(N__27411),
            .I(N__27381));
    Span4Mux_v I__5658 (
            .O(N__27408),
            .I(N__27378));
    LocalMux I__5657 (
            .O(N__27403),
            .I(N__27375));
    LocalMux I__5656 (
            .O(N__27400),
            .I(N__27366));
    LocalMux I__5655 (
            .O(N__27397),
            .I(N__27366));
    LocalMux I__5654 (
            .O(N__27392),
            .I(N__27366));
    Span4Mux_v I__5653 (
            .O(N__27387),
            .I(N__27366));
    LocalMux I__5652 (
            .O(N__27384),
            .I(N__27363));
    InMux I__5651 (
            .O(N__27381),
            .I(N__27360));
    Odrv4 I__5650 (
            .O(N__27378),
            .I(\POWERLED.func_state_RNIZ0Z_1 ));
    Odrv4 I__5649 (
            .O(N__27375),
            .I(\POWERLED.func_state_RNIZ0Z_1 ));
    Odrv4 I__5648 (
            .O(N__27366),
            .I(\POWERLED.func_state_RNIZ0Z_1 ));
    Odrv4 I__5647 (
            .O(N__27363),
            .I(\POWERLED.func_state_RNIZ0Z_1 ));
    LocalMux I__5646 (
            .O(N__27360),
            .I(\POWERLED.func_state_RNIZ0Z_1 ));
    CascadeMux I__5645 (
            .O(N__27349),
            .I(N__27342));
    CascadeMux I__5644 (
            .O(N__27348),
            .I(N__27336));
    InMux I__5643 (
            .O(N__27347),
            .I(N__27326));
    InMux I__5642 (
            .O(N__27346),
            .I(N__27326));
    InMux I__5641 (
            .O(N__27345),
            .I(N__27326));
    InMux I__5640 (
            .O(N__27342),
            .I(N__27323));
    InMux I__5639 (
            .O(N__27341),
            .I(N__27320));
    InMux I__5638 (
            .O(N__27340),
            .I(N__27316));
    CascadeMux I__5637 (
            .O(N__27339),
            .I(N__27312));
    InMux I__5636 (
            .O(N__27336),
            .I(N__27307));
    InMux I__5635 (
            .O(N__27335),
            .I(N__27307));
    CascadeMux I__5634 (
            .O(N__27334),
            .I(N__27304));
    CascadeMux I__5633 (
            .O(N__27333),
            .I(N__27299));
    LocalMux I__5632 (
            .O(N__27326),
            .I(N__27292));
    LocalMux I__5631 (
            .O(N__27323),
            .I(N__27292));
    LocalMux I__5630 (
            .O(N__27320),
            .I(N__27292));
    InMux I__5629 (
            .O(N__27319),
            .I(N__27289));
    LocalMux I__5628 (
            .O(N__27316),
            .I(N__27286));
    InMux I__5627 (
            .O(N__27315),
            .I(N__27281));
    InMux I__5626 (
            .O(N__27312),
            .I(N__27281));
    LocalMux I__5625 (
            .O(N__27307),
            .I(N__27278));
    InMux I__5624 (
            .O(N__27304),
            .I(N__27274));
    InMux I__5623 (
            .O(N__27303),
            .I(N__27269));
    InMux I__5622 (
            .O(N__27302),
            .I(N__27269));
    InMux I__5621 (
            .O(N__27299),
            .I(N__27266));
    Span4Mux_v I__5620 (
            .O(N__27292),
            .I(N__27259));
    LocalMux I__5619 (
            .O(N__27289),
            .I(N__27259));
    Span4Mux_h I__5618 (
            .O(N__27286),
            .I(N__27254));
    LocalMux I__5617 (
            .O(N__27281),
            .I(N__27254));
    Span4Mux_v I__5616 (
            .O(N__27278),
            .I(N__27251));
    InMux I__5615 (
            .O(N__27277),
            .I(N__27248));
    LocalMux I__5614 (
            .O(N__27274),
            .I(N__27243));
    LocalMux I__5613 (
            .O(N__27269),
            .I(N__27243));
    LocalMux I__5612 (
            .O(N__27266),
            .I(N__27240));
    InMux I__5611 (
            .O(N__27265),
            .I(N__27237));
    InMux I__5610 (
            .O(N__27264),
            .I(N__27234));
    Span4Mux_v I__5609 (
            .O(N__27259),
            .I(N__27231));
    Span4Mux_h I__5608 (
            .O(N__27254),
            .I(N__27228));
    Span4Mux_v I__5607 (
            .O(N__27251),
            .I(N__27223));
    LocalMux I__5606 (
            .O(N__27248),
            .I(N__27223));
    Span4Mux_v I__5605 (
            .O(N__27243),
            .I(N__27216));
    Span4Mux_h I__5604 (
            .O(N__27240),
            .I(N__27216));
    LocalMux I__5603 (
            .O(N__27237),
            .I(N__27216));
    LocalMux I__5602 (
            .O(N__27234),
            .I(N__27213));
    IoSpan4Mux I__5601 (
            .O(N__27231),
            .I(N__27210));
    Span4Mux_v I__5600 (
            .O(N__27228),
            .I(N__27207));
    Span4Mux_h I__5599 (
            .O(N__27223),
            .I(N__27204));
    IoSpan4Mux I__5598 (
            .O(N__27216),
            .I(N__27201));
    Span4Mux_h I__5597 (
            .O(N__27213),
            .I(N__27198));
    Odrv4 I__5596 (
            .O(N__27210),
            .I(slp_s3n));
    Odrv4 I__5595 (
            .O(N__27207),
            .I(slp_s3n));
    Odrv4 I__5594 (
            .O(N__27204),
            .I(slp_s3n));
    Odrv4 I__5593 (
            .O(N__27201),
            .I(slp_s3n));
    Odrv4 I__5592 (
            .O(N__27198),
            .I(slp_s3n));
    CascadeMux I__5591 (
            .O(N__27187),
            .I(\POWERLED.un1_clk_100khz_51_and_i_a2_6_0_cascade_ ));
    CascadeMux I__5590 (
            .O(N__27184),
            .I(\POWERLED.un1_clk_100khz_51_and_i_a2_6_sx_cascade_ ));
    CascadeMux I__5589 (
            .O(N__27181),
            .I(\POWERLED.func_state_RNIPUGO_0Z0Z_1_cascade_ ));
    InMux I__5588 (
            .O(N__27178),
            .I(N__27175));
    LocalMux I__5587 (
            .O(N__27175),
            .I(\POWERLED.N_309_N ));
    InMux I__5586 (
            .O(N__27172),
            .I(N__27169));
    LocalMux I__5585 (
            .O(N__27169),
            .I(\POWERLED.count_clk_RNI2O4A1Z0Z_10 ));
    CascadeMux I__5584 (
            .O(N__27166),
            .I(\POWERLED.un1_clk_100khz_51_and_i_o2_4_1_cascade_ ));
    InMux I__5583 (
            .O(N__27163),
            .I(N__27155));
    InMux I__5582 (
            .O(N__27162),
            .I(N__27155));
    InMux I__5581 (
            .O(N__27161),
            .I(N__27146));
    InMux I__5580 (
            .O(N__27160),
            .I(N__27146));
    LocalMux I__5579 (
            .O(N__27155),
            .I(N__27137));
    InMux I__5578 (
            .O(N__27154),
            .I(N__27134));
    InMux I__5577 (
            .O(N__27153),
            .I(N__27129));
    InMux I__5576 (
            .O(N__27152),
            .I(N__27129));
    InMux I__5575 (
            .O(N__27151),
            .I(N__27126));
    LocalMux I__5574 (
            .O(N__27146),
            .I(N__27123));
    CascadeMux I__5573 (
            .O(N__27145),
            .I(N__27120));
    CascadeMux I__5572 (
            .O(N__27144),
            .I(N__27114));
    CascadeMux I__5571 (
            .O(N__27143),
            .I(N__27111));
    InMux I__5570 (
            .O(N__27142),
            .I(N__27105));
    InMux I__5569 (
            .O(N__27141),
            .I(N__27105));
    InMux I__5568 (
            .O(N__27140),
            .I(N__27102));
    Span4Mux_h I__5567 (
            .O(N__27137),
            .I(N__27097));
    LocalMux I__5566 (
            .O(N__27134),
            .I(N__27097));
    LocalMux I__5565 (
            .O(N__27129),
            .I(N__27094));
    LocalMux I__5564 (
            .O(N__27126),
            .I(N__27089));
    Span4Mux_v I__5563 (
            .O(N__27123),
            .I(N__27089));
    InMux I__5562 (
            .O(N__27120),
            .I(N__27086));
    InMux I__5561 (
            .O(N__27119),
            .I(N__27079));
    InMux I__5560 (
            .O(N__27118),
            .I(N__27079));
    InMux I__5559 (
            .O(N__27117),
            .I(N__27079));
    InMux I__5558 (
            .O(N__27114),
            .I(N__27073));
    InMux I__5557 (
            .O(N__27111),
            .I(N__27073));
    InMux I__5556 (
            .O(N__27110),
            .I(N__27070));
    LocalMux I__5555 (
            .O(N__27105),
            .I(N__27066));
    LocalMux I__5554 (
            .O(N__27102),
            .I(N__27055));
    Span4Mux_v I__5553 (
            .O(N__27097),
            .I(N__27055));
    Span4Mux_h I__5552 (
            .O(N__27094),
            .I(N__27055));
    Span4Mux_h I__5551 (
            .O(N__27089),
            .I(N__27055));
    LocalMux I__5550 (
            .O(N__27086),
            .I(N__27055));
    LocalMux I__5549 (
            .O(N__27079),
            .I(N__27050));
    CascadeMux I__5548 (
            .O(N__27078),
            .I(N__27047));
    LocalMux I__5547 (
            .O(N__27073),
            .I(N__27044));
    LocalMux I__5546 (
            .O(N__27070),
            .I(N__27041));
    InMux I__5545 (
            .O(N__27069),
            .I(N__27038));
    Span4Mux_h I__5544 (
            .O(N__27066),
            .I(N__27035));
    Span4Mux_v I__5543 (
            .O(N__27055),
            .I(N__27032));
    InMux I__5542 (
            .O(N__27054),
            .I(N__27027));
    InMux I__5541 (
            .O(N__27053),
            .I(N__27027));
    Span12Mux_s6_h I__5540 (
            .O(N__27050),
            .I(N__27024));
    InMux I__5539 (
            .O(N__27047),
            .I(N__27021));
    Span4Mux_v I__5538 (
            .O(N__27044),
            .I(N__27014));
    Span4Mux_v I__5537 (
            .O(N__27041),
            .I(N__27014));
    LocalMux I__5536 (
            .O(N__27038),
            .I(N__27014));
    Odrv4 I__5535 (
            .O(N__27035),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__5534 (
            .O(N__27032),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__5533 (
            .O(N__27027),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv12 I__5532 (
            .O(N__27024),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__5531 (
            .O(N__27021),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__5530 (
            .O(N__27014),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    InMux I__5529 (
            .O(N__27001),
            .I(N__26998));
    LocalMux I__5528 (
            .O(N__26998),
            .I(N__26995));
    Odrv12 I__5527 (
            .O(N__26995),
            .I(\POWERLED.N_145_N ));
    InMux I__5526 (
            .O(N__26992),
            .I(N__26989));
    LocalMux I__5525 (
            .O(N__26989),
            .I(\POWERLED.un1_clk_100khz_51_and_i_a2_5_0 ));
    CascadeMux I__5524 (
            .O(N__26986),
            .I(\POWERLED.un1_clk_100khz_51_and_i_a2_5_0_cascade_ ));
    InMux I__5523 (
            .O(N__26983),
            .I(N__26974));
    InMux I__5522 (
            .O(N__26982),
            .I(N__26974));
    InMux I__5521 (
            .O(N__26981),
            .I(N__26974));
    LocalMux I__5520 (
            .O(N__26974),
            .I(N__26971));
    Span4Mux_v I__5519 (
            .O(N__26971),
            .I(N__26966));
    InMux I__5518 (
            .O(N__26970),
            .I(N__26963));
    InMux I__5517 (
            .O(N__26969),
            .I(N__26960));
    Odrv4 I__5516 (
            .O(N__26966),
            .I(RSMRSTn_fast));
    LocalMux I__5515 (
            .O(N__26963),
            .I(RSMRSTn_fast));
    LocalMux I__5514 (
            .O(N__26960),
            .I(RSMRSTn_fast));
    InMux I__5513 (
            .O(N__26953),
            .I(N__26950));
    LocalMux I__5512 (
            .O(N__26950),
            .I(\POWERLED.func_state_RNIPUGOZ0Z_1 ));
    CascadeMux I__5511 (
            .O(N__26947),
            .I(N__26943));
    InMux I__5510 (
            .O(N__26946),
            .I(N__26939));
    InMux I__5509 (
            .O(N__26943),
            .I(N__26934));
    InMux I__5508 (
            .O(N__26942),
            .I(N__26934));
    LocalMux I__5507 (
            .O(N__26939),
            .I(\POWERLED.N_340 ));
    LocalMux I__5506 (
            .O(N__26934),
            .I(\POWERLED.N_340 ));
    CascadeMux I__5505 (
            .O(N__26929),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_ ));
    InMux I__5504 (
            .O(N__26926),
            .I(N__26923));
    LocalMux I__5503 (
            .O(N__26923),
            .I(\POWERLED.N_284 ));
    InMux I__5502 (
            .O(N__26920),
            .I(N__26896));
    InMux I__5501 (
            .O(N__26919),
            .I(N__26896));
    InMux I__5500 (
            .O(N__26918),
            .I(N__26896));
    InMux I__5499 (
            .O(N__26917),
            .I(N__26896));
    InMux I__5498 (
            .O(N__26916),
            .I(N__26887));
    InMux I__5497 (
            .O(N__26915),
            .I(N__26887));
    InMux I__5496 (
            .O(N__26914),
            .I(N__26887));
    InMux I__5495 (
            .O(N__26913),
            .I(N__26887));
    InMux I__5494 (
            .O(N__26912),
            .I(N__26880));
    InMux I__5493 (
            .O(N__26911),
            .I(N__26880));
    InMux I__5492 (
            .O(N__26910),
            .I(N__26880));
    InMux I__5491 (
            .O(N__26909),
            .I(N__26875));
    InMux I__5490 (
            .O(N__26908),
            .I(N__26875));
    InMux I__5489 (
            .O(N__26907),
            .I(N__26868));
    InMux I__5488 (
            .O(N__26906),
            .I(N__26868));
    InMux I__5487 (
            .O(N__26905),
            .I(N__26868));
    LocalMux I__5486 (
            .O(N__26896),
            .I(N__26865));
    LocalMux I__5485 (
            .O(N__26887),
            .I(N__26856));
    LocalMux I__5484 (
            .O(N__26880),
            .I(N__26856));
    LocalMux I__5483 (
            .O(N__26875),
            .I(N__26853));
    LocalMux I__5482 (
            .O(N__26868),
            .I(N__26848));
    Span4Mux_h I__5481 (
            .O(N__26865),
            .I(N__26848));
    InMux I__5480 (
            .O(N__26864),
            .I(N__26839));
    InMux I__5479 (
            .O(N__26863),
            .I(N__26839));
    InMux I__5478 (
            .O(N__26862),
            .I(N__26839));
    InMux I__5477 (
            .O(N__26861),
            .I(N__26839));
    Span4Mux_v I__5476 (
            .O(N__26856),
            .I(N__26836));
    Span4Mux_h I__5475 (
            .O(N__26853),
            .I(N__26833));
    Span4Mux_h I__5474 (
            .O(N__26848),
            .I(N__26828));
    LocalMux I__5473 (
            .O(N__26839),
            .I(N__26828));
    Span4Mux_h I__5472 (
            .O(N__26836),
            .I(N__26825));
    Span4Mux_v I__5471 (
            .O(N__26833),
            .I(N__26820));
    Span4Mux_v I__5470 (
            .O(N__26828),
            .I(N__26820));
    Odrv4 I__5469 (
            .O(N__26825),
            .I(\POWERLED.func_state_RNIBQDB2Z0Z_0 ));
    Odrv4 I__5468 (
            .O(N__26820),
            .I(\POWERLED.func_state_RNIBQDB2Z0Z_0 ));
    InMux I__5467 (
            .O(N__26815),
            .I(N__26809));
    InMux I__5466 (
            .O(N__26814),
            .I(N__26809));
    LocalMux I__5465 (
            .O(N__26809),
            .I(N__26806));
    Odrv4 I__5464 (
            .O(N__26806),
            .I(\POWERLED.N_340_N ));
    InMux I__5463 (
            .O(N__26803),
            .I(N__26799));
    CascadeMux I__5462 (
            .O(N__26802),
            .I(N__26796));
    LocalMux I__5461 (
            .O(N__26799),
            .I(N__26793));
    InMux I__5460 (
            .O(N__26796),
            .I(N__26790));
    Odrv4 I__5459 (
            .O(N__26793),
            .I(\POWERLED.func_state_RNI_1Z0Z_0 ));
    LocalMux I__5458 (
            .O(N__26790),
            .I(\POWERLED.func_state_RNI_1Z0Z_0 ));
    InMux I__5457 (
            .O(N__26785),
            .I(N__26782));
    LocalMux I__5456 (
            .O(N__26782),
            .I(\POWERLED.un1_func_state25_6_0_o_N_294_N ));
    InMux I__5455 (
            .O(N__26779),
            .I(N__26776));
    LocalMux I__5454 (
            .O(N__26776),
            .I(N__26773));
    Odrv12 I__5453 (
            .O(N__26773),
            .I(\POWERLED.func_state_1_m2_am_1_1 ));
    InMux I__5452 (
            .O(N__26770),
            .I(N__26760));
    InMux I__5451 (
            .O(N__26769),
            .I(N__26760));
    CascadeMux I__5450 (
            .O(N__26768),
            .I(N__26756));
    InMux I__5449 (
            .O(N__26767),
            .I(N__26752));
    InMux I__5448 (
            .O(N__26766),
            .I(N__26749));
    InMux I__5447 (
            .O(N__26765),
            .I(N__26746));
    LocalMux I__5446 (
            .O(N__26760),
            .I(N__26743));
    CascadeMux I__5445 (
            .O(N__26759),
            .I(N__26738));
    InMux I__5444 (
            .O(N__26756),
            .I(N__26733));
    InMux I__5443 (
            .O(N__26755),
            .I(N__26733));
    LocalMux I__5442 (
            .O(N__26752),
            .I(N__26728));
    LocalMux I__5441 (
            .O(N__26749),
            .I(N__26728));
    LocalMux I__5440 (
            .O(N__26746),
            .I(N__26725));
    Span4Mux_v I__5439 (
            .O(N__26743),
            .I(N__26722));
    InMux I__5438 (
            .O(N__26742),
            .I(N__26717));
    InMux I__5437 (
            .O(N__26741),
            .I(N__26717));
    InMux I__5436 (
            .O(N__26738),
            .I(N__26712));
    LocalMux I__5435 (
            .O(N__26733),
            .I(N__26701));
    Span4Mux_v I__5434 (
            .O(N__26728),
            .I(N__26701));
    Span4Mux_v I__5433 (
            .O(N__26725),
            .I(N__26701));
    Span4Mux_h I__5432 (
            .O(N__26722),
            .I(N__26701));
    LocalMux I__5431 (
            .O(N__26717),
            .I(N__26701));
    InMux I__5430 (
            .O(N__26716),
            .I(N__26695));
    InMux I__5429 (
            .O(N__26715),
            .I(N__26695));
    LocalMux I__5428 (
            .O(N__26712),
            .I(N__26686));
    Span4Mux_h I__5427 (
            .O(N__26701),
            .I(N__26683));
    InMux I__5426 (
            .O(N__26700),
            .I(N__26679));
    LocalMux I__5425 (
            .O(N__26695),
            .I(N__26674));
    InMux I__5424 (
            .O(N__26694),
            .I(N__26667));
    InMux I__5423 (
            .O(N__26693),
            .I(N__26667));
    InMux I__5422 (
            .O(N__26692),
            .I(N__26667));
    InMux I__5421 (
            .O(N__26691),
            .I(N__26660));
    InMux I__5420 (
            .O(N__26690),
            .I(N__26660));
    InMux I__5419 (
            .O(N__26689),
            .I(N__26660));
    Span4Mux_v I__5418 (
            .O(N__26686),
            .I(N__26655));
    Span4Mux_s3_h I__5417 (
            .O(N__26683),
            .I(N__26655));
    InMux I__5416 (
            .O(N__26682),
            .I(N__26652));
    LocalMux I__5415 (
            .O(N__26679),
            .I(N__26649));
    InMux I__5414 (
            .O(N__26678),
            .I(N__26644));
    InMux I__5413 (
            .O(N__26677),
            .I(N__26644));
    Sp12to4 I__5412 (
            .O(N__26674),
            .I(N__26639));
    LocalMux I__5411 (
            .O(N__26667),
            .I(N__26639));
    LocalMux I__5410 (
            .O(N__26660),
            .I(\POWERLED.func_N_5_mux_0 ));
    Odrv4 I__5409 (
            .O(N__26655),
            .I(\POWERLED.func_N_5_mux_0 ));
    LocalMux I__5408 (
            .O(N__26652),
            .I(\POWERLED.func_N_5_mux_0 ));
    Odrv12 I__5407 (
            .O(N__26649),
            .I(\POWERLED.func_N_5_mux_0 ));
    LocalMux I__5406 (
            .O(N__26644),
            .I(\POWERLED.func_N_5_mux_0 ));
    Odrv12 I__5405 (
            .O(N__26639),
            .I(\POWERLED.func_N_5_mux_0 ));
    InMux I__5404 (
            .O(N__26626),
            .I(N__26623));
    LocalMux I__5403 (
            .O(N__26623),
            .I(N__26620));
    Odrv12 I__5402 (
            .O(N__26620),
            .I(\POWERLED.func_state_RNIBL3Q3Z0Z_1 ));
    InMux I__5401 (
            .O(N__26617),
            .I(N__26614));
    LocalMux I__5400 (
            .O(N__26614),
            .I(N__26611));
    Span4Mux_v I__5399 (
            .O(N__26611),
            .I(N__26608));
    Odrv4 I__5398 (
            .O(N__26608),
            .I(\POWERLED.func_state_1_m2s2_i_a2_0_0 ));
    CascadeMux I__5397 (
            .O(N__26605),
            .I(N__26596));
    InMux I__5396 (
            .O(N__26604),
            .I(N__26591));
    InMux I__5395 (
            .O(N__26603),
            .I(N__26588));
    InMux I__5394 (
            .O(N__26602),
            .I(N__26583));
    InMux I__5393 (
            .O(N__26601),
            .I(N__26583));
    CascadeMux I__5392 (
            .O(N__26600),
            .I(N__26580));
    InMux I__5391 (
            .O(N__26599),
            .I(N__26571));
    InMux I__5390 (
            .O(N__26596),
            .I(N__26566));
    InMux I__5389 (
            .O(N__26595),
            .I(N__26566));
    InMux I__5388 (
            .O(N__26594),
            .I(N__26563));
    LocalMux I__5387 (
            .O(N__26591),
            .I(N__26560));
    LocalMux I__5386 (
            .O(N__26588),
            .I(N__26555));
    LocalMux I__5385 (
            .O(N__26583),
            .I(N__26555));
    InMux I__5384 (
            .O(N__26580),
            .I(N__26552));
    InMux I__5383 (
            .O(N__26579),
            .I(N__26549));
    InMux I__5382 (
            .O(N__26578),
            .I(N__26546));
    InMux I__5381 (
            .O(N__26577),
            .I(N__26540));
    InMux I__5380 (
            .O(N__26576),
            .I(N__26540));
    InMux I__5379 (
            .O(N__26575),
            .I(N__26535));
    InMux I__5378 (
            .O(N__26574),
            .I(N__26535));
    LocalMux I__5377 (
            .O(N__26571),
            .I(N__26532));
    LocalMux I__5376 (
            .O(N__26566),
            .I(N__26527));
    LocalMux I__5375 (
            .O(N__26563),
            .I(N__26527));
    Span4Mux_s3_h I__5374 (
            .O(N__26560),
            .I(N__26522));
    Span4Mux_v I__5373 (
            .O(N__26555),
            .I(N__26522));
    LocalMux I__5372 (
            .O(N__26552),
            .I(N__26517));
    LocalMux I__5371 (
            .O(N__26549),
            .I(N__26517));
    LocalMux I__5370 (
            .O(N__26546),
            .I(N__26513));
    InMux I__5369 (
            .O(N__26545),
            .I(N__26510));
    LocalMux I__5368 (
            .O(N__26540),
            .I(N__26505));
    LocalMux I__5367 (
            .O(N__26535),
            .I(N__26505));
    Span12Mux_s10_v I__5366 (
            .O(N__26532),
            .I(N__26502));
    Span4Mux_v I__5365 (
            .O(N__26527),
            .I(N__26499));
    Span4Mux_h I__5364 (
            .O(N__26522),
            .I(N__26494));
    Span4Mux_v I__5363 (
            .O(N__26517),
            .I(N__26494));
    InMux I__5362 (
            .O(N__26516),
            .I(N__26491));
    Odrv4 I__5361 (
            .O(N__26513),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__5360 (
            .O(N__26510),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5359 (
            .O(N__26505),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv12 I__5358 (
            .O(N__26502),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5357 (
            .O(N__26499),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5356 (
            .O(N__26494),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__5355 (
            .O(N__26491),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    InMux I__5354 (
            .O(N__26476),
            .I(N__26471));
    InMux I__5353 (
            .O(N__26475),
            .I(N__26463));
    InMux I__5352 (
            .O(N__26474),
            .I(N__26463));
    LocalMux I__5351 (
            .O(N__26471),
            .I(N__26460));
    InMux I__5350 (
            .O(N__26470),
            .I(N__26457));
    InMux I__5349 (
            .O(N__26469),
            .I(N__26451));
    InMux I__5348 (
            .O(N__26468),
            .I(N__26451));
    LocalMux I__5347 (
            .O(N__26463),
            .I(N__26448));
    Span4Mux_v I__5346 (
            .O(N__26460),
            .I(N__26445));
    LocalMux I__5345 (
            .O(N__26457),
            .I(N__26442));
    InMux I__5344 (
            .O(N__26456),
            .I(N__26439));
    LocalMux I__5343 (
            .O(N__26451),
            .I(N__26432));
    Span4Mux_v I__5342 (
            .O(N__26448),
            .I(N__26432));
    Span4Mux_v I__5341 (
            .O(N__26445),
            .I(N__26432));
    Span4Mux_h I__5340 (
            .O(N__26442),
            .I(N__26427));
    LocalMux I__5339 (
            .O(N__26439),
            .I(N__26427));
    Odrv4 I__5338 (
            .O(N__26432),
            .I(func_state_RNI_7_1));
    Odrv4 I__5337 (
            .O(N__26427),
            .I(func_state_RNI_7_1));
    InMux I__5336 (
            .O(N__26422),
            .I(N__26419));
    LocalMux I__5335 (
            .O(N__26419),
            .I(N__26416));
    Odrv4 I__5334 (
            .O(N__26416),
            .I(N_7));
    IoInMux I__5333 (
            .O(N__26413),
            .I(N__26408));
    InMux I__5332 (
            .O(N__26412),
            .I(N__26405));
    CascadeMux I__5331 (
            .O(N__26411),
            .I(N__26401));
    LocalMux I__5330 (
            .O(N__26408),
            .I(N__26398));
    LocalMux I__5329 (
            .O(N__26405),
            .I(N__26394));
    InMux I__5328 (
            .O(N__26404),
            .I(N__26391));
    InMux I__5327 (
            .O(N__26401),
            .I(N__26388));
    IoSpan4Mux I__5326 (
            .O(N__26398),
            .I(N__26383));
    InMux I__5325 (
            .O(N__26397),
            .I(N__26380));
    Span4Mux_h I__5324 (
            .O(N__26394),
            .I(N__26373));
    LocalMux I__5323 (
            .O(N__26391),
            .I(N__26373));
    LocalMux I__5322 (
            .O(N__26388),
            .I(N__26373));
    InMux I__5321 (
            .O(N__26387),
            .I(N__26370));
    InMux I__5320 (
            .O(N__26386),
            .I(N__26367));
    Span4Mux_s1_v I__5319 (
            .O(N__26383),
            .I(N__26362));
    LocalMux I__5318 (
            .O(N__26380),
            .I(N__26362));
    Span4Mux_h I__5317 (
            .O(N__26373),
            .I(N__26359));
    LocalMux I__5316 (
            .O(N__26370),
            .I(N__26356));
    LocalMux I__5315 (
            .O(N__26367),
            .I(N__26348));
    Span4Mux_h I__5314 (
            .O(N__26362),
            .I(N__26341));
    Span4Mux_s3_h I__5313 (
            .O(N__26359),
            .I(N__26341));
    Span4Mux_s1_v I__5312 (
            .O(N__26356),
            .I(N__26341));
    InMux I__5311 (
            .O(N__26355),
            .I(N__26338));
    InMux I__5310 (
            .O(N__26354),
            .I(N__26333));
    InMux I__5309 (
            .O(N__26353),
            .I(N__26333));
    InMux I__5308 (
            .O(N__26352),
            .I(N__26328));
    InMux I__5307 (
            .O(N__26351),
            .I(N__26328));
    Span4Mux_h I__5306 (
            .O(N__26348),
            .I(N__26325));
    Sp12to4 I__5305 (
            .O(N__26341),
            .I(N__26318));
    LocalMux I__5304 (
            .O(N__26338),
            .I(N__26318));
    LocalMux I__5303 (
            .O(N__26333),
            .I(N__26318));
    LocalMux I__5302 (
            .O(N__26328),
            .I(rsmrstn));
    Odrv4 I__5301 (
            .O(N__26325),
            .I(rsmrstn));
    Odrv12 I__5300 (
            .O(N__26318),
            .I(rsmrstn));
    CascadeMux I__5299 (
            .O(N__26311),
            .I(G_34_0_a4_0_2_cascade_));
    CascadeMux I__5298 (
            .O(N__26308),
            .I(N__26305));
    InMux I__5297 (
            .O(N__26305),
            .I(N__26299));
    InMux I__5296 (
            .O(N__26304),
            .I(N__26299));
    LocalMux I__5295 (
            .O(N__26299),
            .I(POWERLED_un1_dutycycle_172_m3_0_0));
    InMux I__5294 (
            .O(N__26296),
            .I(N__26290));
    InMux I__5293 (
            .O(N__26295),
            .I(N__26290));
    LocalMux I__5292 (
            .O(N__26290),
            .I(\POWERLED.N_8_0 ));
    InMux I__5291 (
            .O(N__26287),
            .I(N__26282));
    InMux I__5290 (
            .O(N__26286),
            .I(N__26277));
    InMux I__5289 (
            .O(N__26285),
            .I(N__26277));
    LocalMux I__5288 (
            .O(N__26282),
            .I(N__26274));
    LocalMux I__5287 (
            .O(N__26277),
            .I(N__26271));
    Span4Mux_h I__5286 (
            .O(N__26274),
            .I(N__26268));
    Odrv4 I__5285 (
            .O(N__26271),
            .I(\POWERLED.un1_dutycycle_172_m1_ns_1 ));
    Odrv4 I__5284 (
            .O(N__26268),
            .I(\POWERLED.un1_dutycycle_172_m1_ns_1 ));
    CascadeMux I__5283 (
            .O(N__26263),
            .I(N__26260));
    InMux I__5282 (
            .O(N__26260),
            .I(N__26254));
    InMux I__5281 (
            .O(N__26259),
            .I(N__26254));
    LocalMux I__5280 (
            .O(N__26254),
            .I(N__26251));
    Span4Mux_v I__5279 (
            .O(N__26251),
            .I(N__26246));
    InMux I__5278 (
            .O(N__26250),
            .I(N__26243));
    CascadeMux I__5277 (
            .O(N__26249),
            .I(N__26240));
    Sp12to4 I__5276 (
            .O(N__26246),
            .I(N__26234));
    LocalMux I__5275 (
            .O(N__26243),
            .I(N__26234));
    InMux I__5274 (
            .O(N__26240),
            .I(N__26231));
    InMux I__5273 (
            .O(N__26239),
            .I(N__26228));
    Span12Mux_s5_h I__5272 (
            .O(N__26234),
            .I(N__26223));
    LocalMux I__5271 (
            .O(N__26231),
            .I(N__26223));
    LocalMux I__5270 (
            .O(N__26228),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_3 ));
    Odrv12 I__5269 (
            .O(N__26223),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_3 ));
    InMux I__5268 (
            .O(N__26218),
            .I(N__26215));
    LocalMux I__5267 (
            .O(N__26215),
            .I(N_11));
    InMux I__5266 (
            .O(N__26212),
            .I(N__26206));
    InMux I__5265 (
            .O(N__26211),
            .I(N__26203));
    InMux I__5264 (
            .O(N__26210),
            .I(N__26200));
    InMux I__5263 (
            .O(N__26209),
            .I(N__26196));
    LocalMux I__5262 (
            .O(N__26206),
            .I(N__26193));
    LocalMux I__5261 (
            .O(N__26203),
            .I(N__26190));
    LocalMux I__5260 (
            .O(N__26200),
            .I(N__26187));
    InMux I__5259 (
            .O(N__26199),
            .I(N__26184));
    LocalMux I__5258 (
            .O(N__26196),
            .I(N__26181));
    Span4Mux_h I__5257 (
            .O(N__26193),
            .I(N__26178));
    Span12Mux_s10_v I__5256 (
            .O(N__26190),
            .I(N__26175));
    Odrv12 I__5255 (
            .O(N__26187),
            .I(\POWERLED.N_319_0 ));
    LocalMux I__5254 (
            .O(N__26184),
            .I(\POWERLED.N_319_0 ));
    Odrv4 I__5253 (
            .O(N__26181),
            .I(\POWERLED.N_319_0 ));
    Odrv4 I__5252 (
            .O(N__26178),
            .I(\POWERLED.N_319_0 ));
    Odrv12 I__5251 (
            .O(N__26175),
            .I(\POWERLED.N_319_0 ));
    InMux I__5250 (
            .O(N__26164),
            .I(N__26158));
    InMux I__5249 (
            .O(N__26163),
            .I(N__26158));
    LocalMux I__5248 (
            .O(N__26158),
            .I(N__26152));
    CascadeMux I__5247 (
            .O(N__26157),
            .I(N__26148));
    CascadeMux I__5246 (
            .O(N__26156),
            .I(N__26144));
    InMux I__5245 (
            .O(N__26155),
            .I(N__26141));
    Span4Mux_v I__5244 (
            .O(N__26152),
            .I(N__26138));
    InMux I__5243 (
            .O(N__26151),
            .I(N__26135));
    InMux I__5242 (
            .O(N__26148),
            .I(N__26130));
    InMux I__5241 (
            .O(N__26147),
            .I(N__26130));
    InMux I__5240 (
            .O(N__26144),
            .I(N__26127));
    LocalMux I__5239 (
            .O(N__26141),
            .I(N__26124));
    Odrv4 I__5238 (
            .O(N__26138),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__5237 (
            .O(N__26135),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__5236 (
            .O(N__26130),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__5235 (
            .O(N__26127),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv12 I__5234 (
            .O(N__26124),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__5233 (
            .O(N__26113),
            .I(N__26110));
    LocalMux I__5232 (
            .O(N__26110),
            .I(\POWERLED.N_297 ));
    InMux I__5231 (
            .O(N__26107),
            .I(N__26104));
    LocalMux I__5230 (
            .O(N__26104),
            .I(N__26101));
    Odrv4 I__5229 (
            .O(N__26101),
            .I(\POWERLED.un1_func_state25_6_0_a2_1 ));
    CascadeMux I__5228 (
            .O(N__26098),
            .I(\POWERLED.un1_func_state25_6_0_o_N_296_N_cascade_ ));
    CascadeMux I__5227 (
            .O(N__26095),
            .I(\POWERLED.un1_func_state25_6_0_1_cascade_ ));
    CascadeMux I__5226 (
            .O(N__26092),
            .I(N__26089));
    InMux I__5225 (
            .O(N__26089),
            .I(N__26086));
    LocalMux I__5224 (
            .O(N__26086),
            .I(N__26083));
    Span4Mux_h I__5223 (
            .O(N__26083),
            .I(N__26080));
    Span4Mux_v I__5222 (
            .O(N__26080),
            .I(N__26077));
    Odrv4 I__5221 (
            .O(N__26077),
            .I(\POWERLED.un1_func_state25_6_0_2 ));
    InMux I__5220 (
            .O(N__26074),
            .I(N__26071));
    LocalMux I__5219 (
            .O(N__26071),
            .I(N__26065));
    InMux I__5218 (
            .O(N__26070),
            .I(N__26060));
    InMux I__5217 (
            .O(N__26069),
            .I(N__26060));
    InMux I__5216 (
            .O(N__26068),
            .I(N__26057));
    Odrv12 I__5215 (
            .O(N__26065),
            .I(RSMRSTn_rep1));
    LocalMux I__5214 (
            .O(N__26060),
            .I(RSMRSTn_rep1));
    LocalMux I__5213 (
            .O(N__26057),
            .I(RSMRSTn_rep1));
    InMux I__5212 (
            .O(N__26050),
            .I(N__26043));
    InMux I__5211 (
            .O(N__26049),
            .I(N__26038));
    InMux I__5210 (
            .O(N__26048),
            .I(N__26038));
    InMux I__5209 (
            .O(N__26047),
            .I(N__26031));
    InMux I__5208 (
            .O(N__26046),
            .I(N__26031));
    LocalMux I__5207 (
            .O(N__26043),
            .I(N__26026));
    LocalMux I__5206 (
            .O(N__26038),
            .I(N__26026));
    InMux I__5205 (
            .O(N__26037),
            .I(N__26021));
    InMux I__5204 (
            .O(N__26036),
            .I(N__26021));
    LocalMux I__5203 (
            .O(N__26031),
            .I(N__26018));
    Span4Mux_v I__5202 (
            .O(N__26026),
            .I(N__26013));
    LocalMux I__5201 (
            .O(N__26021),
            .I(N__26013));
    Span4Mux_h I__5200 (
            .O(N__26018),
            .I(N__26010));
    Span4Mux_h I__5199 (
            .O(N__26013),
            .I(N__26007));
    Odrv4 I__5198 (
            .O(N__26010),
            .I(\POWERLED.N_4_0_3 ));
    Odrv4 I__5197 (
            .O(N__26007),
            .I(\POWERLED.N_4_0_3 ));
    InMux I__5196 (
            .O(N__26002),
            .I(N__25998));
    CascadeMux I__5195 (
            .O(N__26001),
            .I(N__25993));
    LocalMux I__5194 (
            .O(N__25998),
            .I(N__25990));
    InMux I__5193 (
            .O(N__25997),
            .I(N__25987));
    InMux I__5192 (
            .O(N__25996),
            .I(N__25984));
    InMux I__5191 (
            .O(N__25993),
            .I(N__25981));
    Span4Mux_v I__5190 (
            .O(N__25990),
            .I(N__25978));
    LocalMux I__5189 (
            .O(N__25987),
            .I(N__25975));
    LocalMux I__5188 (
            .O(N__25984),
            .I(N__25970));
    LocalMux I__5187 (
            .O(N__25981),
            .I(N__25970));
    Odrv4 I__5186 (
            .O(N__25978),
            .I(\POWERLED.func_state_RNIOGRSZ0Z_0 ));
    Odrv4 I__5185 (
            .O(N__25975),
            .I(\POWERLED.func_state_RNIOGRSZ0Z_0 ));
    Odrv4 I__5184 (
            .O(N__25970),
            .I(\POWERLED.func_state_RNIOGRSZ0Z_0 ));
    CascadeMux I__5183 (
            .O(N__25963),
            .I(N__25959));
    CascadeMux I__5182 (
            .O(N__25962),
            .I(N__25956));
    InMux I__5181 (
            .O(N__25959),
            .I(N__25953));
    InMux I__5180 (
            .O(N__25956),
            .I(N__25950));
    LocalMux I__5179 (
            .O(N__25953),
            .I(N__25947));
    LocalMux I__5178 (
            .O(N__25950),
            .I(N__25942));
    Span4Mux_h I__5177 (
            .O(N__25947),
            .I(N__25942));
    Odrv4 I__5176 (
            .O(N__25942),
            .I(\POWERLED.func_state_1_ss0_i_0_o2_1 ));
    InMux I__5175 (
            .O(N__25939),
            .I(N__25935));
    InMux I__5174 (
            .O(N__25938),
            .I(N__25932));
    LocalMux I__5173 (
            .O(N__25935),
            .I(N__25927));
    LocalMux I__5172 (
            .O(N__25932),
            .I(N__25927));
    Odrv4 I__5171 (
            .O(N__25927),
            .I(\POWERLED.N_76 ));
    CascadeMux I__5170 (
            .O(N__25924),
            .I(\POWERLED.func_state_RNI91IA4Z0Z_1_cascade_ ));
    InMux I__5169 (
            .O(N__25921),
            .I(N__25918));
    LocalMux I__5168 (
            .O(N__25918),
            .I(\POWERLED.func_state_1_m2_1 ));
    InMux I__5167 (
            .O(N__25915),
            .I(N__25909));
    InMux I__5166 (
            .O(N__25914),
            .I(N__25909));
    LocalMux I__5165 (
            .O(N__25909),
            .I(\POWERLED.func_stateZ0Z_1 ));
    CascadeMux I__5164 (
            .O(N__25906),
            .I(\POWERLED.func_state_1_m2_1_cascade_ ));
    CascadeMux I__5163 (
            .O(N__25903),
            .I(N__25900));
    InMux I__5162 (
            .O(N__25900),
            .I(N__25897));
    LocalMux I__5161 (
            .O(N__25897),
            .I(N__25891));
    InMux I__5160 (
            .O(N__25896),
            .I(N__25888));
    InMux I__5159 (
            .O(N__25895),
            .I(N__25883));
    InMux I__5158 (
            .O(N__25894),
            .I(N__25883));
    Span4Mux_h I__5157 (
            .O(N__25891),
            .I(N__25876));
    LocalMux I__5156 (
            .O(N__25888),
            .I(N__25876));
    LocalMux I__5155 (
            .O(N__25883),
            .I(N__25876));
    Odrv4 I__5154 (
            .O(N__25876),
            .I(\POWERLED.func_state_enZ0 ));
    CascadeMux I__5153 (
            .O(N__25873),
            .I(N__25869));
    CascadeMux I__5152 (
            .O(N__25872),
            .I(N__25866));
    InMux I__5151 (
            .O(N__25869),
            .I(N__25857));
    InMux I__5150 (
            .O(N__25866),
            .I(N__25854));
    InMux I__5149 (
            .O(N__25865),
            .I(N__25849));
    InMux I__5148 (
            .O(N__25864),
            .I(N__25849));
    InMux I__5147 (
            .O(N__25863),
            .I(N__25843));
    InMux I__5146 (
            .O(N__25862),
            .I(N__25843));
    InMux I__5145 (
            .O(N__25861),
            .I(N__25840));
    InMux I__5144 (
            .O(N__25860),
            .I(N__25837));
    LocalMux I__5143 (
            .O(N__25857),
            .I(N__25830));
    LocalMux I__5142 (
            .O(N__25854),
            .I(N__25830));
    LocalMux I__5141 (
            .O(N__25849),
            .I(N__25830));
    InMux I__5140 (
            .O(N__25848),
            .I(N__25827));
    LocalMux I__5139 (
            .O(N__25843),
            .I(N__25824));
    LocalMux I__5138 (
            .O(N__25840),
            .I(N__25821));
    LocalMux I__5137 (
            .O(N__25837),
            .I(N__25818));
    Span4Mux_v I__5136 (
            .O(N__25830),
            .I(N__25814));
    LocalMux I__5135 (
            .O(N__25827),
            .I(N__25809));
    Span4Mux_h I__5134 (
            .O(N__25824),
            .I(N__25809));
    Span4Mux_h I__5133 (
            .O(N__25821),
            .I(N__25804));
    Span4Mux_v I__5132 (
            .O(N__25818),
            .I(N__25804));
    InMux I__5131 (
            .O(N__25817),
            .I(N__25801));
    Odrv4 I__5130 (
            .O(N__25814),
            .I(\POWERLED.un1_N_3_mux_0 ));
    Odrv4 I__5129 (
            .O(N__25809),
            .I(\POWERLED.un1_N_3_mux_0 ));
    Odrv4 I__5128 (
            .O(N__25804),
            .I(\POWERLED.un1_N_3_mux_0 ));
    LocalMux I__5127 (
            .O(N__25801),
            .I(\POWERLED.un1_N_3_mux_0 ));
    CascadeMux I__5126 (
            .O(N__25792),
            .I(N_4_1_cascade_));
    InMux I__5125 (
            .O(N__25789),
            .I(N__25786));
    LocalMux I__5124 (
            .O(N__25786),
            .I(\POWERLED.count_clk_0_7 ));
    InMux I__5123 (
            .O(N__25783),
            .I(N__25780));
    LocalMux I__5122 (
            .O(N__25780),
            .I(\POWERLED.count_clk_0_9 ));
    InMux I__5121 (
            .O(N__25777),
            .I(N__25774));
    LocalMux I__5120 (
            .O(N__25774),
            .I(N__25771));
    Span4Mux_v I__5119 (
            .O(N__25771),
            .I(N__25768));
    Span4Mux_h I__5118 (
            .O(N__25768),
            .I(N__25765));
    Span4Mux_h I__5117 (
            .O(N__25765),
            .I(N__25762));
    Odrv4 I__5116 (
            .O(N__25762),
            .I(\POWERLED.count_off_0_5 ));
    InMux I__5115 (
            .O(N__25759),
            .I(N__25756));
    LocalMux I__5114 (
            .O(N__25756),
            .I(N__25752));
    InMux I__5113 (
            .O(N__25755),
            .I(N__25749));
    Span4Mux_v I__5112 (
            .O(N__25752),
            .I(N__25746));
    LocalMux I__5111 (
            .O(N__25749),
            .I(N__25743));
    Span4Mux_h I__5110 (
            .O(N__25746),
            .I(N__25740));
    Odrv12 I__5109 (
            .O(N__25743),
            .I(\POWERLED.count_off_1_5 ));
    Odrv4 I__5108 (
            .O(N__25740),
            .I(\POWERLED.count_off_1_5 ));
    InMux I__5107 (
            .O(N__25735),
            .I(N__25731));
    InMux I__5106 (
            .O(N__25734),
            .I(N__25728));
    LocalMux I__5105 (
            .O(N__25731),
            .I(N__25725));
    LocalMux I__5104 (
            .O(N__25728),
            .I(N__25722));
    Span4Mux_h I__5103 (
            .O(N__25725),
            .I(N__25719));
    Sp12to4 I__5102 (
            .O(N__25722),
            .I(N__25716));
    Span4Mux_v I__5101 (
            .O(N__25719),
            .I(N__25713));
    Odrv12 I__5100 (
            .O(N__25716),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__5099 (
            .O(N__25713),
            .I(\POWERLED.count_offZ0Z_5 ));
    InMux I__5098 (
            .O(N__25708),
            .I(N__25705));
    LocalMux I__5097 (
            .O(N__25705),
            .I(N__25702));
    Span4Mux_h I__5096 (
            .O(N__25702),
            .I(N__25699));
    Span4Mux_h I__5095 (
            .O(N__25699),
            .I(N__25696));
    Span4Mux_v I__5094 (
            .O(N__25696),
            .I(N__25693));
    Odrv4 I__5093 (
            .O(N__25693),
            .I(\POWERLED.count_off_0_6 ));
    InMux I__5092 (
            .O(N__25690),
            .I(N__25686));
    InMux I__5091 (
            .O(N__25689),
            .I(N__25683));
    LocalMux I__5090 (
            .O(N__25686),
            .I(N__25680));
    LocalMux I__5089 (
            .O(N__25683),
            .I(N__25677));
    Span12Mux_s6_h I__5088 (
            .O(N__25680),
            .I(N__25674));
    Odrv12 I__5087 (
            .O(N__25677),
            .I(\POWERLED.count_off_1_6 ));
    Odrv12 I__5086 (
            .O(N__25674),
            .I(\POWERLED.count_off_1_6 ));
    InMux I__5085 (
            .O(N__25669),
            .I(N__25665));
    InMux I__5084 (
            .O(N__25668),
            .I(N__25662));
    LocalMux I__5083 (
            .O(N__25665),
            .I(N__25659));
    LocalMux I__5082 (
            .O(N__25662),
            .I(N__25656));
    Span4Mux_h I__5081 (
            .O(N__25659),
            .I(N__25653));
    Span12Mux_s8_v I__5080 (
            .O(N__25656),
            .I(N__25650));
    Span4Mux_v I__5079 (
            .O(N__25653),
            .I(N__25647));
    Odrv12 I__5078 (
            .O(N__25650),
            .I(\POWERLED.count_offZ0Z_6 ));
    Odrv4 I__5077 (
            .O(N__25647),
            .I(\POWERLED.count_offZ0Z_6 ));
    InMux I__5076 (
            .O(N__25642),
            .I(N__25639));
    LocalMux I__5075 (
            .O(N__25639),
            .I(N__25636));
    Span4Mux_h I__5074 (
            .O(N__25636),
            .I(N__25633));
    Span4Mux_h I__5073 (
            .O(N__25633),
            .I(N__25630));
    Span4Mux_v I__5072 (
            .O(N__25630),
            .I(N__25627));
    Odrv4 I__5071 (
            .O(N__25627),
            .I(\POWERLED.count_off_0_2 ));
    InMux I__5070 (
            .O(N__25624),
            .I(N__25621));
    LocalMux I__5069 (
            .O(N__25621),
            .I(N__25617));
    InMux I__5068 (
            .O(N__25620),
            .I(N__25614));
    Span4Mux_v I__5067 (
            .O(N__25617),
            .I(N__25611));
    LocalMux I__5066 (
            .O(N__25614),
            .I(N__25608));
    Span4Mux_v I__5065 (
            .O(N__25611),
            .I(N__25605));
    Span4Mux_h I__5064 (
            .O(N__25608),
            .I(N__25602));
    Odrv4 I__5063 (
            .O(N__25605),
            .I(\POWERLED.count_off_1_2 ));
    Odrv4 I__5062 (
            .O(N__25602),
            .I(\POWERLED.count_off_1_2 ));
    CEMux I__5061 (
            .O(N__25597),
            .I(N__25593));
    CEMux I__5060 (
            .O(N__25596),
            .I(N__25587));
    LocalMux I__5059 (
            .O(N__25593),
            .I(N__25584));
    CEMux I__5058 (
            .O(N__25592),
            .I(N__25580));
    CascadeMux I__5057 (
            .O(N__25591),
            .I(N__25575));
    CEMux I__5056 (
            .O(N__25590),
            .I(N__25571));
    LocalMux I__5055 (
            .O(N__25587),
            .I(N__25565));
    Span4Mux_v I__5054 (
            .O(N__25584),
            .I(N__25562));
    CEMux I__5053 (
            .O(N__25583),
            .I(N__25559));
    LocalMux I__5052 (
            .O(N__25580),
            .I(N__25554));
    InMux I__5051 (
            .O(N__25579),
            .I(N__25541));
    InMux I__5050 (
            .O(N__25578),
            .I(N__25541));
    InMux I__5049 (
            .O(N__25575),
            .I(N__25541));
    InMux I__5048 (
            .O(N__25574),
            .I(N__25541));
    LocalMux I__5047 (
            .O(N__25571),
            .I(N__25538));
    InMux I__5046 (
            .O(N__25570),
            .I(N__25531));
    InMux I__5045 (
            .O(N__25569),
            .I(N__25531));
    InMux I__5044 (
            .O(N__25568),
            .I(N__25531));
    Span4Mux_v I__5043 (
            .O(N__25565),
            .I(N__25528));
    Span4Mux_h I__5042 (
            .O(N__25562),
            .I(N__25523));
    LocalMux I__5041 (
            .O(N__25559),
            .I(N__25523));
    InMux I__5040 (
            .O(N__25558),
            .I(N__25518));
    CEMux I__5039 (
            .O(N__25557),
            .I(N__25518));
    Span4Mux_h I__5038 (
            .O(N__25554),
            .I(N__25514));
    InMux I__5037 (
            .O(N__25553),
            .I(N__25505));
    InMux I__5036 (
            .O(N__25552),
            .I(N__25505));
    InMux I__5035 (
            .O(N__25551),
            .I(N__25505));
    InMux I__5034 (
            .O(N__25550),
            .I(N__25505));
    LocalMux I__5033 (
            .O(N__25541),
            .I(N__25502));
    Span4Mux_h I__5032 (
            .O(N__25538),
            .I(N__25497));
    LocalMux I__5031 (
            .O(N__25531),
            .I(N__25497));
    Span4Mux_h I__5030 (
            .O(N__25528),
            .I(N__25492));
    Span4Mux_h I__5029 (
            .O(N__25523),
            .I(N__25489));
    LocalMux I__5028 (
            .O(N__25518),
            .I(N__25486));
    InMux I__5027 (
            .O(N__25517),
            .I(N__25483));
    Span4Mux_s3_h I__5026 (
            .O(N__25514),
            .I(N__25474));
    LocalMux I__5025 (
            .O(N__25505),
            .I(N__25474));
    Span4Mux_v I__5024 (
            .O(N__25502),
            .I(N__25474));
    Span4Mux_v I__5023 (
            .O(N__25497),
            .I(N__25474));
    InMux I__5022 (
            .O(N__25496),
            .I(N__25469));
    InMux I__5021 (
            .O(N__25495),
            .I(N__25469));
    Odrv4 I__5020 (
            .O(N__25492),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0 ));
    Odrv4 I__5019 (
            .O(N__25489),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0 ));
    Odrv4 I__5018 (
            .O(N__25486),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0 ));
    LocalMux I__5017 (
            .O(N__25483),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0 ));
    Odrv4 I__5016 (
            .O(N__25474),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0 ));
    LocalMux I__5015 (
            .O(N__25469),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0 ));
    InMux I__5014 (
            .O(N__25456),
            .I(N__25452));
    InMux I__5013 (
            .O(N__25455),
            .I(N__25449));
    LocalMux I__5012 (
            .O(N__25452),
            .I(N__25446));
    LocalMux I__5011 (
            .O(N__25449),
            .I(N__25441));
    Span4Mux_h I__5010 (
            .O(N__25446),
            .I(N__25441));
    Span4Mux_v I__5009 (
            .O(N__25441),
            .I(N__25438));
    Odrv4 I__5008 (
            .O(N__25438),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__5007 (
            .O(N__25435),
            .I(N__25432));
    LocalMux I__5006 (
            .O(N__25432),
            .I(N__25428));
    CascadeMux I__5005 (
            .O(N__25431),
            .I(N__25423));
    Span4Mux_v I__5004 (
            .O(N__25428),
            .I(N__25419));
    InMux I__5003 (
            .O(N__25427),
            .I(N__25416));
    InMux I__5002 (
            .O(N__25426),
            .I(N__25413));
    InMux I__5001 (
            .O(N__25423),
            .I(N__25408));
    InMux I__5000 (
            .O(N__25422),
            .I(N__25408));
    Sp12to4 I__4999 (
            .O(N__25419),
            .I(N__25400));
    LocalMux I__4998 (
            .O(N__25416),
            .I(N__25400));
    LocalMux I__4997 (
            .O(N__25413),
            .I(N__25395));
    LocalMux I__4996 (
            .O(N__25408),
            .I(N__25395));
    InMux I__4995 (
            .O(N__25407),
            .I(N__25390));
    InMux I__4994 (
            .O(N__25406),
            .I(N__25390));
    InMux I__4993 (
            .O(N__25405),
            .I(N__25387));
    Odrv12 I__4992 (
            .O(N__25400),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__4991 (
            .O(N__25395),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4990 (
            .O(N__25390),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4989 (
            .O(N__25387),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    InMux I__4988 (
            .O(N__25378),
            .I(N__25372));
    CascadeMux I__4987 (
            .O(N__25377),
            .I(N__25367));
    InMux I__4986 (
            .O(N__25376),
            .I(N__25362));
    InMux I__4985 (
            .O(N__25375),
            .I(N__25359));
    LocalMux I__4984 (
            .O(N__25372),
            .I(N__25356));
    InMux I__4983 (
            .O(N__25371),
            .I(N__25353));
    CascadeMux I__4982 (
            .O(N__25370),
            .I(N__25350));
    InMux I__4981 (
            .O(N__25367),
            .I(N__25345));
    InMux I__4980 (
            .O(N__25366),
            .I(N__25345));
    InMux I__4979 (
            .O(N__25365),
            .I(N__25342));
    LocalMux I__4978 (
            .O(N__25362),
            .I(N__25338));
    LocalMux I__4977 (
            .O(N__25359),
            .I(N__25331));
    Span4Mux_h I__4976 (
            .O(N__25356),
            .I(N__25331));
    LocalMux I__4975 (
            .O(N__25353),
            .I(N__25331));
    InMux I__4974 (
            .O(N__25350),
            .I(N__25328));
    LocalMux I__4973 (
            .O(N__25345),
            .I(N__25323));
    LocalMux I__4972 (
            .O(N__25342),
            .I(N__25323));
    InMux I__4971 (
            .O(N__25341),
            .I(N__25320));
    Span4Mux_h I__4970 (
            .O(N__25338),
            .I(N__25313));
    Span4Mux_h I__4969 (
            .O(N__25331),
            .I(N__25313));
    LocalMux I__4968 (
            .O(N__25328),
            .I(N__25313));
    Odrv12 I__4967 (
            .O(N__25323),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4966 (
            .O(N__25320),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__4965 (
            .O(N__25313),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    InMux I__4964 (
            .O(N__25306),
            .I(N__25302));
    InMux I__4963 (
            .O(N__25305),
            .I(N__25299));
    LocalMux I__4962 (
            .O(N__25302),
            .I(N__25296));
    LocalMux I__4961 (
            .O(N__25299),
            .I(N__25293));
    Span4Mux_h I__4960 (
            .O(N__25296),
            .I(N__25290));
    Odrv4 I__4959 (
            .O(N__25293),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_13 ));
    Odrv4 I__4958 (
            .O(N__25290),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_13 ));
    InMux I__4957 (
            .O(N__25285),
            .I(N__25282));
    LocalMux I__4956 (
            .O(N__25282),
            .I(N__25279));
    Span4Mux_h I__4955 (
            .O(N__25279),
            .I(N__25276));
    Odrv4 I__4954 (
            .O(N__25276),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_15 ));
    CascadeMux I__4953 (
            .O(N__25273),
            .I(N__25263));
    InMux I__4952 (
            .O(N__25272),
            .I(N__25252));
    InMux I__4951 (
            .O(N__25271),
            .I(N__25252));
    InMux I__4950 (
            .O(N__25270),
            .I(N__25252));
    InMux I__4949 (
            .O(N__25269),
            .I(N__25252));
    InMux I__4948 (
            .O(N__25268),
            .I(N__25252));
    InMux I__4947 (
            .O(N__25267),
            .I(N__25247));
    InMux I__4946 (
            .O(N__25266),
            .I(N__25247));
    InMux I__4945 (
            .O(N__25263),
            .I(N__25244));
    LocalMux I__4944 (
            .O(N__25252),
            .I(N__25241));
    LocalMux I__4943 (
            .O(N__25247),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__4942 (
            .O(N__25244),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv12 I__4941 (
            .O(N__25241),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__4940 (
            .O(N__25234),
            .I(N__25229));
    InMux I__4939 (
            .O(N__25233),
            .I(N__25222));
    InMux I__4938 (
            .O(N__25232),
            .I(N__25222));
    InMux I__4937 (
            .O(N__25229),
            .I(N__25222));
    LocalMux I__4936 (
            .O(N__25222),
            .I(N__25217));
    CascadeMux I__4935 (
            .O(N__25221),
            .I(N__25214));
    CascadeMux I__4934 (
            .O(N__25220),
            .I(N__25211));
    Span4Mux_s3_v I__4933 (
            .O(N__25217),
            .I(N__25204));
    InMux I__4932 (
            .O(N__25214),
            .I(N__25191));
    InMux I__4931 (
            .O(N__25211),
            .I(N__25191));
    InMux I__4930 (
            .O(N__25210),
            .I(N__25191));
    InMux I__4929 (
            .O(N__25209),
            .I(N__25191));
    InMux I__4928 (
            .O(N__25208),
            .I(N__25191));
    InMux I__4927 (
            .O(N__25207),
            .I(N__25191));
    Odrv4 I__4926 (
            .O(N__25204),
            .I(RSMRST_PWRGD_curr_state_0));
    LocalMux I__4925 (
            .O(N__25191),
            .I(RSMRST_PWRGD_curr_state_0));
    InMux I__4924 (
            .O(N__25186),
            .I(N__25183));
    LocalMux I__4923 (
            .O(N__25183),
            .I(\POWERLED.N_301 ));
    SRMux I__4922 (
            .O(N__25180),
            .I(N__25177));
    LocalMux I__4921 (
            .O(N__25177),
            .I(N__25174));
    Span4Mux_v I__4920 (
            .O(N__25174),
            .I(N__25169));
    SRMux I__4919 (
            .O(N__25173),
            .I(N__25166));
    InMux I__4918 (
            .O(N__25172),
            .I(N__25162));
    Span4Mux_s2_v I__4917 (
            .O(N__25169),
            .I(N__25157));
    LocalMux I__4916 (
            .O(N__25166),
            .I(N__25157));
    SRMux I__4915 (
            .O(N__25165),
            .I(N__25154));
    LocalMux I__4914 (
            .O(N__25162),
            .I(N__25151));
    Sp12to4 I__4913 (
            .O(N__25157),
            .I(N__25148));
    LocalMux I__4912 (
            .O(N__25154),
            .I(N__25145));
    Span4Mux_v I__4911 (
            .O(N__25151),
            .I(N__25142));
    Odrv12 I__4910 (
            .O(N__25148),
            .I(G_11));
    Odrv12 I__4909 (
            .O(N__25145),
            .I(G_11));
    Odrv4 I__4908 (
            .O(N__25142),
            .I(G_11));
    CEMux I__4907 (
            .O(N__25135),
            .I(N__25132));
    LocalMux I__4906 (
            .O(N__25132),
            .I(N__25129));
    Span4Mux_h I__4905 (
            .O(N__25129),
            .I(N__25126));
    Odrv4 I__4904 (
            .O(N__25126),
            .I(\RSMRST_PWRGD.N_29_2 ));
    CascadeMux I__4903 (
            .O(N__25123),
            .I(N__25114));
    InMux I__4902 (
            .O(N__25122),
            .I(N__25111));
    InMux I__4901 (
            .O(N__25121),
            .I(N__25107));
    CascadeMux I__4900 (
            .O(N__25120),
            .I(N__25103));
    CascadeMux I__4899 (
            .O(N__25119),
            .I(N__25100));
    InMux I__4898 (
            .O(N__25118),
            .I(N__25093));
    InMux I__4897 (
            .O(N__25117),
            .I(N__25090));
    InMux I__4896 (
            .O(N__25114),
            .I(N__25087));
    LocalMux I__4895 (
            .O(N__25111),
            .I(N__25084));
    InMux I__4894 (
            .O(N__25110),
            .I(N__25081));
    LocalMux I__4893 (
            .O(N__25107),
            .I(N__25078));
    InMux I__4892 (
            .O(N__25106),
            .I(N__25075));
    InMux I__4891 (
            .O(N__25103),
            .I(N__25062));
    InMux I__4890 (
            .O(N__25100),
            .I(N__25062));
    InMux I__4889 (
            .O(N__25099),
            .I(N__25062));
    InMux I__4888 (
            .O(N__25098),
            .I(N__25062));
    InMux I__4887 (
            .O(N__25097),
            .I(N__25062));
    InMux I__4886 (
            .O(N__25096),
            .I(N__25062));
    LocalMux I__4885 (
            .O(N__25093),
            .I(N__25051));
    LocalMux I__4884 (
            .O(N__25090),
            .I(N__25051));
    LocalMux I__4883 (
            .O(N__25087),
            .I(N__25051));
    Span4Mux_s3_v I__4882 (
            .O(N__25084),
            .I(N__25051));
    LocalMux I__4881 (
            .O(N__25081),
            .I(N__25051));
    Span4Mux_v I__4880 (
            .O(N__25078),
            .I(N__25048));
    LocalMux I__4879 (
            .O(N__25075),
            .I(N__25043));
    LocalMux I__4878 (
            .O(N__25062),
            .I(N__25043));
    Span4Mux_v I__4877 (
            .O(N__25051),
            .I(N__25040));
    Span4Mux_v I__4876 (
            .O(N__25048),
            .I(N__25035));
    Span4Mux_s2_v I__4875 (
            .O(N__25043),
            .I(N__25035));
    Span4Mux_v I__4874 (
            .O(N__25040),
            .I(N__25032));
    Odrv4 I__4873 (
            .O(N__25035),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__4872 (
            .O(N__25032),
            .I(COUNTER_un4_counter_7_THRU_CO));
    CascadeMux I__4871 (
            .O(N__25027),
            .I(N__25023));
    CascadeMux I__4870 (
            .O(N__25026),
            .I(N__25020));
    InMux I__4869 (
            .O(N__25023),
            .I(N__25013));
    InMux I__4868 (
            .O(N__25020),
            .I(N__25013));
    InMux I__4867 (
            .O(N__25019),
            .I(N__25010));
    InMux I__4866 (
            .O(N__25018),
            .I(N__25007));
    LocalMux I__4865 (
            .O(N__25013),
            .I(N__25004));
    LocalMux I__4864 (
            .O(N__25010),
            .I(N__25001));
    LocalMux I__4863 (
            .O(N__25007),
            .I(N__24998));
    Span4Mux_h I__4862 (
            .O(N__25004),
            .I(N__24995));
    Span4Mux_h I__4861 (
            .O(N__25001),
            .I(N__24992));
    Span4Mux_v I__4860 (
            .O(N__24998),
            .I(N__24988));
    Span4Mux_v I__4859 (
            .O(N__24995),
            .I(N__24985));
    Span4Mux_s2_h I__4858 (
            .O(N__24992),
            .I(N__24982));
    InMux I__4857 (
            .O(N__24991),
            .I(N__24979));
    Odrv4 I__4856 (
            .O(N__24988),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    Odrv4 I__4855 (
            .O(N__24985),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    Odrv4 I__4854 (
            .O(N__24982),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    LocalMux I__4853 (
            .O(N__24979),
            .I(\POWERLED.dutycycle_N_3_mux_0 ));
    InMux I__4852 (
            .O(N__24970),
            .I(N__24967));
    LocalMux I__4851 (
            .O(N__24967),
            .I(\VPP_VDDQ.count_2_0_8 ));
    InMux I__4850 (
            .O(N__24964),
            .I(N__24961));
    LocalMux I__4849 (
            .O(N__24961),
            .I(\VPP_VDDQ.count_2_0_9 ));
    CascadeMux I__4848 (
            .O(N__24958),
            .I(\VPP_VDDQ.count_2_1_9_cascade_ ));
    InMux I__4847 (
            .O(N__24955),
            .I(N__24952));
    LocalMux I__4846 (
            .O(N__24952),
            .I(\VPP_VDDQ.count_2_0_10 ));
    IoInMux I__4845 (
            .O(N__24949),
            .I(N__24946));
    LocalMux I__4844 (
            .O(N__24946),
            .I(N__24943));
    IoSpan4Mux I__4843 (
            .O(N__24943),
            .I(N__24939));
    IoInMux I__4842 (
            .O(N__24942),
            .I(N__24936));
    IoSpan4Mux I__4841 (
            .O(N__24939),
            .I(N__24930));
    LocalMux I__4840 (
            .O(N__24936),
            .I(N__24930));
    InMux I__4839 (
            .O(N__24935),
            .I(N__24927));
    IoSpan4Mux I__4838 (
            .O(N__24930),
            .I(N__24924));
    LocalMux I__4837 (
            .O(N__24927),
            .I(N__24921));
    Span4Mux_s3_h I__4836 (
            .O(N__24924),
            .I(N__24918));
    Span4Mux_h I__4835 (
            .O(N__24921),
            .I(N__24915));
    Span4Mux_h I__4834 (
            .O(N__24918),
            .I(N__24912));
    Span4Mux_v I__4833 (
            .O(N__24915),
            .I(N__24909));
    Span4Mux_h I__4832 (
            .O(N__24912),
            .I(N__24904));
    Span4Mux_v I__4831 (
            .O(N__24909),
            .I(N__24904));
    Odrv4 I__4830 (
            .O(N__24904),
            .I(v33a_ok));
    InMux I__4829 (
            .O(N__24901),
            .I(N__24898));
    LocalMux I__4828 (
            .O(N__24898),
            .I(N__24895));
    Span4Mux_v I__4827 (
            .O(N__24895),
            .I(N__24892));
    Sp12to4 I__4826 (
            .O(N__24892),
            .I(N__24889));
    Odrv12 I__4825 (
            .O(N__24889),
            .I(v5a_ok));
    InMux I__4824 (
            .O(N__24886),
            .I(N__24883));
    LocalMux I__4823 (
            .O(N__24883),
            .I(N__24879));
    CascadeMux I__4822 (
            .O(N__24882),
            .I(N__24876));
    Span4Mux_v I__4821 (
            .O(N__24879),
            .I(N__24873));
    InMux I__4820 (
            .O(N__24876),
            .I(N__24870));
    Span4Mux_h I__4819 (
            .O(N__24873),
            .I(N__24867));
    LocalMux I__4818 (
            .O(N__24870),
            .I(N__24864));
    Odrv4 I__4817 (
            .O(N__24867),
            .I(slp_susn));
    Odrv12 I__4816 (
            .O(N__24864),
            .I(slp_susn));
    IoInMux I__4815 (
            .O(N__24859),
            .I(N__24856));
    LocalMux I__4814 (
            .O(N__24856),
            .I(N__24852));
    InMux I__4813 (
            .O(N__24855),
            .I(N__24849));
    Span4Mux_s2_h I__4812 (
            .O(N__24852),
            .I(N__24846));
    LocalMux I__4811 (
            .O(N__24849),
            .I(N__24843));
    Sp12to4 I__4810 (
            .O(N__24846),
            .I(N__24838));
    Sp12to4 I__4809 (
            .O(N__24843),
            .I(N__24838));
    Span12Mux_s11_v I__4808 (
            .O(N__24838),
            .I(N__24835));
    Odrv12 I__4807 (
            .O(N__24835),
            .I(v1p8a_ok));
    CascadeMux I__4806 (
            .O(N__24832),
            .I(rsmrst_pwrgd_signal_cascade_));
    CascadeMux I__4805 (
            .O(N__24829),
            .I(\RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ));
    InMux I__4804 (
            .O(N__24826),
            .I(N__24822));
    CascadeMux I__4803 (
            .O(N__24825),
            .I(N__24819));
    LocalMux I__4802 (
            .O(N__24822),
            .I(N__24815));
    InMux I__4801 (
            .O(N__24819),
            .I(N__24810));
    InMux I__4800 (
            .O(N__24818),
            .I(N__24810));
    Odrv12 I__4799 (
            .O(N__24815),
            .I(N_382));
    LocalMux I__4798 (
            .O(N__24810),
            .I(N_382));
    CascadeMux I__4797 (
            .O(N__24805),
            .I(N__24801));
    InMux I__4796 (
            .O(N__24804),
            .I(N__24798));
    InMux I__4795 (
            .O(N__24801),
            .I(N__24795));
    LocalMux I__4794 (
            .O(N__24798),
            .I(N__24792));
    LocalMux I__4793 (
            .O(N__24795),
            .I(N__24789));
    Span4Mux_v I__4792 (
            .O(N__24792),
            .I(N__24784));
    Span4Mux_v I__4791 (
            .O(N__24789),
            .I(N__24784));
    Odrv4 I__4790 (
            .O(N__24784),
            .I(\RSMRST_PWRGD.N_254_i ));
    InMux I__4789 (
            .O(N__24781),
            .I(N__24777));
    InMux I__4788 (
            .O(N__24780),
            .I(N__24774));
    LocalMux I__4787 (
            .O(N__24777),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    LocalMux I__4786 (
            .O(N__24774),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__4785 (
            .O(N__24769),
            .I(N__24765));
    InMux I__4784 (
            .O(N__24768),
            .I(N__24762));
    LocalMux I__4783 (
            .O(N__24765),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__4782 (
            .O(N__24762),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    CascadeMux I__4781 (
            .O(N__24757),
            .I(N__24754));
    InMux I__4780 (
            .O(N__24754),
            .I(N__24751));
    LocalMux I__4779 (
            .O(N__24751),
            .I(N__24748));
    Span4Mux_h I__4778 (
            .O(N__24748),
            .I(N__24745));
    Odrv4 I__4777 (
            .O(N__24745),
            .I(\RSMRST_PWRGD.m4_0_a2_0 ));
    InMux I__4776 (
            .O(N__24742),
            .I(N__24738));
    InMux I__4775 (
            .O(N__24741),
            .I(N__24735));
    LocalMux I__4774 (
            .O(N__24738),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__4773 (
            .O(N__24735),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__4772 (
            .O(N__24730),
            .I(N__24727));
    LocalMux I__4771 (
            .O(N__24727),
            .I(\RSMRST_PWRGD.m4_0_a2_12 ));
    CascadeMux I__4770 (
            .O(N__24724),
            .I(\VPP_VDDQ.count_2_1_10_cascade_ ));
    InMux I__4769 (
            .O(N__24721),
            .I(N__24715));
    InMux I__4768 (
            .O(N__24720),
            .I(N__24715));
    LocalMux I__4767 (
            .O(N__24715),
            .I(N__24712));
    Span4Mux_h I__4766 (
            .O(N__24712),
            .I(N__24707));
    InMux I__4765 (
            .O(N__24711),
            .I(N__24704));
    InMux I__4764 (
            .O(N__24710),
            .I(N__24701));
    Odrv4 I__4763 (
            .O(N__24707),
            .I(\PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0 ));
    LocalMux I__4762 (
            .O(N__24704),
            .I(\PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0 ));
    LocalMux I__4761 (
            .O(N__24701),
            .I(\PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0 ));
    InMux I__4760 (
            .O(N__24694),
            .I(N__24691));
    LocalMux I__4759 (
            .O(N__24691),
            .I(\PCH_PWRGD.curr_state_0_0 ));
    CascadeMux I__4758 (
            .O(N__24688),
            .I(\PCH_PWRGD.m4_0_cascade_ ));
    CascadeMux I__4757 (
            .O(N__24685),
            .I(\VPP_VDDQ.count_2_1_8_cascade_ ));
    CascadeMux I__4756 (
            .O(N__24682),
            .I(\PCH_PWRGD.countZ0Z_0_cascade_ ));
    InMux I__4755 (
            .O(N__24679),
            .I(N__24673));
    InMux I__4754 (
            .O(N__24678),
            .I(N__24673));
    LocalMux I__4753 (
            .O(N__24673),
            .I(\PCH_PWRGD.N_2173_i ));
    InMux I__4752 (
            .O(N__24670),
            .I(N__24666));
    InMux I__4751 (
            .O(N__24669),
            .I(N__24663));
    LocalMux I__4750 (
            .O(N__24666),
            .I(\PCH_PWRGD.count_1_i_a2_11_0 ));
    LocalMux I__4749 (
            .O(N__24663),
            .I(\PCH_PWRGD.count_1_i_a2_11_0 ));
    CascadeMux I__4748 (
            .O(N__24658),
            .I(\PCH_PWRGD.N_2173_i_cascade_ ));
    InMux I__4747 (
            .O(N__24655),
            .I(N__24651));
    InMux I__4746 (
            .O(N__24654),
            .I(N__24648));
    LocalMux I__4745 (
            .O(N__24651),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__4744 (
            .O(N__24648),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__4743 (
            .O(N__24643),
            .I(N__24639));
    InMux I__4742 (
            .O(N__24642),
            .I(N__24636));
    LocalMux I__4741 (
            .O(N__24639),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__4740 (
            .O(N__24636),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__4739 (
            .O(N__24631),
            .I(N__24627));
    InMux I__4738 (
            .O(N__24630),
            .I(N__24624));
    LocalMux I__4737 (
            .O(N__24627),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__4736 (
            .O(N__24624),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    CascadeMux I__4735 (
            .O(N__24619),
            .I(\RSMRST_PWRGD.m4_0_a2_11_cascade_ ));
    InMux I__4734 (
            .O(N__24616),
            .I(N__24612));
    InMux I__4733 (
            .O(N__24615),
            .I(N__24609));
    LocalMux I__4732 (
            .O(N__24612),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__4731 (
            .O(N__24609),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__4730 (
            .O(N__24604),
            .I(N__24600));
    InMux I__4729 (
            .O(N__24603),
            .I(N__24597));
    LocalMux I__4728 (
            .O(N__24600),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__4727 (
            .O(N__24597),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    CascadeMux I__4726 (
            .O(N__24592),
            .I(N__24588));
    InMux I__4725 (
            .O(N__24591),
            .I(N__24585));
    InMux I__4724 (
            .O(N__24588),
            .I(N__24582));
    LocalMux I__4723 (
            .O(N__24585),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__4722 (
            .O(N__24582),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__4721 (
            .O(N__24577),
            .I(N__24573));
    InMux I__4720 (
            .O(N__24576),
            .I(N__24570));
    LocalMux I__4719 (
            .O(N__24573),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__4718 (
            .O(N__24570),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__4717 (
            .O(N__24565),
            .I(N__24562));
    LocalMux I__4716 (
            .O(N__24562),
            .I(\RSMRST_PWRGD.m4_0_a2_10 ));
    InMux I__4715 (
            .O(N__24559),
            .I(N__24555));
    InMux I__4714 (
            .O(N__24558),
            .I(N__24552));
    LocalMux I__4713 (
            .O(N__24555),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__4712 (
            .O(N__24552),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    InMux I__4711 (
            .O(N__24547),
            .I(N__24543));
    InMux I__4710 (
            .O(N__24546),
            .I(N__24540));
    LocalMux I__4709 (
            .O(N__24543),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__4708 (
            .O(N__24540),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    CascadeMux I__4707 (
            .O(N__24535),
            .I(N__24531));
    InMux I__4706 (
            .O(N__24534),
            .I(N__24528));
    InMux I__4705 (
            .O(N__24531),
            .I(N__24525));
    LocalMux I__4704 (
            .O(N__24528),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__4703 (
            .O(N__24525),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__4702 (
            .O(N__24520),
            .I(N__24516));
    InMux I__4701 (
            .O(N__24519),
            .I(N__24513));
    LocalMux I__4700 (
            .O(N__24516),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__4699 (
            .O(N__24513),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__4698 (
            .O(N__24508),
            .I(N__24505));
    LocalMux I__4697 (
            .O(N__24505),
            .I(\RSMRST_PWRGD.m4_0_a2_9 ));
    InMux I__4696 (
            .O(N__24502),
            .I(N__24499));
    LocalMux I__4695 (
            .O(N__24499),
            .I(N__24496));
    Odrv4 I__4694 (
            .O(N__24496),
            .I(\PCH_PWRGD.count_0_6 ));
    InMux I__4693 (
            .O(N__24493),
            .I(N__24487));
    InMux I__4692 (
            .O(N__24492),
            .I(N__24487));
    LocalMux I__4691 (
            .O(N__24487),
            .I(\PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ));
    InMux I__4690 (
            .O(N__24484),
            .I(N__24481));
    LocalMux I__4689 (
            .O(N__24481),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__4688 (
            .O(N__24478),
            .I(N__24472));
    InMux I__4687 (
            .O(N__24477),
            .I(N__24472));
    LocalMux I__4686 (
            .O(N__24472),
            .I(\PCH_PWRGD.count_0_10 ));
    CascadeMux I__4685 (
            .O(N__24469),
            .I(\PCH_PWRGD.countZ0Z_6_cascade_ ));
    InMux I__4684 (
            .O(N__24466),
            .I(N__24461));
    InMux I__4683 (
            .O(N__24465),
            .I(N__24456));
    InMux I__4682 (
            .O(N__24464),
            .I(N__24456));
    LocalMux I__4681 (
            .O(N__24461),
            .I(\PCH_PWRGD.count_rst_4 ));
    LocalMux I__4680 (
            .O(N__24456),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__4679 (
            .O(N__24451),
            .I(N__24448));
    LocalMux I__4678 (
            .O(N__24448),
            .I(N__24445));
    Odrv4 I__4677 (
            .O(N__24445),
            .I(\PCH_PWRGD.count_1_i_a2_1_0 ));
    InMux I__4676 (
            .O(N__24442),
            .I(N__24439));
    LocalMux I__4675 (
            .O(N__24439),
            .I(N__24435));
    InMux I__4674 (
            .O(N__24438),
            .I(N__24432));
    Odrv4 I__4673 (
            .O(N__24435),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    LocalMux I__4672 (
            .O(N__24432),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    CascadeMux I__4671 (
            .O(N__24427),
            .I(\PCH_PWRGD.count_1_i_a2_0_0_cascade_ ));
    InMux I__4670 (
            .O(N__24424),
            .I(N__24421));
    LocalMux I__4669 (
            .O(N__24421),
            .I(N__24418));
    Span4Mux_v I__4668 (
            .O(N__24418),
            .I(N__24415));
    Odrv4 I__4667 (
            .O(N__24415),
            .I(\PCH_PWRGD.count_1_i_a2_2_0 ));
    CascadeMux I__4666 (
            .O(N__24412),
            .I(\PCH_PWRGD.count_1_i_a2_11_0_cascade_ ));
    CascadeMux I__4665 (
            .O(N__24409),
            .I(\PCH_PWRGD.count_rst_3_cascade_ ));
    CascadeMux I__4664 (
            .O(N__24406),
            .I(N_253_cascade_));
    InMux I__4663 (
            .O(N__24403),
            .I(N__24400));
    LocalMux I__4662 (
            .O(N__24400),
            .I(\PCH_PWRGD.count_0_0 ));
    InMux I__4661 (
            .O(N__24397),
            .I(N__24394));
    LocalMux I__4660 (
            .O(N__24394),
            .I(\PCH_PWRGD.count_RNIM6A821Z0Z_1 ));
    CascadeMux I__4659 (
            .O(N__24391),
            .I(\PCH_PWRGD.countZ0Z_3_cascade_ ));
    InMux I__4658 (
            .O(N__24388),
            .I(N__24382));
    InMux I__4657 (
            .O(N__24387),
            .I(N__24382));
    LocalMux I__4656 (
            .O(N__24382),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    InMux I__4655 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__4654 (
            .O(N__24376),
            .I(\PCH_PWRGD.count_0_3 ));
    CascadeMux I__4653 (
            .O(N__24373),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__4652 (
            .O(N__24370),
            .I(\PCH_PWRGD.countZ0Z_8_cascade_ ));
    InMux I__4651 (
            .O(N__24367),
            .I(N__24361));
    InMux I__4650 (
            .O(N__24366),
            .I(N__24361));
    LocalMux I__4649 (
            .O(N__24361),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__4648 (
            .O(N__24358),
            .I(N__24355));
    LocalMux I__4647 (
            .O(N__24355),
            .I(\PCH_PWRGD.count_0_8 ));
    InMux I__4646 (
            .O(N__24352),
            .I(N__24349));
    LocalMux I__4645 (
            .O(N__24349),
            .I(\PCH_PWRGD.un2_count_1_axb_10 ));
    InMux I__4644 (
            .O(N__24346),
            .I(N__24343));
    LocalMux I__4643 (
            .O(N__24343),
            .I(N__24339));
    InMux I__4642 (
            .O(N__24342),
            .I(N__24336));
    Odrv4 I__4641 (
            .O(N__24339),
            .I(\POWERLED.dutycycle_RNIZ0Z_6 ));
    LocalMux I__4640 (
            .O(N__24336),
            .I(\POWERLED.dutycycle_RNIZ0Z_6 ));
    InMux I__4639 (
            .O(N__24331),
            .I(N__24327));
    InMux I__4638 (
            .O(N__24330),
            .I(N__24324));
    LocalMux I__4637 (
            .O(N__24327),
            .I(N__24319));
    LocalMux I__4636 (
            .O(N__24324),
            .I(N__24319));
    Span12Mux_s10_v I__4635 (
            .O(N__24319),
            .I(N__24316));
    Odrv12 I__4634 (
            .O(N__24316),
            .I(\POWERLED.un1_dutycycle_172_m3s4_1 ));
    InMux I__4633 (
            .O(N__24313),
            .I(N__24307));
    InMux I__4632 (
            .O(N__24312),
            .I(N__24307));
    LocalMux I__4631 (
            .O(N__24307),
            .I(N__24302));
    InMux I__4630 (
            .O(N__24306),
            .I(N__24297));
    InMux I__4629 (
            .O(N__24305),
            .I(N__24297));
    Odrv12 I__4628 (
            .O(N__24302),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_6 ));
    LocalMux I__4627 (
            .O(N__24297),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_6 ));
    InMux I__4626 (
            .O(N__24292),
            .I(N__24289));
    LocalMux I__4625 (
            .O(N__24289),
            .I(\POWERLED.N_239 ));
    InMux I__4624 (
            .O(N__24286),
            .I(N__24283));
    LocalMux I__4623 (
            .O(N__24283),
            .I(N__24279));
    InMux I__4622 (
            .O(N__24282),
            .I(N__24276));
    Span4Mux_v I__4621 (
            .O(N__24279),
            .I(N__24273));
    LocalMux I__4620 (
            .O(N__24276),
            .I(N__24270));
    Odrv4 I__4619 (
            .O(N__24273),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    Odrv12 I__4618 (
            .O(N__24270),
            .I(\POWERLED.func_state_RNI_0Z0Z_0 ));
    CascadeMux I__4617 (
            .O(N__24265),
            .I(N__24262));
    InMux I__4616 (
            .O(N__24262),
            .I(N__24259));
    LocalMux I__4615 (
            .O(N__24259),
            .I(N__24256));
    Odrv4 I__4614 (
            .O(N__24256),
            .I(\POWERLED.N_271 ));
    InMux I__4613 (
            .O(N__24253),
            .I(N__24250));
    LocalMux I__4612 (
            .O(N__24250),
            .I(N__24247));
    Span4Mux_v I__4611 (
            .O(N__24247),
            .I(N__24243));
    InMux I__4610 (
            .O(N__24246),
            .I(N__24240));
    Odrv4 I__4609 (
            .O(N__24243),
            .I(\POWERLED.N_366 ));
    LocalMux I__4608 (
            .O(N__24240),
            .I(\POWERLED.N_366 ));
    CascadeMux I__4607 (
            .O(N__24235),
            .I(N__24230));
    InMux I__4606 (
            .O(N__24234),
            .I(N__24221));
    InMux I__4605 (
            .O(N__24233),
            .I(N__24221));
    InMux I__4604 (
            .O(N__24230),
            .I(N__24221));
    CascadeMux I__4603 (
            .O(N__24229),
            .I(N__24218));
    InMux I__4602 (
            .O(N__24228),
            .I(N__24214));
    LocalMux I__4601 (
            .O(N__24221),
            .I(N__24211));
    InMux I__4600 (
            .O(N__24218),
            .I(N__24208));
    InMux I__4599 (
            .O(N__24217),
            .I(N__24205));
    LocalMux I__4598 (
            .O(N__24214),
            .I(N__24202));
    Span4Mux_v I__4597 (
            .O(N__24211),
            .I(N__24197));
    LocalMux I__4596 (
            .O(N__24208),
            .I(N__24197));
    LocalMux I__4595 (
            .O(N__24205),
            .I(\POWERLED.N_331 ));
    Odrv4 I__4594 (
            .O(N__24202),
            .I(\POWERLED.N_331 ));
    Odrv4 I__4593 (
            .O(N__24197),
            .I(\POWERLED.N_331 ));
    InMux I__4592 (
            .O(N__24190),
            .I(N__24187));
    LocalMux I__4591 (
            .O(N__24187),
            .I(\POWERLED.N_272 ));
    CascadeMux I__4590 (
            .O(N__24184),
            .I(N__24181));
    InMux I__4589 (
            .O(N__24181),
            .I(N__24178));
    LocalMux I__4588 (
            .O(N__24178),
            .I(N__24175));
    Odrv12 I__4587 (
            .O(N__24175),
            .I(\POWERLED.dutycycle_N_3_mux_0_0 ));
    InMux I__4586 (
            .O(N__24172),
            .I(N__24169));
    LocalMux I__4585 (
            .O(N__24169),
            .I(N__24166));
    Odrv12 I__4584 (
            .O(N__24166),
            .I(\PCH_PWRGD.count_rst_10 ));
    InMux I__4583 (
            .O(N__24163),
            .I(N__24160));
    LocalMux I__4582 (
            .O(N__24160),
            .I(N__24156));
    InMux I__4581 (
            .O(N__24159),
            .I(N__24153));
    Odrv4 I__4580 (
            .O(N__24156),
            .I(\PCH_PWRGD.count_0_4 ));
    LocalMux I__4579 (
            .O(N__24153),
            .I(\PCH_PWRGD.count_0_4 ));
    CascadeMux I__4578 (
            .O(N__24148),
            .I(\PCH_PWRGD.count_rst_11_cascade_ ));
    CascadeMux I__4577 (
            .O(N__24145),
            .I(N__24142));
    InMux I__4576 (
            .O(N__24142),
            .I(N__24135));
    InMux I__4575 (
            .O(N__24141),
            .I(N__24135));
    InMux I__4574 (
            .O(N__24140),
            .I(N__24132));
    LocalMux I__4573 (
            .O(N__24135),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__4572 (
            .O(N__24132),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    CascadeMux I__4571 (
            .O(N__24127),
            .I(\POWERLED.count_off_1_sqmuxa_cascade_ ));
    InMux I__4570 (
            .O(N__24124),
            .I(N__24121));
    LocalMux I__4569 (
            .O(N__24121),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_6 ));
    InMux I__4568 (
            .O(N__24118),
            .I(N__24115));
    LocalMux I__4567 (
            .O(N__24115),
            .I(N__24111));
    InMux I__4566 (
            .O(N__24114),
            .I(N__24108));
    Span4Mux_h I__4565 (
            .O(N__24111),
            .I(N__24105));
    LocalMux I__4564 (
            .O(N__24108),
            .I(N__24102));
    Span4Mux_h I__4563 (
            .O(N__24105),
            .I(N__24099));
    Span4Mux_v I__4562 (
            .O(N__24102),
            .I(N__24096));
    Span4Mux_v I__4561 (
            .O(N__24099),
            .I(N__24093));
    Odrv4 I__4560 (
            .O(N__24096),
            .I(\POWERLED.N_325 ));
    Odrv4 I__4559 (
            .O(N__24093),
            .I(\POWERLED.N_325 ));
    CascadeMux I__4558 (
            .O(N__24088),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_6_cascade_ ));
    InMux I__4557 (
            .O(N__24085),
            .I(N__24079));
    InMux I__4556 (
            .O(N__24084),
            .I(N__24074));
    InMux I__4555 (
            .O(N__24083),
            .I(N__24074));
    CascadeMux I__4554 (
            .O(N__24082),
            .I(N__24071));
    LocalMux I__4553 (
            .O(N__24079),
            .I(N__24066));
    LocalMux I__4552 (
            .O(N__24074),
            .I(N__24066));
    InMux I__4551 (
            .O(N__24071),
            .I(N__24063));
    Span4Mux_v I__4550 (
            .O(N__24066),
            .I(N__24060));
    LocalMux I__4549 (
            .O(N__24063),
            .I(N__24057));
    Odrv4 I__4548 (
            .O(N__24060),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    Odrv4 I__4547 (
            .O(N__24057),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    InMux I__4546 (
            .O(N__24052),
            .I(N__24048));
    InMux I__4545 (
            .O(N__24051),
            .I(N__24045));
    LocalMux I__4544 (
            .O(N__24048),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_0 ));
    LocalMux I__4543 (
            .O(N__24045),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_0 ));
    CascadeMux I__4542 (
            .O(N__24040),
            .I(N__24037));
    InMux I__4541 (
            .O(N__24037),
            .I(N__24033));
    InMux I__4540 (
            .O(N__24036),
            .I(N__24030));
    LocalMux I__4539 (
            .O(N__24033),
            .I(N__24027));
    LocalMux I__4538 (
            .O(N__24030),
            .I(N__24024));
    Odrv4 I__4537 (
            .O(N__24027),
            .I(\POWERLED.dutycycle_RNINH5P1Z0Z_2 ));
    Odrv4 I__4536 (
            .O(N__24024),
            .I(\POWERLED.dutycycle_RNINH5P1Z0Z_2 ));
    CascadeMux I__4535 (
            .O(N__24019),
            .I(N__24015));
    InMux I__4534 (
            .O(N__24018),
            .I(N__24010));
    InMux I__4533 (
            .O(N__24015),
            .I(N__24010));
    LocalMux I__4532 (
            .O(N__24010),
            .I(N__24006));
    InMux I__4531 (
            .O(N__24009),
            .I(N__24003));
    Odrv4 I__4530 (
            .O(N__24006),
            .I(\POWERLED.dutycycle_RNI4G9K2Z0Z_5 ));
    LocalMux I__4529 (
            .O(N__24003),
            .I(\POWERLED.dutycycle_RNI4G9K2Z0Z_5 ));
    CascadeMux I__4528 (
            .O(N__23998),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_0_cascade_ ));
    CascadeMux I__4527 (
            .O(N__23995),
            .I(\POWERLED.dutycycle_RNO_2Z0Z_5_cascade_ ));
    InMux I__4526 (
            .O(N__23992),
            .I(N__23989));
    LocalMux I__4525 (
            .O(N__23989),
            .I(N__23986));
    Odrv4 I__4524 (
            .O(N__23986),
            .I(\POWERLED.N_240 ));
    CascadeMux I__4523 (
            .O(N__23983),
            .I(N__23979));
    InMux I__4522 (
            .O(N__23982),
            .I(N__23976));
    InMux I__4521 (
            .O(N__23979),
            .I(N__23973));
    LocalMux I__4520 (
            .O(N__23976),
            .I(N__23968));
    LocalMux I__4519 (
            .O(N__23973),
            .I(N__23968));
    Span4Mux_h I__4518 (
            .O(N__23968),
            .I(N__23965));
    Span4Mux_v I__4517 (
            .O(N__23965),
            .I(N__23962));
    Odrv4 I__4516 (
            .O(N__23962),
            .I(\POWERLED.dutycycle_eena_13 ));
    InMux I__4515 (
            .O(N__23959),
            .I(N__23956));
    LocalMux I__4514 (
            .O(N__23956),
            .I(N__23953));
    Span4Mux_h I__4513 (
            .O(N__23953),
            .I(N__23950));
    Odrv4 I__4512 (
            .O(N__23950),
            .I(\POWERLED.un2_count_clk_17_0_0 ));
    InMux I__4511 (
            .O(N__23947),
            .I(N__23944));
    LocalMux I__4510 (
            .O(N__23944),
            .I(\POWERLED.g3 ));
    CascadeMux I__4509 (
            .O(N__23941),
            .I(\POWERLED.un1_dutycycle_172_m3_1_0_cascade_ ));
    InMux I__4508 (
            .O(N__23938),
            .I(N__23935));
    LocalMux I__4507 (
            .O(N__23935),
            .I(\POWERLED.dutycycle_RNO_3Z0Z_5 ));
    InMux I__4506 (
            .O(N__23932),
            .I(N__23927));
    InMux I__4505 (
            .O(N__23931),
            .I(N__23922));
    InMux I__4504 (
            .O(N__23930),
            .I(N__23922));
    LocalMux I__4503 (
            .O(N__23927),
            .I(\POWERLED.dutycycle_1_0_5 ));
    LocalMux I__4502 (
            .O(N__23922),
            .I(\POWERLED.dutycycle_1_0_5 ));
    CascadeMux I__4501 (
            .O(N__23917),
            .I(N__23914));
    InMux I__4500 (
            .O(N__23914),
            .I(N__23911));
    LocalMux I__4499 (
            .O(N__23911),
            .I(\POWERLED.dutycycle_fb_15_1_1 ));
    InMux I__4498 (
            .O(N__23908),
            .I(N__23905));
    LocalMux I__4497 (
            .O(N__23905),
            .I(N__23902));
    Span4Mux_v I__4496 (
            .O(N__23902),
            .I(N__23899));
    Odrv4 I__4495 (
            .O(N__23899),
            .I(\POWERLED.g2_0 ));
    InMux I__4494 (
            .O(N__23896),
            .I(N__23893));
    LocalMux I__4493 (
            .O(N__23893),
            .I(N__23890));
    Odrv12 I__4492 (
            .O(N__23890),
            .I(\POWERLED.N_398_0 ));
    InMux I__4491 (
            .O(N__23887),
            .I(N__23884));
    LocalMux I__4490 (
            .O(N__23884),
            .I(\POWERLED.g0_1_0 ));
    InMux I__4489 (
            .O(N__23881),
            .I(N__23876));
    InMux I__4488 (
            .O(N__23880),
            .I(N__23870));
    InMux I__4487 (
            .O(N__23879),
            .I(N__23870));
    LocalMux I__4486 (
            .O(N__23876),
            .I(N__23867));
    InMux I__4485 (
            .O(N__23875),
            .I(N__23864));
    LocalMux I__4484 (
            .O(N__23870),
            .I(N__23859));
    Span4Mux_v I__4483 (
            .O(N__23867),
            .I(N__23859));
    LocalMux I__4482 (
            .O(N__23864),
            .I(N__23856));
    Span4Mux_v I__4481 (
            .O(N__23859),
            .I(N__23851));
    Span4Mux_v I__4480 (
            .O(N__23856),
            .I(N__23851));
    Odrv4 I__4479 (
            .O(N__23851),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_10 ));
    InMux I__4478 (
            .O(N__23848),
            .I(N__23845));
    LocalMux I__4477 (
            .O(N__23845),
            .I(N__23842));
    Span4Mux_v I__4476 (
            .O(N__23842),
            .I(N__23839));
    Odrv4 I__4475 (
            .O(N__23839),
            .I(\POWERLED.func_state_1_m2s2_i_a3_0 ));
    CascadeMux I__4474 (
            .O(N__23836),
            .I(N__23833));
    InMux I__4473 (
            .O(N__23833),
            .I(N__23830));
    LocalMux I__4472 (
            .O(N__23830),
            .I(N__23823));
    InMux I__4471 (
            .O(N__23829),
            .I(N__23820));
    InMux I__4470 (
            .O(N__23828),
            .I(N__23813));
    InMux I__4469 (
            .O(N__23827),
            .I(N__23813));
    InMux I__4468 (
            .O(N__23826),
            .I(N__23813));
    Odrv4 I__4467 (
            .O(N__23823),
            .I(\POWERLED.dutycycle_0_5 ));
    LocalMux I__4466 (
            .O(N__23820),
            .I(\POWERLED.dutycycle_0_5 ));
    LocalMux I__4465 (
            .O(N__23813),
            .I(\POWERLED.dutycycle_0_5 ));
    InMux I__4464 (
            .O(N__23806),
            .I(N__23803));
    LocalMux I__4463 (
            .O(N__23803),
            .I(N__23800));
    Odrv4 I__4462 (
            .O(N__23800),
            .I(\POWERLED.dutycycle_fb_14_a4_1 ));
    CascadeMux I__4461 (
            .O(N__23797),
            .I(N__23793));
    CascadeMux I__4460 (
            .O(N__23796),
            .I(N__23787));
    InMux I__4459 (
            .O(N__23793),
            .I(N__23783));
    InMux I__4458 (
            .O(N__23792),
            .I(N__23778));
    InMux I__4457 (
            .O(N__23791),
            .I(N__23778));
    CascadeMux I__4456 (
            .O(N__23790),
            .I(N__23775));
    InMux I__4455 (
            .O(N__23787),
            .I(N__23770));
    InMux I__4454 (
            .O(N__23786),
            .I(N__23770));
    LocalMux I__4453 (
            .O(N__23783),
            .I(N__23765));
    LocalMux I__4452 (
            .O(N__23778),
            .I(N__23765));
    InMux I__4451 (
            .O(N__23775),
            .I(N__23762));
    LocalMux I__4450 (
            .O(N__23770),
            .I(N__23752));
    Span4Mux_v I__4449 (
            .O(N__23765),
            .I(N__23752));
    LocalMux I__4448 (
            .O(N__23762),
            .I(N__23749));
    InMux I__4447 (
            .O(N__23761),
            .I(N__23746));
    InMux I__4446 (
            .O(N__23760),
            .I(N__23741));
    InMux I__4445 (
            .O(N__23759),
            .I(N__23741));
    InMux I__4444 (
            .O(N__23758),
            .I(N__23738));
    InMux I__4443 (
            .O(N__23757),
            .I(N__23735));
    Span4Mux_h I__4442 (
            .O(N__23752),
            .I(N__23730));
    Span4Mux_v I__4441 (
            .O(N__23749),
            .I(N__23730));
    LocalMux I__4440 (
            .O(N__23746),
            .I(\POWERLED.dutycycle ));
    LocalMux I__4439 (
            .O(N__23741),
            .I(\POWERLED.dutycycle ));
    LocalMux I__4438 (
            .O(N__23738),
            .I(\POWERLED.dutycycle ));
    LocalMux I__4437 (
            .O(N__23735),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__4436 (
            .O(N__23730),
            .I(\POWERLED.dutycycle ));
    InMux I__4435 (
            .O(N__23719),
            .I(N__23716));
    LocalMux I__4434 (
            .O(N__23716),
            .I(\POWERLED.count_off_1_sqmuxa ));
    CascadeMux I__4433 (
            .O(N__23713),
            .I(\POWERLED.g0_9_1_cascade_ ));
    CascadeMux I__4432 (
            .O(N__23710),
            .I(\POWERLED.dutycycle_fb_15_4_0_cascade_ ));
    InMux I__4431 (
            .O(N__23707),
            .I(N__23704));
    LocalMux I__4430 (
            .O(N__23704),
            .I(\POWERLED.dutycycle_fb_15_0 ));
    CascadeMux I__4429 (
            .O(N__23701),
            .I(\POWERLED.dutycycle_en_14_cascade_ ));
    SRMux I__4428 (
            .O(N__23698),
            .I(N__23692));
    SRMux I__4427 (
            .O(N__23697),
            .I(N__23689));
    SRMux I__4426 (
            .O(N__23696),
            .I(N__23686));
    SRMux I__4425 (
            .O(N__23695),
            .I(N__23682));
    LocalMux I__4424 (
            .O(N__23692),
            .I(N__23677));
    LocalMux I__4423 (
            .O(N__23689),
            .I(N__23677));
    LocalMux I__4422 (
            .O(N__23686),
            .I(N__23674));
    SRMux I__4421 (
            .O(N__23685),
            .I(N__23671));
    LocalMux I__4420 (
            .O(N__23682),
            .I(N__23665));
    Span4Mux_v I__4419 (
            .O(N__23677),
            .I(N__23661));
    Span4Mux_v I__4418 (
            .O(N__23674),
            .I(N__23656));
    LocalMux I__4417 (
            .O(N__23671),
            .I(N__23656));
    SRMux I__4416 (
            .O(N__23670),
            .I(N__23653));
    SRMux I__4415 (
            .O(N__23669),
            .I(N__23650));
    SRMux I__4414 (
            .O(N__23668),
            .I(N__23647));
    Span4Mux_v I__4413 (
            .O(N__23665),
            .I(N__23643));
    SRMux I__4412 (
            .O(N__23664),
            .I(N__23640));
    Span4Mux_v I__4411 (
            .O(N__23661),
            .I(N__23637));
    Span4Mux_v I__4410 (
            .O(N__23656),
            .I(N__23634));
    LocalMux I__4409 (
            .O(N__23653),
            .I(N__23631));
    LocalMux I__4408 (
            .O(N__23650),
            .I(N__23628));
    LocalMux I__4407 (
            .O(N__23647),
            .I(N__23625));
    SRMux I__4406 (
            .O(N__23646),
            .I(N__23622));
    Span4Mux_v I__4405 (
            .O(N__23643),
            .I(N__23617));
    LocalMux I__4404 (
            .O(N__23640),
            .I(N__23617));
    Sp12to4 I__4403 (
            .O(N__23637),
            .I(N__23612));
    Span4Mux_h I__4402 (
            .O(N__23634),
            .I(N__23607));
    Span4Mux_v I__4401 (
            .O(N__23631),
            .I(N__23607));
    Span4Mux_v I__4400 (
            .O(N__23628),
            .I(N__23600));
    Span4Mux_h I__4399 (
            .O(N__23625),
            .I(N__23600));
    LocalMux I__4398 (
            .O(N__23622),
            .I(N__23600));
    Span4Mux_v I__4397 (
            .O(N__23617),
            .I(N__23597));
    SRMux I__4396 (
            .O(N__23616),
            .I(N__23594));
    SRMux I__4395 (
            .O(N__23615),
            .I(N__23591));
    Odrv12 I__4394 (
            .O(N__23612),
            .I(\POWERLED.func_m2_0_a2_isoZ0 ));
    Odrv4 I__4393 (
            .O(N__23607),
            .I(\POWERLED.func_m2_0_a2_isoZ0 ));
    Odrv4 I__4392 (
            .O(N__23600),
            .I(\POWERLED.func_m2_0_a2_isoZ0 ));
    Odrv4 I__4391 (
            .O(N__23597),
            .I(\POWERLED.func_m2_0_a2_isoZ0 ));
    LocalMux I__4390 (
            .O(N__23594),
            .I(\POWERLED.func_m2_0_a2_isoZ0 ));
    LocalMux I__4389 (
            .O(N__23591),
            .I(\POWERLED.func_m2_0_a2_isoZ0 ));
    InMux I__4388 (
            .O(N__23578),
            .I(N__23569));
    InMux I__4387 (
            .O(N__23577),
            .I(N__23569));
    InMux I__4386 (
            .O(N__23576),
            .I(N__23569));
    LocalMux I__4385 (
            .O(N__23569),
            .I(\POWERLED.dutycycle_eena_14_0Z0Z_0 ));
    InMux I__4384 (
            .O(N__23566),
            .I(N__23563));
    LocalMux I__4383 (
            .O(N__23563),
            .I(N__23560));
    Odrv4 I__4382 (
            .O(N__23560),
            .I(\POWERLED.dutycycle_fb_15_1 ));
    InMux I__4381 (
            .O(N__23557),
            .I(N__23554));
    LocalMux I__4380 (
            .O(N__23554),
            .I(\POWERLED.g1_0 ));
    InMux I__4379 (
            .O(N__23551),
            .I(N__23548));
    LocalMux I__4378 (
            .O(N__23548),
            .I(N__23545));
    Odrv12 I__4377 (
            .O(N__23545),
            .I(\POWERLED.g1 ));
    InMux I__4376 (
            .O(N__23542),
            .I(N__23539));
    LocalMux I__4375 (
            .O(N__23539),
            .I(\POWERLED.dutycycle_fb_15_2_0 ));
    CascadeMux I__4374 (
            .O(N__23536),
            .I(N__23529));
    InMux I__4373 (
            .O(N__23535),
            .I(N__23524));
    InMux I__4372 (
            .O(N__23534),
            .I(N__23524));
    InMux I__4371 (
            .O(N__23533),
            .I(N__23521));
    InMux I__4370 (
            .O(N__23532),
            .I(N__23518));
    InMux I__4369 (
            .O(N__23529),
            .I(N__23515));
    LocalMux I__4368 (
            .O(N__23524),
            .I(SUSWARN_N_rep1));
    LocalMux I__4367 (
            .O(N__23521),
            .I(SUSWARN_N_rep1));
    LocalMux I__4366 (
            .O(N__23518),
            .I(SUSWARN_N_rep1));
    LocalMux I__4365 (
            .O(N__23515),
            .I(SUSWARN_N_rep1));
    CascadeMux I__4364 (
            .O(N__23506),
            .I(\POWERLED.N_340_cascade_ ));
    InMux I__4363 (
            .O(N__23503),
            .I(N__23500));
    LocalMux I__4362 (
            .O(N__23500),
            .I(N__23497));
    Odrv4 I__4361 (
            .O(N__23497),
            .I(\POWERLED.func_state_RNIRAVV2Z0Z_0 ));
    InMux I__4360 (
            .O(N__23494),
            .I(N__23491));
    LocalMux I__4359 (
            .O(N__23491),
            .I(N__23488));
    Span4Mux_v I__4358 (
            .O(N__23488),
            .I(N__23485));
    Sp12to4 I__4357 (
            .O(N__23485),
            .I(N__23482));
    Odrv12 I__4356 (
            .O(N__23482),
            .I(\POWERLED.m18_e_5 ));
    InMux I__4355 (
            .O(N__23479),
            .I(N__23476));
    LocalMux I__4354 (
            .O(N__23476),
            .I(\POWERLED.m18_e_6 ));
    InMux I__4353 (
            .O(N__23473),
            .I(N__23470));
    LocalMux I__4352 (
            .O(N__23470),
            .I(\POWERLED.func_m2_0_a2Z0Z_0 ));
    CascadeMux I__4351 (
            .O(N__23467),
            .I(\POWERLED.func_m2_0_a2Z0Z_0_cascade_ ));
    InMux I__4350 (
            .O(N__23464),
            .I(N__23452));
    InMux I__4349 (
            .O(N__23463),
            .I(N__23452));
    InMux I__4348 (
            .O(N__23462),
            .I(N__23449));
    InMux I__4347 (
            .O(N__23461),
            .I(N__23444));
    InMux I__4346 (
            .O(N__23460),
            .I(N__23444));
    InMux I__4345 (
            .O(N__23459),
            .I(N__23441));
    InMux I__4344 (
            .O(N__23458),
            .I(N__23438));
    CascadeMux I__4343 (
            .O(N__23457),
            .I(N__23435));
    LocalMux I__4342 (
            .O(N__23452),
            .I(N__23432));
    LocalMux I__4341 (
            .O(N__23449),
            .I(N__23427));
    LocalMux I__4340 (
            .O(N__23444),
            .I(N__23427));
    LocalMux I__4339 (
            .O(N__23441),
            .I(N__23422));
    LocalMux I__4338 (
            .O(N__23438),
            .I(N__23422));
    InMux I__4337 (
            .O(N__23435),
            .I(N__23419));
    Span4Mux_h I__4336 (
            .O(N__23432),
            .I(N__23416));
    Span4Mux_v I__4335 (
            .O(N__23427),
            .I(N__23413));
    Span4Mux_h I__4334 (
            .O(N__23422),
            .I(N__23408));
    LocalMux I__4333 (
            .O(N__23419),
            .I(N__23408));
    Odrv4 I__4332 (
            .O(N__23416),
            .I(\POWERLED.count_clk_RNI2O4A1_0Z0Z_10 ));
    Odrv4 I__4331 (
            .O(N__23413),
            .I(\POWERLED.count_clk_RNI2O4A1_0Z0Z_10 ));
    Odrv4 I__4330 (
            .O(N__23408),
            .I(\POWERLED.count_clk_RNI2O4A1_0Z0Z_10 ));
    CascadeMux I__4329 (
            .O(N__23401),
            .I(\POWERLED.func_state_RNI91IA4_0Z0Z_1_cascade_ ));
    InMux I__4328 (
            .O(N__23398),
            .I(N__23395));
    LocalMux I__4327 (
            .O(N__23395),
            .I(\POWERLED.func_state_1_m2_0 ));
    InMux I__4326 (
            .O(N__23392),
            .I(N__23386));
    InMux I__4325 (
            .O(N__23391),
            .I(N__23386));
    LocalMux I__4324 (
            .O(N__23386),
            .I(\POWERLED.func_stateZ1Z_0 ));
    CascadeMux I__4323 (
            .O(N__23383),
            .I(\POWERLED.func_state_1_m2_0_cascade_ ));
    CascadeMux I__4322 (
            .O(N__23380),
            .I(N__23377));
    InMux I__4321 (
            .O(N__23377),
            .I(N__23366));
    InMux I__4320 (
            .O(N__23376),
            .I(N__23366));
    InMux I__4319 (
            .O(N__23375),
            .I(N__23361));
    InMux I__4318 (
            .O(N__23374),
            .I(N__23361));
    InMux I__4317 (
            .O(N__23373),
            .I(N__23358));
    InMux I__4316 (
            .O(N__23372),
            .I(N__23353));
    InMux I__4315 (
            .O(N__23371),
            .I(N__23353));
    LocalMux I__4314 (
            .O(N__23366),
            .I(N__23350));
    LocalMux I__4313 (
            .O(N__23361),
            .I(N__23347));
    LocalMux I__4312 (
            .O(N__23358),
            .I(N__23342));
    LocalMux I__4311 (
            .O(N__23353),
            .I(N__23339));
    Span4Mux_h I__4310 (
            .O(N__23350),
            .I(N__23336));
    Span4Mux_h I__4309 (
            .O(N__23347),
            .I(N__23333));
    InMux I__4308 (
            .O(N__23346),
            .I(N__23330));
    InMux I__4307 (
            .O(N__23345),
            .I(N__23327));
    Odrv4 I__4306 (
            .O(N__23342),
            .I(\POWERLED.N_335 ));
    Odrv12 I__4305 (
            .O(N__23339),
            .I(\POWERLED.N_335 ));
    Odrv4 I__4304 (
            .O(N__23336),
            .I(\POWERLED.N_335 ));
    Odrv4 I__4303 (
            .O(N__23333),
            .I(\POWERLED.N_335 ));
    LocalMux I__4302 (
            .O(N__23330),
            .I(\POWERLED.N_335 ));
    LocalMux I__4301 (
            .O(N__23327),
            .I(\POWERLED.N_335 ));
    CascadeMux I__4300 (
            .O(N__23314),
            .I(\POWERLED.func_state_RNI2O4A1Z0Z_1_cascade_ ));
    InMux I__4299 (
            .O(N__23311),
            .I(N__23305));
    InMux I__4298 (
            .O(N__23310),
            .I(N__23305));
    LocalMux I__4297 (
            .O(N__23305),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__4296 (
            .O(N__23302),
            .I(N__23299));
    InMux I__4295 (
            .O(N__23299),
            .I(N__23293));
    InMux I__4294 (
            .O(N__23298),
            .I(N__23293));
    LocalMux I__4293 (
            .O(N__23293),
            .I(\POWERLED.dutycycle_en_9 ));
    CascadeMux I__4292 (
            .O(N__23290),
            .I(\POWERLED.func_state_RNI2O4A1_1Z0Z_1_cascade_ ));
    InMux I__4291 (
            .O(N__23287),
            .I(N__23281));
    InMux I__4290 (
            .O(N__23286),
            .I(N__23281));
    LocalMux I__4289 (
            .O(N__23281),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ));
    InMux I__4288 (
            .O(N__23278),
            .I(N__23275));
    LocalMux I__4287 (
            .O(N__23275),
            .I(N__23270));
    CascadeMux I__4286 (
            .O(N__23274),
            .I(N__23262));
    CascadeMux I__4285 (
            .O(N__23273),
            .I(N__23257));
    Span4Mux_v I__4284 (
            .O(N__23270),
            .I(N__23254));
    InMux I__4283 (
            .O(N__23269),
            .I(N__23251));
    CascadeMux I__4282 (
            .O(N__23268),
            .I(N__23248));
    InMux I__4281 (
            .O(N__23267),
            .I(N__23244));
    InMux I__4280 (
            .O(N__23266),
            .I(N__23241));
    InMux I__4279 (
            .O(N__23265),
            .I(N__23230));
    InMux I__4278 (
            .O(N__23262),
            .I(N__23230));
    InMux I__4277 (
            .O(N__23261),
            .I(N__23230));
    InMux I__4276 (
            .O(N__23260),
            .I(N__23230));
    InMux I__4275 (
            .O(N__23257),
            .I(N__23230));
    Span4Mux_h I__4274 (
            .O(N__23254),
            .I(N__23224));
    LocalMux I__4273 (
            .O(N__23251),
            .I(N__23224));
    InMux I__4272 (
            .O(N__23248),
            .I(N__23219));
    InMux I__4271 (
            .O(N__23247),
            .I(N__23219));
    LocalMux I__4270 (
            .O(N__23244),
            .I(N__23214));
    LocalMux I__4269 (
            .O(N__23241),
            .I(N__23214));
    LocalMux I__4268 (
            .O(N__23230),
            .I(N__23211));
    CascadeMux I__4267 (
            .O(N__23229),
            .I(N__23208));
    Span4Mux_v I__4266 (
            .O(N__23224),
            .I(N__23205));
    LocalMux I__4265 (
            .O(N__23219),
            .I(N__23202));
    Span4Mux_h I__4264 (
            .O(N__23214),
            .I(N__23199));
    Span4Mux_h I__4263 (
            .O(N__23211),
            .I(N__23196));
    InMux I__4262 (
            .O(N__23208),
            .I(N__23193));
    Odrv4 I__4261 (
            .O(N__23205),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv12 I__4260 (
            .O(N__23202),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__4259 (
            .O(N__23199),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__4258 (
            .O(N__23196),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__4257 (
            .O(N__23193),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    CascadeMux I__4256 (
            .O(N__23182),
            .I(\POWERLED.dutycycleZ0Z_11_cascade_ ));
    InMux I__4255 (
            .O(N__23179),
            .I(N__23176));
    LocalMux I__4254 (
            .O(N__23176),
            .I(\POWERLED.un1_clk_100khz_42_and_i_0_0 ));
    InMux I__4253 (
            .O(N__23173),
            .I(N__23167));
    InMux I__4252 (
            .O(N__23172),
            .I(N__23167));
    LocalMux I__4251 (
            .O(N__23167),
            .I(N__23163));
    InMux I__4250 (
            .O(N__23166),
            .I(N__23159));
    Span12Mux_s7_h I__4249 (
            .O(N__23163),
            .I(N__23156));
    InMux I__4248 (
            .O(N__23162),
            .I(N__23153));
    LocalMux I__4247 (
            .O(N__23159),
            .I(\POWERLED.func_state_RNI2O4A1Z0Z_1 ));
    Odrv12 I__4246 (
            .O(N__23156),
            .I(\POWERLED.func_state_RNI2O4A1Z0Z_1 ));
    LocalMux I__4245 (
            .O(N__23153),
            .I(\POWERLED.func_state_RNI2O4A1Z0Z_1 ));
    CascadeMux I__4244 (
            .O(N__23146),
            .I(\POWERLED.un1_clk_100khz_47_and_i_0_0_cascade_ ));
    InMux I__4243 (
            .O(N__23143),
            .I(N__23137));
    InMux I__4242 (
            .O(N__23142),
            .I(N__23137));
    LocalMux I__4241 (
            .O(N__23137),
            .I(N__23133));
    CascadeMux I__4240 (
            .O(N__23136),
            .I(N__23130));
    Span4Mux_h I__4239 (
            .O(N__23133),
            .I(N__23126));
    InMux I__4238 (
            .O(N__23130),
            .I(N__23121));
    InMux I__4237 (
            .O(N__23129),
            .I(N__23121));
    Odrv4 I__4236 (
            .O(N__23126),
            .I(\POWERLED.N_399_N ));
    LocalMux I__4235 (
            .O(N__23121),
            .I(\POWERLED.N_399_N ));
    CascadeMux I__4234 (
            .O(N__23116),
            .I(N__23112));
    InMux I__4233 (
            .O(N__23115),
            .I(N__23109));
    InMux I__4232 (
            .O(N__23112),
            .I(N__23106));
    LocalMux I__4231 (
            .O(N__23109),
            .I(N__23101));
    LocalMux I__4230 (
            .O(N__23106),
            .I(N__23101));
    Span4Mux_h I__4229 (
            .O(N__23101),
            .I(N__23098));
    Odrv4 I__4228 (
            .O(N__23098),
            .I(\POWERLED.dutycycle_en_11 ));
    CascadeMux I__4227 (
            .O(N__23095),
            .I(\POWERLED.N_2216_i_cascade_ ));
    CascadeMux I__4226 (
            .O(N__23092),
            .I(\POWERLED.func_state_1_m2s2_i_1_cascade_ ));
    CascadeMux I__4225 (
            .O(N__23089),
            .I(N__23085));
    InMux I__4224 (
            .O(N__23088),
            .I(N__23080));
    InMux I__4223 (
            .O(N__23085),
            .I(N__23080));
    LocalMux I__4222 (
            .O(N__23080),
            .I(N__23077));
    Odrv4 I__4221 (
            .O(N__23077),
            .I(\POWERLED.N_160 ));
    CascadeMux I__4220 (
            .O(N__23074),
            .I(N__23065));
    InMux I__4219 (
            .O(N__23073),
            .I(N__23060));
    InMux I__4218 (
            .O(N__23072),
            .I(N__23060));
    InMux I__4217 (
            .O(N__23071),
            .I(N__23057));
    InMux I__4216 (
            .O(N__23070),
            .I(N__23052));
    InMux I__4215 (
            .O(N__23069),
            .I(N__23052));
    InMux I__4214 (
            .O(N__23068),
            .I(N__23047));
    InMux I__4213 (
            .O(N__23065),
            .I(N__23047));
    LocalMux I__4212 (
            .O(N__23060),
            .I(N__23044));
    LocalMux I__4211 (
            .O(N__23057),
            .I(N__23037));
    LocalMux I__4210 (
            .O(N__23052),
            .I(N__23037));
    LocalMux I__4209 (
            .O(N__23047),
            .I(N__23037));
    Span4Mux_h I__4208 (
            .O(N__23044),
            .I(N__23032));
    Span4Mux_v I__4207 (
            .O(N__23037),
            .I(N__23032));
    Odrv4 I__4206 (
            .O(N__23032),
            .I(\POWERLED.N_3_0 ));
    CascadeMux I__4205 (
            .O(N__23029),
            .I(slp_s3n_signal_cascade_));
    InMux I__4204 (
            .O(N__23026),
            .I(N__23020));
    InMux I__4203 (
            .O(N__23025),
            .I(N__23020));
    LocalMux I__4202 (
            .O(N__23020),
            .I(\POWERLED.N_183 ));
    CascadeMux I__4201 (
            .O(N__23017),
            .I(\POWERLED.func_state_RNIZ0Z_1_cascade_ ));
    InMux I__4200 (
            .O(N__23014),
            .I(N__22994));
    InMux I__4199 (
            .O(N__23013),
            .I(N__22994));
    InMux I__4198 (
            .O(N__23012),
            .I(N__22994));
    InMux I__4197 (
            .O(N__23011),
            .I(N__22987));
    InMux I__4196 (
            .O(N__23010),
            .I(N__22987));
    InMux I__4195 (
            .O(N__23009),
            .I(N__22987));
    InMux I__4194 (
            .O(N__23008),
            .I(N__22978));
    InMux I__4193 (
            .O(N__23007),
            .I(N__22978));
    InMux I__4192 (
            .O(N__23006),
            .I(N__22978));
    InMux I__4191 (
            .O(N__23005),
            .I(N__22978));
    InMux I__4190 (
            .O(N__23004),
            .I(N__22969));
    InMux I__4189 (
            .O(N__23003),
            .I(N__22969));
    InMux I__4188 (
            .O(N__23002),
            .I(N__22969));
    InMux I__4187 (
            .O(N__23001),
            .I(N__22969));
    LocalMux I__4186 (
            .O(N__22994),
            .I(\POWERLED.N_162_i ));
    LocalMux I__4185 (
            .O(N__22987),
            .I(\POWERLED.N_162_i ));
    LocalMux I__4184 (
            .O(N__22978),
            .I(\POWERLED.N_162_i ));
    LocalMux I__4183 (
            .O(N__22969),
            .I(\POWERLED.N_162_i ));
    InMux I__4182 (
            .O(N__22960),
            .I(N__22957));
    LocalMux I__4181 (
            .O(N__22957),
            .I(\POWERLED.count_off_0_1 ));
    CascadeMux I__4180 (
            .O(N__22954),
            .I(N__22951));
    InMux I__4179 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__4178 (
            .O(N__22948),
            .I(\POWERLED.count_off_RNIZ0Z_1 ));
    InMux I__4177 (
            .O(N__22945),
            .I(N__22942));
    LocalMux I__4176 (
            .O(N__22942),
            .I(N__22938));
    InMux I__4175 (
            .O(N__22941),
            .I(N__22935));
    Span4Mux_h I__4174 (
            .O(N__22938),
            .I(N__22932));
    LocalMux I__4173 (
            .O(N__22935),
            .I(\POWERLED.count_offZ0Z_1 ));
    Odrv4 I__4172 (
            .O(N__22932),
            .I(\POWERLED.count_offZ0Z_1 ));
    CascadeMux I__4171 (
            .O(N__22927),
            .I(\POWERLED.count_offZ0Z_1_cascade_ ));
    InMux I__4170 (
            .O(N__22924),
            .I(N__22921));
    LocalMux I__4169 (
            .O(N__22921),
            .I(\POWERLED.un34_clk_100khz_10 ));
    InMux I__4168 (
            .O(N__22918),
            .I(N__22915));
    LocalMux I__4167 (
            .O(N__22915),
            .I(N__22912));
    Span12Mux_v I__4166 (
            .O(N__22912),
            .I(N__22909));
    Odrv12 I__4165 (
            .O(N__22909),
            .I(\POWERLED.un34_clk_100khz_8 ));
    CascadeMux I__4164 (
            .O(N__22906),
            .I(\POWERLED.un34_clk_100khz_9_cascade_ ));
    InMux I__4163 (
            .O(N__22903),
            .I(N__22900));
    LocalMux I__4162 (
            .O(N__22900),
            .I(N__22897));
    Span4Mux_v I__4161 (
            .O(N__22897),
            .I(N__22894));
    Odrv4 I__4160 (
            .O(N__22894),
            .I(\POWERLED.un34_clk_100khz_11 ));
    InMux I__4159 (
            .O(N__22891),
            .I(N__22888));
    LocalMux I__4158 (
            .O(N__22888),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ));
    CascadeMux I__4157 (
            .O(N__22885),
            .I(\POWERLED.N_220_cascade_ ));
    InMux I__4156 (
            .O(N__22882),
            .I(N__22878));
    InMux I__4155 (
            .O(N__22881),
            .I(N__22875));
    LocalMux I__4154 (
            .O(N__22878),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823 ));
    LocalMux I__4153 (
            .O(N__22875),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823 ));
    CascadeMux I__4152 (
            .O(N__22870),
            .I(\POWERLED.N_304_cascade_ ));
    InMux I__4151 (
            .O(N__22867),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__4150 (
            .O(N__22864),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__4149 (
            .O(N__22861),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    InMux I__4148 (
            .O(N__22858),
            .I(bfn_8_5_0_));
    CascadeMux I__4147 (
            .O(N__22855),
            .I(\POWERLED.count_off_RNIBQDB2Z0Z_0_cascade_ ));
    CascadeMux I__4146 (
            .O(N__22852),
            .I(\POWERLED.count_offZ0Z_0_cascade_ ));
    CascadeMux I__4145 (
            .O(N__22849),
            .I(\POWERLED.count_off_RNIZ0Z_1_cascade_ ));
    CascadeMux I__4144 (
            .O(N__22846),
            .I(N__22843));
    InMux I__4143 (
            .O(N__22843),
            .I(N__22840));
    LocalMux I__4142 (
            .O(N__22840),
            .I(N__22834));
    InMux I__4141 (
            .O(N__22839),
            .I(N__22831));
    InMux I__4140 (
            .O(N__22838),
            .I(N__22826));
    InMux I__4139 (
            .O(N__22837),
            .I(N__22826));
    Span4Mux_h I__4138 (
            .O(N__22834),
            .I(N__22823));
    LocalMux I__4137 (
            .O(N__22831),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__4136 (
            .O(N__22826),
            .I(\POWERLED.count_offZ0Z_0 ));
    Odrv4 I__4135 (
            .O(N__22823),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__4134 (
            .O(N__22816),
            .I(N__22813));
    LocalMux I__4133 (
            .O(N__22813),
            .I(\POWERLED.count_off_0_0 ));
    InMux I__4132 (
            .O(N__22810),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__4131 (
            .O(N__22807),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__4130 (
            .O(N__22804),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__4129 (
            .O(N__22801),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__4128 (
            .O(N__22798),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    InMux I__4127 (
            .O(N__22795),
            .I(bfn_8_4_0_));
    InMux I__4126 (
            .O(N__22792),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__4125 (
            .O(N__22789),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__4124 (
            .O(N__22786),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    InMux I__4123 (
            .O(N__22783),
            .I(N__22777));
    InMux I__4122 (
            .O(N__22782),
            .I(N__22777));
    LocalMux I__4121 (
            .O(N__22777),
            .I(\PCH_PWRGD.count_rst_2 ));
    InMux I__4120 (
            .O(N__22774),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__4119 (
            .O(N__22771),
            .I(N__22768));
    LocalMux I__4118 (
            .O(N__22768),
            .I(\PCH_PWRGD.un2_count_1_axb_13 ));
    InMux I__4117 (
            .O(N__22765),
            .I(N__22758));
    InMux I__4116 (
            .O(N__22764),
            .I(N__22758));
    InMux I__4115 (
            .O(N__22763),
            .I(N__22755));
    LocalMux I__4114 (
            .O(N__22758),
            .I(\PCH_PWRGD.count_rst_1 ));
    LocalMux I__4113 (
            .O(N__22755),
            .I(\PCH_PWRGD.count_rst_1 ));
    InMux I__4112 (
            .O(N__22750),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    InMux I__4111 (
            .O(N__22747),
            .I(N__22744));
    LocalMux I__4110 (
            .O(N__22744),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__4109 (
            .O(N__22741),
            .I(N__22735));
    InMux I__4108 (
            .O(N__22740),
            .I(N__22735));
    LocalMux I__4107 (
            .O(N__22735),
            .I(N__22732));
    Odrv4 I__4106 (
            .O(N__22732),
            .I(\PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ));
    InMux I__4105 (
            .O(N__22729),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__4104 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__4103 (
            .O(N__22723),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    InMux I__4102 (
            .O(N__22720),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__4101 (
            .O(N__22717),
            .I(N__22711));
    InMux I__4100 (
            .O(N__22716),
            .I(N__22711));
    LocalMux I__4099 (
            .O(N__22711),
            .I(\PCH_PWRGD.count_rst ));
    InMux I__4098 (
            .O(N__22708),
            .I(N__22704));
    InMux I__4097 (
            .O(N__22707),
            .I(N__22701));
    LocalMux I__4096 (
            .O(N__22704),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__4095 (
            .O(N__22701),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    InMux I__4094 (
            .O(N__22696),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__4093 (
            .O(N__22693),
            .I(N__22689));
    InMux I__4092 (
            .O(N__22692),
            .I(N__22686));
    LocalMux I__4091 (
            .O(N__22689),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__4090 (
            .O(N__22686),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__4089 (
            .O(N__22681),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    InMux I__4088 (
            .O(N__22678),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    CascadeMux I__4087 (
            .O(N__22675),
            .I(N__22672));
    InMux I__4086 (
            .O(N__22672),
            .I(N__22668));
    InMux I__4085 (
            .O(N__22671),
            .I(N__22665));
    LocalMux I__4084 (
            .O(N__22668),
            .I(\PCH_PWRGD.un2_count_1_axb_4 ));
    LocalMux I__4083 (
            .O(N__22665),
            .I(\PCH_PWRGD.un2_count_1_axb_4 ));
    InMux I__4082 (
            .O(N__22660),
            .I(N__22654));
    InMux I__4081 (
            .O(N__22659),
            .I(N__22654));
    LocalMux I__4080 (
            .O(N__22654),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__4079 (
            .O(N__22651),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    InMux I__4078 (
            .O(N__22648),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    InMux I__4077 (
            .O(N__22645),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    InMux I__4076 (
            .O(N__22642),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    InMux I__4075 (
            .O(N__22639),
            .I(\PCH_PWRGD.un2_count_1_cry_7 ));
    InMux I__4074 (
            .O(N__22636),
            .I(bfn_8_2_0_));
    InMux I__4073 (
            .O(N__22633),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    InMux I__4072 (
            .O(N__22630),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__4071 (
            .O(N__22627),
            .I(N__22624));
    LocalMux I__4070 (
            .O(N__22624),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    CascadeMux I__4069 (
            .O(N__22621),
            .I(N__22618));
    InMux I__4068 (
            .O(N__22618),
            .I(N__22615));
    LocalMux I__4067 (
            .O(N__22615),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__4066 (
            .O(N__22612),
            .I(N__22609));
    LocalMux I__4065 (
            .O(N__22609),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    CascadeMux I__4064 (
            .O(N__22606),
            .I(N__22603));
    InMux I__4063 (
            .O(N__22603),
            .I(N__22593));
    InMux I__4062 (
            .O(N__22602),
            .I(N__22593));
    InMux I__4061 (
            .O(N__22601),
            .I(N__22593));
    InMux I__4060 (
            .O(N__22600),
            .I(N__22590));
    LocalMux I__4059 (
            .O(N__22593),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__4058 (
            .O(N__22590),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__4057 (
            .O(N__22585),
            .I(N__22581));
    InMux I__4056 (
            .O(N__22584),
            .I(N__22573));
    InMux I__4055 (
            .O(N__22581),
            .I(N__22573));
    InMux I__4054 (
            .O(N__22580),
            .I(N__22573));
    LocalMux I__4053 (
            .O(N__22573),
            .I(G_2078));
    CascadeMux I__4052 (
            .O(N__22570),
            .I(N__22567));
    InMux I__4051 (
            .O(N__22567),
            .I(N__22564));
    LocalMux I__4050 (
            .O(N__22564),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__4049 (
            .O(N__22561),
            .I(N__22558));
    LocalMux I__4048 (
            .O(N__22558),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__4047 (
            .O(N__22555),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    InMux I__4046 (
            .O(N__22552),
            .I(N__22549));
    LocalMux I__4045 (
            .O(N__22549),
            .I(N__22546));
    Span4Mux_v I__4044 (
            .O(N__22546),
            .I(N__22543));
    Span4Mux_h I__4043 (
            .O(N__22543),
            .I(N__22540));
    Odrv4 I__4042 (
            .O(N__22540),
            .I(\POWERLED.un85_clk_100khz_0 ));
    IoInMux I__4041 (
            .O(N__22537),
            .I(N__22534));
    LocalMux I__4040 (
            .O(N__22534),
            .I(G_9));
    InMux I__4039 (
            .O(N__22531),
            .I(N__22528));
    LocalMux I__4038 (
            .O(N__22528),
            .I(\PCH_PWRGD.un2_count_1_axb_2 ));
    InMux I__4037 (
            .O(N__22525),
            .I(N__22516));
    InMux I__4036 (
            .O(N__22524),
            .I(N__22516));
    InMux I__4035 (
            .O(N__22523),
            .I(N__22516));
    LocalMux I__4034 (
            .O(N__22516),
            .I(\PCH_PWRGD.count_rst_12 ));
    InMux I__4033 (
            .O(N__22513),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    CascadeMux I__4032 (
            .O(N__22510),
            .I(N__22507));
    InMux I__4031 (
            .O(N__22507),
            .I(N__22504));
    LocalMux I__4030 (
            .O(N__22504),
            .I(N__22501));
    Span4Mux_v I__4029 (
            .O(N__22501),
            .I(N__22498));
    Odrv4 I__4028 (
            .O(N__22498),
            .I(\POWERLED.mult1_un152_sum_i ));
    InMux I__4027 (
            .O(N__22495),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__4026 (
            .O(N__22492),
            .I(N__22489));
    LocalMux I__4025 (
            .O(N__22489),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__4024 (
            .O(N__22486),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    CascadeMux I__4023 (
            .O(N__22483),
            .I(N__22480));
    InMux I__4022 (
            .O(N__22480),
            .I(N__22477));
    LocalMux I__4021 (
            .O(N__22477),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__4020 (
            .O(N__22474),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__4019 (
            .O(N__22471),
            .I(N__22468));
    LocalMux I__4018 (
            .O(N__22468),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    CascadeMux I__4017 (
            .O(N__22465),
            .I(N__22462));
    InMux I__4016 (
            .O(N__22462),
            .I(N__22454));
    InMux I__4015 (
            .O(N__22461),
            .I(N__22454));
    InMux I__4014 (
            .O(N__22460),
            .I(N__22451));
    InMux I__4013 (
            .O(N__22459),
            .I(N__22448));
    LocalMux I__4012 (
            .O(N__22454),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__4011 (
            .O(N__22451),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__4010 (
            .O(N__22448),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    InMux I__4009 (
            .O(N__22441),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    CascadeMux I__4008 (
            .O(N__22438),
            .I(N__22434));
    InMux I__4007 (
            .O(N__22437),
            .I(N__22426));
    InMux I__4006 (
            .O(N__22434),
            .I(N__22426));
    InMux I__4005 (
            .O(N__22433),
            .I(N__22426));
    LocalMux I__4004 (
            .O(N__22426),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    CascadeMux I__4003 (
            .O(N__22423),
            .I(N__22420));
    InMux I__4002 (
            .O(N__22420),
            .I(N__22417));
    LocalMux I__4001 (
            .O(N__22417),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__4000 (
            .O(N__22414),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__3999 (
            .O(N__22411),
            .I(N__22408));
    LocalMux I__3998 (
            .O(N__22408),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__3997 (
            .O(N__22405),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__3996 (
            .O(N__22402),
            .I(\POWERLED.mult1_un159_sum_s_7_cascade_ ));
    InMux I__3995 (
            .O(N__22399),
            .I(N__22396));
    LocalMux I__3994 (
            .O(N__22396),
            .I(N__22393));
    Span4Mux_v I__3993 (
            .O(N__22393),
            .I(N__22390));
    Span4Mux_h I__3992 (
            .O(N__22390),
            .I(N__22387));
    Odrv4 I__3991 (
            .O(N__22387),
            .I(\POWERLED.un85_clk_100khz_1 ));
    CascadeMux I__3990 (
            .O(N__22384),
            .I(N__22379));
    InMux I__3989 (
            .O(N__22383),
            .I(N__22373));
    InMux I__3988 (
            .O(N__22382),
            .I(N__22370));
    InMux I__3987 (
            .O(N__22379),
            .I(N__22367));
    InMux I__3986 (
            .O(N__22378),
            .I(N__22361));
    InMux I__3985 (
            .O(N__22377),
            .I(N__22361));
    CascadeMux I__3984 (
            .O(N__22376),
            .I(N__22358));
    LocalMux I__3983 (
            .O(N__22373),
            .I(N__22353));
    LocalMux I__3982 (
            .O(N__22370),
            .I(N__22350));
    LocalMux I__3981 (
            .O(N__22367),
            .I(N__22347));
    InMux I__3980 (
            .O(N__22366),
            .I(N__22344));
    LocalMux I__3979 (
            .O(N__22361),
            .I(N__22339));
    InMux I__3978 (
            .O(N__22358),
            .I(N__22334));
    InMux I__3977 (
            .O(N__22357),
            .I(N__22334));
    CascadeMux I__3976 (
            .O(N__22356),
            .I(N__22331));
    Span4Mux_v I__3975 (
            .O(N__22353),
            .I(N__22328));
    Span4Mux_h I__3974 (
            .O(N__22350),
            .I(N__22323));
    Span4Mux_v I__3973 (
            .O(N__22347),
            .I(N__22323));
    LocalMux I__3972 (
            .O(N__22344),
            .I(N__22319));
    InMux I__3971 (
            .O(N__22343),
            .I(N__22314));
    InMux I__3970 (
            .O(N__22342),
            .I(N__22314));
    Span4Mux_v I__3969 (
            .O(N__22339),
            .I(N__22309));
    LocalMux I__3968 (
            .O(N__22334),
            .I(N__22309));
    InMux I__3967 (
            .O(N__22331),
            .I(N__22306));
    Span4Mux_h I__3966 (
            .O(N__22328),
            .I(N__22301));
    Span4Mux_v I__3965 (
            .O(N__22323),
            .I(N__22301));
    InMux I__3964 (
            .O(N__22322),
            .I(N__22298));
    Span12Mux_s4_v I__3963 (
            .O(N__22319),
            .I(N__22289));
    LocalMux I__3962 (
            .O(N__22314),
            .I(N__22289));
    Sp12to4 I__3961 (
            .O(N__22309),
            .I(N__22289));
    LocalMux I__3960 (
            .O(N__22306),
            .I(N__22289));
    Odrv4 I__3959 (
            .O(N__22301),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__3958 (
            .O(N__22298),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv12 I__3957 (
            .O(N__22289),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    CascadeMux I__3956 (
            .O(N__22282),
            .I(N__22279));
    InMux I__3955 (
            .O(N__22279),
            .I(N__22276));
    LocalMux I__3954 (
            .O(N__22276),
            .I(N__22273));
    Span12Mux_s8_h I__3953 (
            .O(N__22273),
            .I(N__22270));
    Odrv12 I__3952 (
            .O(N__22270),
            .I(\POWERLED.mult1_un159_sum_i ));
    InMux I__3951 (
            .O(N__22267),
            .I(N__22264));
    LocalMux I__3950 (
            .O(N__22264),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__3949 (
            .O(N__22261),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    CascadeMux I__3948 (
            .O(N__22258),
            .I(N__22255));
    InMux I__3947 (
            .O(N__22255),
            .I(N__22252));
    LocalMux I__3946 (
            .O(N__22252),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__3945 (
            .O(N__22249),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    InMux I__3944 (
            .O(N__22246),
            .I(N__22243));
    LocalMux I__3943 (
            .O(N__22243),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__3942 (
            .O(N__22240),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__3941 (
            .O(N__22237),
            .I(N__22234));
    LocalMux I__3940 (
            .O(N__22234),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__3939 (
            .O(N__22231),
            .I(N__22228));
    LocalMux I__3938 (
            .O(N__22228),
            .I(N__22225));
    Span4Mux_s2_v I__3937 (
            .O(N__22225),
            .I(N__22220));
    CascadeMux I__3936 (
            .O(N__22224),
            .I(N__22217));
    CascadeMux I__3935 (
            .O(N__22223),
            .I(N__22214));
    Span4Mux_h I__3934 (
            .O(N__22220),
            .I(N__22210));
    InMux I__3933 (
            .O(N__22217),
            .I(N__22207));
    InMux I__3932 (
            .O(N__22214),
            .I(N__22204));
    InMux I__3931 (
            .O(N__22213),
            .I(N__22201));
    Odrv4 I__3930 (
            .O(N__22210),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3929 (
            .O(N__22207),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3928 (
            .O(N__22204),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__3927 (
            .O(N__22201),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    InMux I__3926 (
            .O(N__22192),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    InMux I__3925 (
            .O(N__22189),
            .I(N__22186));
    LocalMux I__3924 (
            .O(N__22186),
            .I(N__22183));
    Odrv4 I__3923 (
            .O(N__22183),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    CascadeMux I__3922 (
            .O(N__22180),
            .I(N__22176));
    CascadeMux I__3921 (
            .O(N__22179),
            .I(N__22172));
    InMux I__3920 (
            .O(N__22176),
            .I(N__22165));
    InMux I__3919 (
            .O(N__22175),
            .I(N__22165));
    InMux I__3918 (
            .O(N__22172),
            .I(N__22165));
    LocalMux I__3917 (
            .O(N__22165),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    InMux I__3916 (
            .O(N__22162),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__3915 (
            .O(N__22159),
            .I(N__22156));
    LocalMux I__3914 (
            .O(N__22156),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__3913 (
            .O(N__22153),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__3912 (
            .O(N__22150),
            .I(\POWERLED.mult1_un152_sum_s_8_cascade_ ));
    InMux I__3911 (
            .O(N__22147),
            .I(N__22136));
    InMux I__3910 (
            .O(N__22146),
            .I(N__22133));
    CascadeMux I__3909 (
            .O(N__22145),
            .I(N__22130));
    InMux I__3908 (
            .O(N__22144),
            .I(N__22126));
    InMux I__3907 (
            .O(N__22143),
            .I(N__22121));
    InMux I__3906 (
            .O(N__22142),
            .I(N__22121));
    InMux I__3905 (
            .O(N__22141),
            .I(N__22118));
    InMux I__3904 (
            .O(N__22140),
            .I(N__22113));
    InMux I__3903 (
            .O(N__22139),
            .I(N__22113));
    LocalMux I__3902 (
            .O(N__22136),
            .I(N__22107));
    LocalMux I__3901 (
            .O(N__22133),
            .I(N__22107));
    InMux I__3900 (
            .O(N__22130),
            .I(N__22103));
    InMux I__3899 (
            .O(N__22129),
            .I(N__22100));
    LocalMux I__3898 (
            .O(N__22126),
            .I(N__22095));
    LocalMux I__3897 (
            .O(N__22121),
            .I(N__22095));
    LocalMux I__3896 (
            .O(N__22118),
            .I(N__22090));
    LocalMux I__3895 (
            .O(N__22113),
            .I(N__22087));
    CascadeMux I__3894 (
            .O(N__22112),
            .I(N__22083));
    Sp12to4 I__3893 (
            .O(N__22107),
            .I(N__22080));
    CascadeMux I__3892 (
            .O(N__22106),
            .I(N__22077));
    LocalMux I__3891 (
            .O(N__22103),
            .I(N__22074));
    LocalMux I__3890 (
            .O(N__22100),
            .I(N__22069));
    Span4Mux_v I__3889 (
            .O(N__22095),
            .I(N__22069));
    InMux I__3888 (
            .O(N__22094),
            .I(N__22064));
    InMux I__3887 (
            .O(N__22093),
            .I(N__22064));
    Span4Mux_v I__3886 (
            .O(N__22090),
            .I(N__22059));
    Span4Mux_s2_h I__3885 (
            .O(N__22087),
            .I(N__22059));
    InMux I__3884 (
            .O(N__22086),
            .I(N__22056));
    InMux I__3883 (
            .O(N__22083),
            .I(N__22053));
    Span12Mux_v I__3882 (
            .O(N__22080),
            .I(N__22050));
    InMux I__3881 (
            .O(N__22077),
            .I(N__22047));
    Span4Mux_v I__3880 (
            .O(N__22074),
            .I(N__22044));
    Span4Mux_v I__3879 (
            .O(N__22069),
            .I(N__22033));
    LocalMux I__3878 (
            .O(N__22064),
            .I(N__22033));
    Span4Mux_h I__3877 (
            .O(N__22059),
            .I(N__22033));
    LocalMux I__3876 (
            .O(N__22056),
            .I(N__22033));
    LocalMux I__3875 (
            .O(N__22053),
            .I(N__22033));
    Odrv12 I__3874 (
            .O(N__22050),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__3873 (
            .O(N__22047),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__3872 (
            .O(N__22044),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__3871 (
            .O(N__22033),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    CascadeMux I__3870 (
            .O(N__22024),
            .I(G_155_cascade_));
    InMux I__3869 (
            .O(N__22021),
            .I(N__22018));
    LocalMux I__3868 (
            .O(N__22018),
            .I(\POWERLED.N_73 ));
    InMux I__3867 (
            .O(N__22015),
            .I(N__22009));
    InMux I__3866 (
            .O(N__22014),
            .I(N__22009));
    LocalMux I__3865 (
            .O(N__22009),
            .I(\POWERLED.dutycycle_eena_1 ));
    CascadeMux I__3864 (
            .O(N__22006),
            .I(\POWERLED.N_73_cascade_ ));
    InMux I__3863 (
            .O(N__22003),
            .I(N__21997));
    InMux I__3862 (
            .O(N__22002),
            .I(N__21997));
    LocalMux I__3861 (
            .O(N__21997),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    CascadeMux I__3860 (
            .O(N__21994),
            .I(N__21991));
    InMux I__3859 (
            .O(N__21991),
            .I(N__21988));
    LocalMux I__3858 (
            .O(N__21988),
            .I(\POWERLED.N_277 ));
    InMux I__3857 (
            .O(N__21985),
            .I(N__21982));
    LocalMux I__3856 (
            .O(N__21982),
            .I(N__21979));
    Odrv12 I__3855 (
            .O(N__21979),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ));
    InMux I__3854 (
            .O(N__21976),
            .I(N__21973));
    LocalMux I__3853 (
            .O(N__21973),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_2 ));
    CascadeMux I__3852 (
            .O(N__21970),
            .I(\POWERLED.dutycycle_1_0_iv_0_1_5_cascade_ ));
    InMux I__3851 (
            .O(N__21967),
            .I(N__21958));
    InMux I__3850 (
            .O(N__21966),
            .I(N__21958));
    InMux I__3849 (
            .O(N__21965),
            .I(N__21958));
    LocalMux I__3848 (
            .O(N__21958),
            .I(SUSWARN_N_fast));
    InMux I__3847 (
            .O(N__21955),
            .I(N__21946));
    CascadeMux I__3846 (
            .O(N__21954),
            .I(N__21943));
    InMux I__3845 (
            .O(N__21953),
            .I(N__21940));
    InMux I__3844 (
            .O(N__21952),
            .I(N__21936));
    CascadeMux I__3843 (
            .O(N__21951),
            .I(N__21933));
    InMux I__3842 (
            .O(N__21950),
            .I(N__21930));
    InMux I__3841 (
            .O(N__21949),
            .I(N__21927));
    LocalMux I__3840 (
            .O(N__21946),
            .I(N__21922));
    InMux I__3839 (
            .O(N__21943),
            .I(N__21919));
    LocalMux I__3838 (
            .O(N__21940),
            .I(N__21916));
    InMux I__3837 (
            .O(N__21939),
            .I(N__21913));
    LocalMux I__3836 (
            .O(N__21936),
            .I(N__21910));
    InMux I__3835 (
            .O(N__21933),
            .I(N__21907));
    LocalMux I__3834 (
            .O(N__21930),
            .I(N__21904));
    LocalMux I__3833 (
            .O(N__21927),
            .I(N__21901));
    CascadeMux I__3832 (
            .O(N__21926),
            .I(N__21897));
    InMux I__3831 (
            .O(N__21925),
            .I(N__21885));
    Span4Mux_h I__3830 (
            .O(N__21922),
            .I(N__21880));
    LocalMux I__3829 (
            .O(N__21919),
            .I(N__21880));
    Span4Mux_v I__3828 (
            .O(N__21916),
            .I(N__21875));
    LocalMux I__3827 (
            .O(N__21913),
            .I(N__21875));
    Span4Mux_v I__3826 (
            .O(N__21910),
            .I(N__21870));
    LocalMux I__3825 (
            .O(N__21907),
            .I(N__21870));
    Span4Mux_v I__3824 (
            .O(N__21904),
            .I(N__21865));
    Span4Mux_v I__3823 (
            .O(N__21901),
            .I(N__21865));
    InMux I__3822 (
            .O(N__21900),
            .I(N__21858));
    InMux I__3821 (
            .O(N__21897),
            .I(N__21858));
    InMux I__3820 (
            .O(N__21896),
            .I(N__21858));
    InMux I__3819 (
            .O(N__21895),
            .I(N__21847));
    InMux I__3818 (
            .O(N__21894),
            .I(N__21847));
    InMux I__3817 (
            .O(N__21893),
            .I(N__21847));
    InMux I__3816 (
            .O(N__21892),
            .I(N__21847));
    InMux I__3815 (
            .O(N__21891),
            .I(N__21847));
    InMux I__3814 (
            .O(N__21890),
            .I(N__21840));
    InMux I__3813 (
            .O(N__21889),
            .I(N__21840));
    InMux I__3812 (
            .O(N__21888),
            .I(N__21840));
    LocalMux I__3811 (
            .O(N__21885),
            .I(N__21835));
    Span4Mux_h I__3810 (
            .O(N__21880),
            .I(N__21835));
    Odrv4 I__3809 (
            .O(N__21875),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__3808 (
            .O(N__21870),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__3807 (
            .O(N__21865),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__3806 (
            .O(N__21858),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__3805 (
            .O(N__21847),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__3804 (
            .O(N__21840),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__3803 (
            .O(N__21835),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__3802 (
            .O(N__21820),
            .I(N__21817));
    LocalMux I__3801 (
            .O(N__21817),
            .I(\POWERLED.m18_e_0 ));
    CascadeMux I__3800 (
            .O(N__21814),
            .I(N__21810));
    CascadeMux I__3799 (
            .O(N__21813),
            .I(N__21797));
    InMux I__3798 (
            .O(N__21810),
            .I(N__21793));
    InMux I__3797 (
            .O(N__21809),
            .I(N__21788));
    InMux I__3796 (
            .O(N__21808),
            .I(N__21788));
    InMux I__3795 (
            .O(N__21807),
            .I(N__21785));
    CascadeMux I__3794 (
            .O(N__21806),
            .I(N__21781));
    InMux I__3793 (
            .O(N__21805),
            .I(N__21778));
    CascadeMux I__3792 (
            .O(N__21804),
            .I(N__21772));
    InMux I__3791 (
            .O(N__21803),
            .I(N__21767));
    InMux I__3790 (
            .O(N__21802),
            .I(N__21767));
    CascadeMux I__3789 (
            .O(N__21801),
            .I(N__21763));
    CascadeMux I__3788 (
            .O(N__21800),
            .I(N__21759));
    InMux I__3787 (
            .O(N__21797),
            .I(N__21756));
    InMux I__3786 (
            .O(N__21796),
            .I(N__21753));
    LocalMux I__3785 (
            .O(N__21793),
            .I(N__21750));
    LocalMux I__3784 (
            .O(N__21788),
            .I(N__21747));
    LocalMux I__3783 (
            .O(N__21785),
            .I(N__21744));
    InMux I__3782 (
            .O(N__21784),
            .I(N__21741));
    InMux I__3781 (
            .O(N__21781),
            .I(N__21738));
    LocalMux I__3780 (
            .O(N__21778),
            .I(N__21735));
    InMux I__3779 (
            .O(N__21777),
            .I(N__21730));
    InMux I__3778 (
            .O(N__21776),
            .I(N__21730));
    InMux I__3777 (
            .O(N__21775),
            .I(N__21723));
    InMux I__3776 (
            .O(N__21772),
            .I(N__21723));
    LocalMux I__3775 (
            .O(N__21767),
            .I(N__21720));
    InMux I__3774 (
            .O(N__21766),
            .I(N__21711));
    InMux I__3773 (
            .O(N__21763),
            .I(N__21711));
    InMux I__3772 (
            .O(N__21762),
            .I(N__21711));
    InMux I__3771 (
            .O(N__21759),
            .I(N__21711));
    LocalMux I__3770 (
            .O(N__21756),
            .I(N__21708));
    LocalMux I__3769 (
            .O(N__21753),
            .I(N__21705));
    Span4Mux_h I__3768 (
            .O(N__21750),
            .I(N__21694));
    Span4Mux_v I__3767 (
            .O(N__21747),
            .I(N__21694));
    Span4Mux_h I__3766 (
            .O(N__21744),
            .I(N__21694));
    LocalMux I__3765 (
            .O(N__21741),
            .I(N__21694));
    LocalMux I__3764 (
            .O(N__21738),
            .I(N__21694));
    Span4Mux_v I__3763 (
            .O(N__21735),
            .I(N__21689));
    LocalMux I__3762 (
            .O(N__21730),
            .I(N__21689));
    InMux I__3761 (
            .O(N__21729),
            .I(N__21684));
    InMux I__3760 (
            .O(N__21728),
            .I(N__21684));
    LocalMux I__3759 (
            .O(N__21723),
            .I(N__21681));
    Span4Mux_h I__3758 (
            .O(N__21720),
            .I(N__21676));
    LocalMux I__3757 (
            .O(N__21711),
            .I(N__21676));
    Odrv4 I__3756 (
            .O(N__21708),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3755 (
            .O(N__21705),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3754 (
            .O(N__21694),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3753 (
            .O(N__21689),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__3752 (
            .O(N__21684),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3751 (
            .O(N__21681),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3750 (
            .O(N__21676),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    InMux I__3749 (
            .O(N__21661),
            .I(N__21658));
    LocalMux I__3748 (
            .O(N__21658),
            .I(\POWERLED.un1_dutycycle_94_cry_4_c_RNI919HZ0Z1 ));
    CascadeMux I__3747 (
            .O(N__21655),
            .I(\POWERLED.dutycycle_1_0_5_cascade_ ));
    InMux I__3746 (
            .O(N__21652),
            .I(N__21648));
    InMux I__3745 (
            .O(N__21651),
            .I(N__21645));
    LocalMux I__3744 (
            .O(N__21648),
            .I(\POWERLED.func_state_RNIT69J5Z0Z_1 ));
    LocalMux I__3743 (
            .O(N__21645),
            .I(\POWERLED.func_state_RNIT69J5Z0Z_1 ));
    CascadeMux I__3742 (
            .O(N__21640),
            .I(\POWERLED.N_366_cascade_ ));
    CascadeMux I__3741 (
            .O(N__21637),
            .I(\POWERLED.dutycycle_RNI2O4A1Z0Z_6_cascade_ ));
    InMux I__3740 (
            .O(N__21634),
            .I(N__21631));
    LocalMux I__3739 (
            .O(N__21631),
            .I(\POWERLED.dutycycle_RNI2O4A1_2Z0Z_2 ));
    CascadeMux I__3738 (
            .O(N__21628),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m1_cascade_ ));
    InMux I__3737 (
            .O(N__21625),
            .I(N__21622));
    LocalMux I__3736 (
            .O(N__21622),
            .I(N__21617));
    InMux I__3735 (
            .O(N__21621),
            .I(N__21612));
    InMux I__3734 (
            .O(N__21620),
            .I(N__21612));
    Span4Mux_v I__3733 (
            .O(N__21617),
            .I(N__21607));
    LocalMux I__3732 (
            .O(N__21612),
            .I(N__21607));
    Odrv4 I__3731 (
            .O(N__21607),
            .I(\POWERLED.dutycycle_RNIZ0Z_5 ));
    CascadeMux I__3730 (
            .O(N__21604),
            .I(\POWERLED.func_state_RNI_0Z0Z_0_cascade_ ));
    InMux I__3729 (
            .O(N__21601),
            .I(N__21598));
    LocalMux I__3728 (
            .O(N__21598),
            .I(\POWERLED.func_state_RNI68EU3Z0Z_1 ));
    InMux I__3727 (
            .O(N__21595),
            .I(N__21592));
    LocalMux I__3726 (
            .O(N__21592),
            .I(N__21589));
    Span4Mux_h I__3725 (
            .O(N__21589),
            .I(N__21586));
    Odrv4 I__3724 (
            .O(N__21586),
            .I(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ));
    InMux I__3723 (
            .O(N__21583),
            .I(N__21577));
    InMux I__3722 (
            .O(N__21582),
            .I(N__21577));
    LocalMux I__3721 (
            .O(N__21577),
            .I(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ));
    InMux I__3720 (
            .O(N__21574),
            .I(\POWERLED.un1_dutycycle_94_cry_10 ));
    InMux I__3719 (
            .O(N__21571),
            .I(\POWERLED.un1_dutycycle_94_cry_11 ));
    InMux I__3718 (
            .O(N__21568),
            .I(N__21563));
    InMux I__3717 (
            .O(N__21567),
            .I(N__21559));
    InMux I__3716 (
            .O(N__21566),
            .I(N__21556));
    LocalMux I__3715 (
            .O(N__21563),
            .I(N__21552));
    CascadeMux I__3714 (
            .O(N__21562),
            .I(N__21548));
    LocalMux I__3713 (
            .O(N__21559),
            .I(N__21544));
    LocalMux I__3712 (
            .O(N__21556),
            .I(N__21541));
    InMux I__3711 (
            .O(N__21555),
            .I(N__21538));
    Span4Mux_v I__3710 (
            .O(N__21552),
            .I(N__21535));
    InMux I__3709 (
            .O(N__21551),
            .I(N__21530));
    InMux I__3708 (
            .O(N__21548),
            .I(N__21530));
    CascadeMux I__3707 (
            .O(N__21547),
            .I(N__21525));
    Span4Mux_v I__3706 (
            .O(N__21544),
            .I(N__21518));
    Span4Mux_v I__3705 (
            .O(N__21541),
            .I(N__21518));
    LocalMux I__3704 (
            .O(N__21538),
            .I(N__21518));
    Span4Mux_h I__3703 (
            .O(N__21535),
            .I(N__21513));
    LocalMux I__3702 (
            .O(N__21530),
            .I(N__21513));
    InMux I__3701 (
            .O(N__21529),
            .I(N__21510));
    InMux I__3700 (
            .O(N__21528),
            .I(N__21507));
    InMux I__3699 (
            .O(N__21525),
            .I(N__21504));
    Odrv4 I__3698 (
            .O(N__21518),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__3697 (
            .O(N__21513),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3696 (
            .O(N__21510),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3695 (
            .O(N__21507),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3694 (
            .O(N__21504),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    InMux I__3693 (
            .O(N__21493),
            .I(N__21487));
    InMux I__3692 (
            .O(N__21492),
            .I(N__21487));
    LocalMux I__3691 (
            .O(N__21487),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    InMux I__3690 (
            .O(N__21484),
            .I(\POWERLED.un1_dutycycle_94_cry_12 ));
    InMux I__3689 (
            .O(N__21481),
            .I(N__21475));
    InMux I__3688 (
            .O(N__21480),
            .I(N__21475));
    LocalMux I__3687 (
            .O(N__21475),
            .I(N__21472));
    Odrv4 I__3686 (
            .O(N__21472),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    InMux I__3685 (
            .O(N__21469),
            .I(\POWERLED.un1_dutycycle_94_cry_13 ));
    InMux I__3684 (
            .O(N__21466),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    InMux I__3683 (
            .O(N__21463),
            .I(N__21457));
    InMux I__3682 (
            .O(N__21462),
            .I(N__21457));
    LocalMux I__3681 (
            .O(N__21457),
            .I(N__21454));
    Odrv4 I__3680 (
            .O(N__21454),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    InMux I__3679 (
            .O(N__21451),
            .I(N__21446));
    CascadeMux I__3678 (
            .O(N__21450),
            .I(N__21443));
    CascadeMux I__3677 (
            .O(N__21449),
            .I(N__21440));
    LocalMux I__3676 (
            .O(N__21446),
            .I(N__21435));
    InMux I__3675 (
            .O(N__21443),
            .I(N__21430));
    InMux I__3674 (
            .O(N__21440),
            .I(N__21427));
    InMux I__3673 (
            .O(N__21439),
            .I(N__21424));
    CascadeMux I__3672 (
            .O(N__21438),
            .I(N__21421));
    Span4Mux_v I__3671 (
            .O(N__21435),
            .I(N__21418));
    InMux I__3670 (
            .O(N__21434),
            .I(N__21415));
    InMux I__3669 (
            .O(N__21433),
            .I(N__21412));
    LocalMux I__3668 (
            .O(N__21430),
            .I(N__21409));
    LocalMux I__3667 (
            .O(N__21427),
            .I(N__21404));
    LocalMux I__3666 (
            .O(N__21424),
            .I(N__21404));
    InMux I__3665 (
            .O(N__21421),
            .I(N__21401));
    Odrv4 I__3664 (
            .O(N__21418),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3663 (
            .O(N__21415),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3662 (
            .O(N__21412),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv12 I__3661 (
            .O(N__21409),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__3660 (
            .O(N__21404),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3659 (
            .O(N__21401),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    CascadeMux I__3658 (
            .O(N__21388),
            .I(N__21382));
    CascadeMux I__3657 (
            .O(N__21387),
            .I(N__21377));
    InMux I__3656 (
            .O(N__21386),
            .I(N__21374));
    InMux I__3655 (
            .O(N__21385),
            .I(N__21369));
    InMux I__3654 (
            .O(N__21382),
            .I(N__21369));
    InMux I__3653 (
            .O(N__21381),
            .I(N__21362));
    InMux I__3652 (
            .O(N__21380),
            .I(N__21362));
    InMux I__3651 (
            .O(N__21377),
            .I(N__21362));
    LocalMux I__3650 (
            .O(N__21374),
            .I(N__21355));
    LocalMux I__3649 (
            .O(N__21369),
            .I(N__21352));
    LocalMux I__3648 (
            .O(N__21362),
            .I(N__21349));
    InMux I__3647 (
            .O(N__21361),
            .I(N__21340));
    InMux I__3646 (
            .O(N__21360),
            .I(N__21340));
    InMux I__3645 (
            .O(N__21359),
            .I(N__21340));
    InMux I__3644 (
            .O(N__21358),
            .I(N__21340));
    Span4Mux_h I__3643 (
            .O(N__21355),
            .I(N__21335));
    Span4Mux_h I__3642 (
            .O(N__21352),
            .I(N__21335));
    Odrv12 I__3641 (
            .O(N__21349),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    LocalMux I__3640 (
            .O(N__21340),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    Odrv4 I__3639 (
            .O(N__21335),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    InMux I__3638 (
            .O(N__21328),
            .I(N__21322));
    InMux I__3637 (
            .O(N__21327),
            .I(N__21322));
    LocalMux I__3636 (
            .O(N__21322),
            .I(N__21319));
    Odrv12 I__3635 (
            .O(N__21319),
            .I(\POWERLED.N_115_f0_1 ));
    CascadeMux I__3634 (
            .O(N__21316),
            .I(N__21311));
    CascadeMux I__3633 (
            .O(N__21315),
            .I(N__21308));
    InMux I__3632 (
            .O(N__21314),
            .I(N__21302));
    InMux I__3631 (
            .O(N__21311),
            .I(N__21302));
    InMux I__3630 (
            .O(N__21308),
            .I(N__21293));
    InMux I__3629 (
            .O(N__21307),
            .I(N__21290));
    LocalMux I__3628 (
            .O(N__21302),
            .I(N__21287));
    CascadeMux I__3627 (
            .O(N__21301),
            .I(N__21284));
    InMux I__3626 (
            .O(N__21300),
            .I(N__21281));
    InMux I__3625 (
            .O(N__21299),
            .I(N__21275));
    InMux I__3624 (
            .O(N__21298),
            .I(N__21268));
    InMux I__3623 (
            .O(N__21297),
            .I(N__21268));
    InMux I__3622 (
            .O(N__21296),
            .I(N__21268));
    LocalMux I__3621 (
            .O(N__21293),
            .I(N__21264));
    LocalMux I__3620 (
            .O(N__21290),
            .I(N__21259));
    Span4Mux_v I__3619 (
            .O(N__21287),
            .I(N__21259));
    InMux I__3618 (
            .O(N__21284),
            .I(N__21256));
    LocalMux I__3617 (
            .O(N__21281),
            .I(N__21253));
    InMux I__3616 (
            .O(N__21280),
            .I(N__21250));
    CascadeMux I__3615 (
            .O(N__21279),
            .I(N__21246));
    CascadeMux I__3614 (
            .O(N__21278),
            .I(N__21243));
    LocalMux I__3613 (
            .O(N__21275),
            .I(N__21237));
    LocalMux I__3612 (
            .O(N__21268),
            .I(N__21234));
    InMux I__3611 (
            .O(N__21267),
            .I(N__21231));
    Span4Mux_h I__3610 (
            .O(N__21264),
            .I(N__21228));
    Span4Mux_h I__3609 (
            .O(N__21259),
            .I(N__21223));
    LocalMux I__3608 (
            .O(N__21256),
            .I(N__21223));
    Span4Mux_h I__3607 (
            .O(N__21253),
            .I(N__21218));
    LocalMux I__3606 (
            .O(N__21250),
            .I(N__21218));
    InMux I__3605 (
            .O(N__21249),
            .I(N__21213));
    InMux I__3604 (
            .O(N__21246),
            .I(N__21213));
    InMux I__3603 (
            .O(N__21243),
            .I(N__21204));
    InMux I__3602 (
            .O(N__21242),
            .I(N__21204));
    InMux I__3601 (
            .O(N__21241),
            .I(N__21204));
    InMux I__3600 (
            .O(N__21240),
            .I(N__21204));
    Span4Mux_h I__3599 (
            .O(N__21237),
            .I(N__21199));
    Span4Mux_v I__3598 (
            .O(N__21234),
            .I(N__21199));
    LocalMux I__3597 (
            .O(N__21231),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__3596 (
            .O(N__21228),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__3595 (
            .O(N__21223),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__3594 (
            .O(N__21218),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__3593 (
            .O(N__21213),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__3592 (
            .O(N__21204),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__3591 (
            .O(N__21199),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    InMux I__3590 (
            .O(N__21184),
            .I(N__21178));
    InMux I__3589 (
            .O(N__21183),
            .I(N__21178));
    LocalMux I__3588 (
            .O(N__21178),
            .I(N__21175));
    Span4Mux_h I__3587 (
            .O(N__21175),
            .I(N__21172));
    Odrv4 I__3586 (
            .O(N__21172),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI765BZ0Z1 ));
    InMux I__3585 (
            .O(N__21169),
            .I(\POWERLED.un1_dutycycle_94_cry_2 ));
    InMux I__3584 (
            .O(N__21166),
            .I(N__21163));
    LocalMux I__3583 (
            .O(N__21163),
            .I(N__21159));
    InMux I__3582 (
            .O(N__21162),
            .I(N__21156));
    Sp12to4 I__3581 (
            .O(N__21159),
            .I(N__21151));
    LocalMux I__3580 (
            .O(N__21156),
            .I(N__21151));
    Odrv12 I__3579 (
            .O(N__21151),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI886BZ0Z1 ));
    InMux I__3578 (
            .O(N__21148),
            .I(\POWERLED.un1_dutycycle_94_cry_3 ));
    InMux I__3577 (
            .O(N__21145),
            .I(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ));
    InMux I__3576 (
            .O(N__21142),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__3575 (
            .O(N__21139),
            .I(N__21132));
    InMux I__3574 (
            .O(N__21138),
            .I(N__21132));
    CascadeMux I__3573 (
            .O(N__21137),
            .I(N__21126));
    LocalMux I__3572 (
            .O(N__21132),
            .I(N__21118));
    InMux I__3571 (
            .O(N__21131),
            .I(N__21115));
    InMux I__3570 (
            .O(N__21130),
            .I(N__21110));
    InMux I__3569 (
            .O(N__21129),
            .I(N__21110));
    InMux I__3568 (
            .O(N__21126),
            .I(N__21095));
    InMux I__3567 (
            .O(N__21125),
            .I(N__21095));
    InMux I__3566 (
            .O(N__21124),
            .I(N__21095));
    CascadeMux I__3565 (
            .O(N__21123),
            .I(N__21092));
    CascadeMux I__3564 (
            .O(N__21122),
            .I(N__21089));
    CascadeMux I__3563 (
            .O(N__21121),
            .I(N__21086));
    Span4Mux_h I__3562 (
            .O(N__21118),
            .I(N__21083));
    LocalMux I__3561 (
            .O(N__21115),
            .I(N__21078));
    LocalMux I__3560 (
            .O(N__21110),
            .I(N__21078));
    InMux I__3559 (
            .O(N__21109),
            .I(N__21073));
    InMux I__3558 (
            .O(N__21108),
            .I(N__21073));
    InMux I__3557 (
            .O(N__21107),
            .I(N__21068));
    InMux I__3556 (
            .O(N__21106),
            .I(N__21068));
    InMux I__3555 (
            .O(N__21105),
            .I(N__21054));
    InMux I__3554 (
            .O(N__21104),
            .I(N__21054));
    InMux I__3553 (
            .O(N__21103),
            .I(N__21054));
    InMux I__3552 (
            .O(N__21102),
            .I(N__21051));
    LocalMux I__3551 (
            .O(N__21095),
            .I(N__21048));
    InMux I__3550 (
            .O(N__21092),
            .I(N__21045));
    InMux I__3549 (
            .O(N__21089),
            .I(N__21040));
    InMux I__3548 (
            .O(N__21086),
            .I(N__21040));
    Span4Mux_v I__3547 (
            .O(N__21083),
            .I(N__21035));
    Span4Mux_h I__3546 (
            .O(N__21078),
            .I(N__21035));
    LocalMux I__3545 (
            .O(N__21073),
            .I(N__21030));
    LocalMux I__3544 (
            .O(N__21068),
            .I(N__21030));
    InMux I__3543 (
            .O(N__21067),
            .I(N__21023));
    InMux I__3542 (
            .O(N__21066),
            .I(N__21023));
    InMux I__3541 (
            .O(N__21065),
            .I(N__21023));
    InMux I__3540 (
            .O(N__21064),
            .I(N__21016));
    InMux I__3539 (
            .O(N__21063),
            .I(N__21016));
    InMux I__3538 (
            .O(N__21062),
            .I(N__21016));
    InMux I__3537 (
            .O(N__21061),
            .I(N__21013));
    LocalMux I__3536 (
            .O(N__21054),
            .I(N__21010));
    LocalMux I__3535 (
            .O(N__21051),
            .I(N__21003));
    Span4Mux_s3_h I__3534 (
            .O(N__21048),
            .I(N__21003));
    LocalMux I__3533 (
            .O(N__21045),
            .I(N__21003));
    LocalMux I__3532 (
            .O(N__21040),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__3531 (
            .O(N__21035),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__3530 (
            .O(N__21030),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__3529 (
            .O(N__21023),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__3528 (
            .O(N__21016),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__3527 (
            .O(N__21013),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__3526 (
            .O(N__21010),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__3525 (
            .O(N__21003),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    InMux I__3524 (
            .O(N__20986),
            .I(N__20980));
    InMux I__3523 (
            .O(N__20985),
            .I(N__20980));
    LocalMux I__3522 (
            .O(N__20980),
            .I(N__20977));
    Odrv4 I__3521 (
            .O(N__20977),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4AZ0Z1 ));
    InMux I__3520 (
            .O(N__20974),
            .I(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ));
    CascadeMux I__3519 (
            .O(N__20971),
            .I(N__20965));
    InMux I__3518 (
            .O(N__20970),
            .I(N__20959));
    InMux I__3517 (
            .O(N__20969),
            .I(N__20952));
    InMux I__3516 (
            .O(N__20968),
            .I(N__20952));
    InMux I__3515 (
            .O(N__20965),
            .I(N__20952));
    InMux I__3514 (
            .O(N__20964),
            .I(N__20944));
    InMux I__3513 (
            .O(N__20963),
            .I(N__20944));
    CascadeMux I__3512 (
            .O(N__20962),
            .I(N__20934));
    LocalMux I__3511 (
            .O(N__20959),
            .I(N__20928));
    LocalMux I__3510 (
            .O(N__20952),
            .I(N__20925));
    CascadeMux I__3509 (
            .O(N__20951),
            .I(N__20921));
    InMux I__3508 (
            .O(N__20950),
            .I(N__20914));
    InMux I__3507 (
            .O(N__20949),
            .I(N__20914));
    LocalMux I__3506 (
            .O(N__20944),
            .I(N__20910));
    InMux I__3505 (
            .O(N__20943),
            .I(N__20907));
    InMux I__3504 (
            .O(N__20942),
            .I(N__20898));
    InMux I__3503 (
            .O(N__20941),
            .I(N__20898));
    InMux I__3502 (
            .O(N__20940),
            .I(N__20898));
    InMux I__3501 (
            .O(N__20939),
            .I(N__20898));
    InMux I__3500 (
            .O(N__20938),
            .I(N__20895));
    InMux I__3499 (
            .O(N__20937),
            .I(N__20892));
    InMux I__3498 (
            .O(N__20934),
            .I(N__20889));
    InMux I__3497 (
            .O(N__20933),
            .I(N__20882));
    InMux I__3496 (
            .O(N__20932),
            .I(N__20882));
    InMux I__3495 (
            .O(N__20931),
            .I(N__20882));
    Span4Mux_h I__3494 (
            .O(N__20928),
            .I(N__20877));
    Span4Mux_s3_h I__3493 (
            .O(N__20925),
            .I(N__20877));
    InMux I__3492 (
            .O(N__20924),
            .I(N__20868));
    InMux I__3491 (
            .O(N__20921),
            .I(N__20868));
    InMux I__3490 (
            .O(N__20920),
            .I(N__20868));
    InMux I__3489 (
            .O(N__20919),
            .I(N__20868));
    LocalMux I__3488 (
            .O(N__20914),
            .I(N__20865));
    InMux I__3487 (
            .O(N__20913),
            .I(N__20862));
    Span4Mux_h I__3486 (
            .O(N__20910),
            .I(N__20859));
    LocalMux I__3485 (
            .O(N__20907),
            .I(N__20854));
    LocalMux I__3484 (
            .O(N__20898),
            .I(N__20854));
    LocalMux I__3483 (
            .O(N__20895),
            .I(N__20847));
    LocalMux I__3482 (
            .O(N__20892),
            .I(N__20847));
    LocalMux I__3481 (
            .O(N__20889),
            .I(N__20847));
    LocalMux I__3480 (
            .O(N__20882),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__3479 (
            .O(N__20877),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3478 (
            .O(N__20868),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__3477 (
            .O(N__20865),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3476 (
            .O(N__20862),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__3475 (
            .O(N__20859),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv12 I__3474 (
            .O(N__20854),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv12 I__3473 (
            .O(N__20847),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    InMux I__3472 (
            .O(N__20830),
            .I(N__20824));
    InMux I__3471 (
            .O(N__20829),
            .I(N__20824));
    LocalMux I__3470 (
            .O(N__20824),
            .I(N__20821));
    Odrv12 I__3469 (
            .O(N__20821),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNICGABZ0Z1 ));
    InMux I__3468 (
            .O(N__20818),
            .I(bfn_7_8_0_));
    InMux I__3467 (
            .O(N__20815),
            .I(N__20802));
    CascadeMux I__3466 (
            .O(N__20814),
            .I(N__20799));
    InMux I__3465 (
            .O(N__20813),
            .I(N__20794));
    InMux I__3464 (
            .O(N__20812),
            .I(N__20794));
    InMux I__3463 (
            .O(N__20811),
            .I(N__20785));
    InMux I__3462 (
            .O(N__20810),
            .I(N__20785));
    InMux I__3461 (
            .O(N__20809),
            .I(N__20785));
    InMux I__3460 (
            .O(N__20808),
            .I(N__20785));
    InMux I__3459 (
            .O(N__20807),
            .I(N__20780));
    InMux I__3458 (
            .O(N__20806),
            .I(N__20780));
    InMux I__3457 (
            .O(N__20805),
            .I(N__20777));
    LocalMux I__3456 (
            .O(N__20802),
            .I(N__20768));
    InMux I__3455 (
            .O(N__20799),
            .I(N__20765));
    LocalMux I__3454 (
            .O(N__20794),
            .I(N__20759));
    LocalMux I__3453 (
            .O(N__20785),
            .I(N__20756));
    LocalMux I__3452 (
            .O(N__20780),
            .I(N__20751));
    LocalMux I__3451 (
            .O(N__20777),
            .I(N__20751));
    InMux I__3450 (
            .O(N__20776),
            .I(N__20746));
    InMux I__3449 (
            .O(N__20775),
            .I(N__20746));
    CascadeMux I__3448 (
            .O(N__20774),
            .I(N__20743));
    InMux I__3447 (
            .O(N__20773),
            .I(N__20740));
    InMux I__3446 (
            .O(N__20772),
            .I(N__20735));
    InMux I__3445 (
            .O(N__20771),
            .I(N__20735));
    Span4Mux_h I__3444 (
            .O(N__20768),
            .I(N__20732));
    LocalMux I__3443 (
            .O(N__20765),
            .I(N__20729));
    InMux I__3442 (
            .O(N__20764),
            .I(N__20722));
    InMux I__3441 (
            .O(N__20763),
            .I(N__20722));
    InMux I__3440 (
            .O(N__20762),
            .I(N__20722));
    Span4Mux_v I__3439 (
            .O(N__20759),
            .I(N__20713));
    Span4Mux_s3_h I__3438 (
            .O(N__20756),
            .I(N__20713));
    Span4Mux_v I__3437 (
            .O(N__20751),
            .I(N__20713));
    LocalMux I__3436 (
            .O(N__20746),
            .I(N__20713));
    InMux I__3435 (
            .O(N__20743),
            .I(N__20710));
    LocalMux I__3434 (
            .O(N__20740),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__3433 (
            .O(N__20735),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__3432 (
            .O(N__20732),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__3431 (
            .O(N__20729),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__3430 (
            .O(N__20722),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__3429 (
            .O(N__20713),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__3428 (
            .O(N__20710),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    InMux I__3427 (
            .O(N__20695),
            .I(N__20689));
    InMux I__3426 (
            .O(N__20694),
            .I(N__20689));
    LocalMux I__3425 (
            .O(N__20689),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ));
    InMux I__3424 (
            .O(N__20686),
            .I(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ));
    InMux I__3423 (
            .O(N__20683),
            .I(N__20677));
    InMux I__3422 (
            .O(N__20682),
            .I(N__20677));
    LocalMux I__3421 (
            .O(N__20677),
            .I(N__20674));
    Span4Mux_v I__3420 (
            .O(N__20674),
            .I(N__20671));
    Odrv4 I__3419 (
            .O(N__20671),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCBZ0Z1 ));
    InMux I__3418 (
            .O(N__20668),
            .I(\POWERLED.un1_dutycycle_94_cry_9 ));
    InMux I__3417 (
            .O(N__20665),
            .I(N__20659));
    InMux I__3416 (
            .O(N__20664),
            .I(N__20659));
    LocalMux I__3415 (
            .O(N__20659),
            .I(N__20656));
    Odrv4 I__3414 (
            .O(N__20656),
            .I(\POWERLED.dutycycle_0_6 ));
    CascadeMux I__3413 (
            .O(N__20653),
            .I(\POWERLED.dutycycleZ1Z_6_cascade_ ));
    CascadeMux I__3412 (
            .O(N__20650),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_0_cascade_ ));
    CascadeMux I__3411 (
            .O(N__20647),
            .I(N__20644));
    InMux I__3410 (
            .O(N__20644),
            .I(N__20641));
    LocalMux I__3409 (
            .O(N__20641),
            .I(\POWERLED.un1_dutycycle_96_0_a3_0 ));
    CascadeMux I__3408 (
            .O(N__20638),
            .I(N__20635));
    InMux I__3407 (
            .O(N__20635),
            .I(N__20632));
    LocalMux I__3406 (
            .O(N__20632),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_0 ));
    CascadeMux I__3405 (
            .O(N__20629),
            .I(\POWERLED.un2_count_clk_17_0_cascade_ ));
    InMux I__3404 (
            .O(N__20626),
            .I(N__20623));
    LocalMux I__3403 (
            .O(N__20623),
            .I(N__20620));
    Odrv4 I__3402 (
            .O(N__20620),
            .I(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ));
    InMux I__3401 (
            .O(N__20617),
            .I(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__3400 (
            .O(N__20614),
            .I(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ));
    CascadeMux I__3399 (
            .O(N__20611),
            .I(\POWERLED.func_state_RNISKPU6Z0Z_0_cascade_ ));
    InMux I__3398 (
            .O(N__20608),
            .I(N__20602));
    InMux I__3397 (
            .O(N__20607),
            .I(N__20602));
    LocalMux I__3396 (
            .O(N__20602),
            .I(\POWERLED.count_off_1_13 ));
    InMux I__3395 (
            .O(N__20599),
            .I(N__20596));
    LocalMux I__3394 (
            .O(N__20596),
            .I(\POWERLED.count_off_0_13 ));
    InMux I__3393 (
            .O(N__20593),
            .I(N__20587));
    InMux I__3392 (
            .O(N__20592),
            .I(N__20587));
    LocalMux I__3391 (
            .O(N__20587),
            .I(\POWERLED.count_off_1_14 ));
    InMux I__3390 (
            .O(N__20584),
            .I(N__20581));
    LocalMux I__3389 (
            .O(N__20581),
            .I(\POWERLED.count_off_0_14 ));
    InMux I__3388 (
            .O(N__20578),
            .I(N__20574));
    InMux I__3387 (
            .O(N__20577),
            .I(N__20571));
    LocalMux I__3386 (
            .O(N__20574),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2 ));
    LocalMux I__3385 (
            .O(N__20571),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2 ));
    InMux I__3384 (
            .O(N__20566),
            .I(N__20563));
    LocalMux I__3383 (
            .O(N__20563),
            .I(\POWERLED.count_off_0_15 ));
    InMux I__3382 (
            .O(N__20560),
            .I(N__20557));
    LocalMux I__3381 (
            .O(N__20557),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__3380 (
            .O(N__20554),
            .I(N__20550));
    InMux I__3379 (
            .O(N__20553),
            .I(N__20547));
    LocalMux I__3378 (
            .O(N__20550),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__3377 (
            .O(N__20547),
            .I(\POWERLED.count_offZ0Z_13 ));
    CascadeMux I__3376 (
            .O(N__20542),
            .I(\POWERLED.count_offZ0Z_15_cascade_ ));
    InMux I__3375 (
            .O(N__20539),
            .I(N__20535));
    InMux I__3374 (
            .O(N__20538),
            .I(N__20532));
    LocalMux I__3373 (
            .O(N__20535),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__3372 (
            .O(N__20532),
            .I(\POWERLED.count_offZ0Z_14 ));
    CascadeMux I__3371 (
            .O(N__20527),
            .I(\POWERLED.dutycycleZ0Z_1_cascade_ ));
    InMux I__3370 (
            .O(N__20524),
            .I(N__20521));
    LocalMux I__3369 (
            .O(N__20521),
            .I(\POWERLED.dutycycle_eena ));
    CascadeMux I__3368 (
            .O(N__20518),
            .I(\POWERLED.dutycycle_eena_cascade_ ));
    CascadeMux I__3367 (
            .O(N__20515),
            .I(N__20511));
    InMux I__3366 (
            .O(N__20514),
            .I(N__20508));
    InMux I__3365 (
            .O(N__20511),
            .I(N__20505));
    LocalMux I__3364 (
            .O(N__20508),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    LocalMux I__3363 (
            .O(N__20505),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    CascadeMux I__3362 (
            .O(N__20500),
            .I(\POWERLED.dutycycle_1_0_1_cascade_ ));
    InMux I__3361 (
            .O(N__20497),
            .I(N__20494));
    LocalMux I__3360 (
            .O(N__20494),
            .I(\POWERLED.dutycycle_eena_0 ));
    InMux I__3359 (
            .O(N__20491),
            .I(N__20488));
    LocalMux I__3358 (
            .O(N__20488),
            .I(\POWERLED.dutycycle_1_0_1 ));
    InMux I__3357 (
            .O(N__20485),
            .I(N__20479));
    InMux I__3356 (
            .O(N__20484),
            .I(N__20479));
    LocalMux I__3355 (
            .O(N__20479),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    CascadeMux I__3354 (
            .O(N__20476),
            .I(\POWERLED.dutycycle_eena_0_cascade_ ));
    InMux I__3353 (
            .O(N__20473),
            .I(N__20467));
    InMux I__3352 (
            .O(N__20472),
            .I(N__20467));
    LocalMux I__3351 (
            .O(N__20467),
            .I(\POWERLED.dutycycle_1_0_0 ));
    CascadeMux I__3350 (
            .O(N__20464),
            .I(N__20461));
    InMux I__3349 (
            .O(N__20461),
            .I(N__20458));
    LocalMux I__3348 (
            .O(N__20458),
            .I(\PCH_PWRGD.count_0_14 ));
    InMux I__3347 (
            .O(N__20455),
            .I(N__20449));
    InMux I__3346 (
            .O(N__20454),
            .I(N__20449));
    LocalMux I__3345 (
            .O(N__20449),
            .I(\PCH_PWRGD.count_0_2 ));
    CascadeMux I__3344 (
            .O(N__20446),
            .I(\PCH_PWRGD.countZ0Z_14_cascade_ ));
    InMux I__3343 (
            .O(N__20443),
            .I(N__20440));
    LocalMux I__3342 (
            .O(N__20440),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__3341 (
            .O(N__20437),
            .I(N__20431));
    InMux I__3340 (
            .O(N__20436),
            .I(N__20431));
    LocalMux I__3339 (
            .O(N__20431),
            .I(N__20427));
    InMux I__3338 (
            .O(N__20430),
            .I(N__20424));
    Span4Mux_s3_h I__3337 (
            .O(N__20427),
            .I(N__20419));
    LocalMux I__3336 (
            .O(N__20424),
            .I(N__20419));
    Odrv4 I__3335 (
            .O(N__20419),
            .I(PCH_PWRGD_delayed_vccin_ok));
    InMux I__3334 (
            .O(N__20416),
            .I(N__20413));
    LocalMux I__3333 (
            .O(N__20413),
            .I(\PCH_PWRGD.N_250_0 ));
    CascadeMux I__3332 (
            .O(N__20410),
            .I(\PCH_PWRGD.N_250_0_cascade_ ));
    InMux I__3331 (
            .O(N__20407),
            .I(N__20401));
    InMux I__3330 (
            .O(N__20406),
            .I(N__20401));
    LocalMux I__3329 (
            .O(N__20401),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    InMux I__3328 (
            .O(N__20398),
            .I(N__20395));
    LocalMux I__3327 (
            .O(N__20395),
            .I(\PCH_PWRGD.count_0_15 ));
    InMux I__3326 (
            .O(N__20392),
            .I(N__20386));
    InMux I__3325 (
            .O(N__20391),
            .I(N__20386));
    LocalMux I__3324 (
            .O(N__20386),
            .I(\PCH_PWRGD.count_0_13 ));
    CascadeMux I__3323 (
            .O(N__20383),
            .I(\PCH_PWRGD.countZ0Z_15_cascade_ ));
    CascadeMux I__3322 (
            .O(N__20380),
            .I(\PCH_PWRGD.count_rst_10_cascade_ ));
    CascadeMux I__3321 (
            .O(N__20377),
            .I(\PCH_PWRGD.un2_count_1_axb_4_cascade_ ));
    InMux I__3320 (
            .O(N__20374),
            .I(N__20371));
    LocalMux I__3319 (
            .O(N__20371),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__3318 (
            .O(N__20368),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    CascadeMux I__3317 (
            .O(N__20365),
            .I(N__20362));
    InMux I__3316 (
            .O(N__20362),
            .I(N__20359));
    LocalMux I__3315 (
            .O(N__20359),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__3314 (
            .O(N__20356),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    CascadeMux I__3313 (
            .O(N__20353),
            .I(N__20350));
    InMux I__3312 (
            .O(N__20350),
            .I(N__20347));
    LocalMux I__3311 (
            .O(N__20347),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__3310 (
            .O(N__20344),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    InMux I__3309 (
            .O(N__20341),
            .I(N__20338));
    LocalMux I__3308 (
            .O(N__20338),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__3307 (
            .O(N__20335),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__3306 (
            .O(N__20332),
            .I(\POWERLED.mult1_un145_sum_s_8_cascade_ ));
    CascadeMux I__3305 (
            .O(N__20329),
            .I(N__20325));
    InMux I__3304 (
            .O(N__20328),
            .I(N__20318));
    InMux I__3303 (
            .O(N__20325),
            .I(N__20318));
    InMux I__3302 (
            .O(N__20324),
            .I(N__20315));
    InMux I__3301 (
            .O(N__20323),
            .I(N__20312));
    LocalMux I__3300 (
            .O(N__20318),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__3299 (
            .O(N__20315),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__3298 (
            .O(N__20312),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__3297 (
            .O(N__20305),
            .I(N__20301));
    InMux I__3296 (
            .O(N__20304),
            .I(N__20293));
    InMux I__3295 (
            .O(N__20301),
            .I(N__20293));
    InMux I__3294 (
            .O(N__20300),
            .I(N__20293));
    LocalMux I__3293 (
            .O(N__20293),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    InMux I__3292 (
            .O(N__20290),
            .I(N__20287));
    LocalMux I__3291 (
            .O(N__20287),
            .I(N__20284));
    Span4Mux_s3_v I__3290 (
            .O(N__20284),
            .I(N__20280));
    InMux I__3289 (
            .O(N__20283),
            .I(N__20277));
    Span4Mux_v I__3288 (
            .O(N__20280),
            .I(N__20274));
    LocalMux I__3287 (
            .O(N__20277),
            .I(N__20271));
    Odrv4 I__3286 (
            .O(N__20274),
            .I(\POWERLED.mult1_un131_sum ));
    Odrv12 I__3285 (
            .O(N__20271),
            .I(\POWERLED.mult1_un131_sum ));
    CascadeMux I__3284 (
            .O(N__20266),
            .I(N__20263));
    InMux I__3283 (
            .O(N__20263),
            .I(N__20260));
    LocalMux I__3282 (
            .O(N__20260),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__3281 (
            .O(N__20257),
            .I(N__20254));
    LocalMux I__3280 (
            .O(N__20254),
            .I(N__20251));
    Span4Mux_h I__3279 (
            .O(N__20251),
            .I(N__20247));
    InMux I__3278 (
            .O(N__20250),
            .I(N__20244));
    Sp12to4 I__3277 (
            .O(N__20247),
            .I(N__20239));
    LocalMux I__3276 (
            .O(N__20244),
            .I(N__20239));
    Odrv12 I__3275 (
            .O(N__20239),
            .I(\POWERLED.mult1_un89_sum ));
    CascadeMux I__3274 (
            .O(N__20236),
            .I(N__20233));
    InMux I__3273 (
            .O(N__20233),
            .I(N__20230));
    LocalMux I__3272 (
            .O(N__20230),
            .I(N__20227));
    Span4Mux_h I__3271 (
            .O(N__20227),
            .I(N__20224));
    Odrv4 I__3270 (
            .O(N__20224),
            .I(\POWERLED.mult1_un89_sum_i ));
    CascadeMux I__3269 (
            .O(N__20221),
            .I(N__20217));
    CascadeMux I__3268 (
            .O(N__20220),
            .I(N__20214));
    InMux I__3267 (
            .O(N__20217),
            .I(N__20208));
    InMux I__3266 (
            .O(N__20214),
            .I(N__20203));
    InMux I__3265 (
            .O(N__20213),
            .I(N__20203));
    InMux I__3264 (
            .O(N__20212),
            .I(N__20200));
    InMux I__3263 (
            .O(N__20211),
            .I(N__20197));
    LocalMux I__3262 (
            .O(N__20208),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3261 (
            .O(N__20203),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3260 (
            .O(N__20200),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__3259 (
            .O(N__20197),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__3258 (
            .O(N__20188),
            .I(N__20185));
    InMux I__3257 (
            .O(N__20185),
            .I(N__20182));
    LocalMux I__3256 (
            .O(N__20182),
            .I(N__20179));
    Span4Mux_s1_h I__3255 (
            .O(N__20179),
            .I(N__20176));
    Span4Mux_h I__3254 (
            .O(N__20176),
            .I(N__20173));
    Odrv4 I__3253 (
            .O(N__20173),
            .I(\POWERLED.mult1_un68_sum_i_8 ));
    CascadeMux I__3252 (
            .O(N__20170),
            .I(N__20167));
    InMux I__3251 (
            .O(N__20167),
            .I(N__20163));
    InMux I__3250 (
            .O(N__20166),
            .I(N__20160));
    LocalMux I__3249 (
            .O(N__20163),
            .I(N__20155));
    LocalMux I__3248 (
            .O(N__20160),
            .I(N__20155));
    Odrv4 I__3247 (
            .O(N__20155),
            .I(\POWERLED.mult1_un75_sum ));
    CascadeMux I__3246 (
            .O(N__20152),
            .I(N__20149));
    InMux I__3245 (
            .O(N__20149),
            .I(N__20146));
    LocalMux I__3244 (
            .O(N__20146),
            .I(\POWERLED.mult1_un75_sum_i ));
    InMux I__3243 (
            .O(N__20143),
            .I(N__20140));
    LocalMux I__3242 (
            .O(N__20140),
            .I(N__20136));
    InMux I__3241 (
            .O(N__20139),
            .I(N__20133));
    Sp12to4 I__3240 (
            .O(N__20136),
            .I(N__20128));
    LocalMux I__3239 (
            .O(N__20133),
            .I(N__20128));
    Odrv12 I__3238 (
            .O(N__20128),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__3237 (
            .O(N__20125),
            .I(N__20122));
    LocalMux I__3236 (
            .O(N__20122),
            .I(N__20119));
    Odrv12 I__3235 (
            .O(N__20119),
            .I(\POWERLED.un85_clk_100khz_2 ));
    InMux I__3234 (
            .O(N__20116),
            .I(N__20112));
    InMux I__3233 (
            .O(N__20115),
            .I(N__20109));
    LocalMux I__3232 (
            .O(N__20112),
            .I(N__20106));
    LocalMux I__3231 (
            .O(N__20109),
            .I(N__20103));
    Span12Mux_s5_h I__3230 (
            .O(N__20106),
            .I(N__20100));
    Span4Mux_v I__3229 (
            .O(N__20103),
            .I(N__20097));
    Odrv12 I__3228 (
            .O(N__20100),
            .I(\POWERLED.mult1_un96_sum ));
    Odrv4 I__3227 (
            .O(N__20097),
            .I(\POWERLED.mult1_un96_sum ));
    CascadeMux I__3226 (
            .O(N__20092),
            .I(N__20089));
    InMux I__3225 (
            .O(N__20089),
            .I(N__20086));
    LocalMux I__3224 (
            .O(N__20086),
            .I(N__20083));
    Span4Mux_s3_v I__3223 (
            .O(N__20083),
            .I(N__20080));
    Odrv4 I__3222 (
            .O(N__20080),
            .I(\POWERLED.mult1_un96_sum_i ));
    InMux I__3221 (
            .O(N__20077),
            .I(N__20074));
    LocalMux I__3220 (
            .O(N__20074),
            .I(N__20070));
    InMux I__3219 (
            .O(N__20073),
            .I(N__20067));
    Span4Mux_v I__3218 (
            .O(N__20070),
            .I(N__20062));
    LocalMux I__3217 (
            .O(N__20067),
            .I(N__20062));
    Span4Mux_v I__3216 (
            .O(N__20062),
            .I(N__20059));
    Odrv4 I__3215 (
            .O(N__20059),
            .I(\POWERLED.mult1_un145_sum ));
    CascadeMux I__3214 (
            .O(N__20056),
            .I(N__20053));
    InMux I__3213 (
            .O(N__20053),
            .I(N__20050));
    LocalMux I__3212 (
            .O(N__20050),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__3211 (
            .O(N__20047),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    InMux I__3210 (
            .O(N__20044),
            .I(N__20041));
    LocalMux I__3209 (
            .O(N__20041),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__3208 (
            .O(N__20038),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    CascadeMux I__3207 (
            .O(N__20035),
            .I(N__20032));
    InMux I__3206 (
            .O(N__20032),
            .I(N__20029));
    LocalMux I__3205 (
            .O(N__20029),
            .I(N__20026));
    Span4Mux_v I__3204 (
            .O(N__20026),
            .I(N__20023));
    Span4Mux_h I__3203 (
            .O(N__20023),
            .I(N__20020));
    Odrv4 I__3202 (
            .O(N__20020),
            .I(\POWERLED.g2_1 ));
    InMux I__3201 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__3200 (
            .O(N__20014),
            .I(N__20011));
    Odrv4 I__3199 (
            .O(N__20011),
            .I(\POWERLED.g2_5 ));
    InMux I__3198 (
            .O(N__20008),
            .I(N__20005));
    LocalMux I__3197 (
            .O(N__20005),
            .I(N__20002));
    Span4Mux_h I__3196 (
            .O(N__20002),
            .I(N__19999));
    Span4Mux_v I__3195 (
            .O(N__19999),
            .I(N__19996));
    Odrv4 I__3194 (
            .O(N__19996),
            .I(\POWERLED.g0_4_4 ));
    CascadeMux I__3193 (
            .O(N__19993),
            .I(\POWERLED.g0_4_5_cascade_ ));
    CascadeMux I__3192 (
            .O(N__19990),
            .I(N__19986));
    InMux I__3191 (
            .O(N__19989),
            .I(N__19983));
    InMux I__3190 (
            .O(N__19986),
            .I(N__19980));
    LocalMux I__3189 (
            .O(N__19983),
            .I(N__19975));
    LocalMux I__3188 (
            .O(N__19980),
            .I(N__19975));
    Odrv4 I__3187 (
            .O(N__19975),
            .I(\POWERLED.mult1_un68_sum ));
    CascadeMux I__3186 (
            .O(N__19972),
            .I(N__19969));
    InMux I__3185 (
            .O(N__19969),
            .I(N__19966));
    LocalMux I__3184 (
            .O(N__19966),
            .I(N__19963));
    Odrv4 I__3183 (
            .O(N__19963),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__3182 (
            .O(N__19960),
            .I(N__19957));
    LocalMux I__3181 (
            .O(N__19957),
            .I(\POWERLED.g3_1_0 ));
    CascadeMux I__3180 (
            .O(N__19954),
            .I(\POWERLED.g3_1_4_cascade_ ));
    CascadeMux I__3179 (
            .O(N__19951),
            .I(\POWERLED.g3_1_6_cascade_ ));
    CascadeMux I__3178 (
            .O(N__19948),
            .I(N__19945));
    InMux I__3177 (
            .O(N__19945),
            .I(N__19938));
    InMux I__3176 (
            .O(N__19944),
            .I(N__19938));
    CascadeMux I__3175 (
            .O(N__19943),
            .I(N__19935));
    LocalMux I__3174 (
            .O(N__19938),
            .I(N__19932));
    InMux I__3173 (
            .O(N__19935),
            .I(N__19929));
    Span4Mux_h I__3172 (
            .O(N__19932),
            .I(N__19924));
    LocalMux I__3171 (
            .O(N__19929),
            .I(N__19924));
    Odrv4 I__3170 (
            .O(N__19924),
            .I(\POWERLED.un2_count_clk_17_0_a2_5 ));
    CascadeMux I__3169 (
            .O(N__19921),
            .I(N__19918));
    InMux I__3168 (
            .O(N__19918),
            .I(N__19915));
    LocalMux I__3167 (
            .O(N__19915),
            .I(N__19912));
    Odrv4 I__3166 (
            .O(N__19912),
            .I(\POWERLED.dutycycle_RNIZ0Z_15 ));
    InMux I__3165 (
            .O(N__19909),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    CascadeMux I__3164 (
            .O(N__19906),
            .I(N__19903));
    InMux I__3163 (
            .O(N__19903),
            .I(N__19900));
    LocalMux I__3162 (
            .O(N__19900),
            .I(N__19897));
    Span4Mux_h I__3161 (
            .O(N__19897),
            .I(N__19894));
    Odrv4 I__3160 (
            .O(N__19894),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_13 ));
    InMux I__3159 (
            .O(N__19891),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__3158 (
            .O(N__19888),
            .I(N__19885));
    LocalMux I__3157 (
            .O(N__19885),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    InMux I__3156 (
            .O(N__19882),
            .I(N__19879));
    LocalMux I__3155 (
            .O(N__19879),
            .I(N__19875));
    CascadeMux I__3154 (
            .O(N__19878),
            .I(N__19872));
    Span4Mux_h I__3153 (
            .O(N__19875),
            .I(N__19869));
    InMux I__3152 (
            .O(N__19872),
            .I(N__19866));
    Odrv4 I__3151 (
            .O(N__19869),
            .I(\POWERLED.mult1_un47_sum ));
    LocalMux I__3150 (
            .O(N__19866),
            .I(\POWERLED.mult1_un47_sum ));
    InMux I__3149 (
            .O(N__19861),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    CascadeMux I__3148 (
            .O(N__19858),
            .I(N__19853));
    InMux I__3147 (
            .O(N__19857),
            .I(N__19843));
    InMux I__3146 (
            .O(N__19856),
            .I(N__19843));
    InMux I__3145 (
            .O(N__19853),
            .I(N__19843));
    InMux I__3144 (
            .O(N__19852),
            .I(N__19843));
    LocalMux I__3143 (
            .O(N__19843),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    InMux I__3142 (
            .O(N__19840),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    CascadeMux I__3141 (
            .O(N__19837),
            .I(N__19833));
    InMux I__3140 (
            .O(N__19836),
            .I(N__19825));
    InMux I__3139 (
            .O(N__19833),
            .I(N__19825));
    InMux I__3138 (
            .O(N__19832),
            .I(N__19825));
    LocalMux I__3137 (
            .O(N__19825),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    InMux I__3136 (
            .O(N__19822),
            .I(bfn_6_11_0_));
    InMux I__3135 (
            .O(N__19819),
            .I(\POWERLED.CO2 ));
    CascadeMux I__3134 (
            .O(N__19816),
            .I(N__19813));
    InMux I__3133 (
            .O(N__19813),
            .I(N__19807));
    InMux I__3132 (
            .O(N__19812),
            .I(N__19807));
    LocalMux I__3131 (
            .O(N__19807),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__3130 (
            .O(N__19804),
            .I(N__19801));
    InMux I__3129 (
            .O(N__19801),
            .I(N__19798));
    LocalMux I__3128 (
            .O(N__19798),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    InMux I__3127 (
            .O(N__19795),
            .I(N__19791));
    InMux I__3126 (
            .O(N__19794),
            .I(N__19788));
    LocalMux I__3125 (
            .O(N__19791),
            .I(\POWERLED.mult1_un61_sum ));
    LocalMux I__3124 (
            .O(N__19788),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__3123 (
            .O(N__19783),
            .I(N__19780));
    LocalMux I__3122 (
            .O(N__19780),
            .I(N__19777));
    Span4Mux_h I__3121 (
            .O(N__19777),
            .I(N__19774));
    Odrv4 I__3120 (
            .O(N__19774),
            .I(\POWERLED.mult1_un61_sum_i ));
    CascadeMux I__3119 (
            .O(N__19771),
            .I(N__19768));
    InMux I__3118 (
            .O(N__19768),
            .I(N__19764));
    InMux I__3117 (
            .O(N__19767),
            .I(N__19761));
    LocalMux I__3116 (
            .O(N__19764),
            .I(N__19758));
    LocalMux I__3115 (
            .O(N__19761),
            .I(\POWERLED.mult1_un54_sum ));
    Odrv4 I__3114 (
            .O(N__19758),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__3113 (
            .O(N__19753),
            .I(N__19750));
    LocalMux I__3112 (
            .O(N__19750),
            .I(N__19747));
    Odrv4 I__3111 (
            .O(N__19747),
            .I(\POWERLED.mult1_un54_sum_i ));
    InMux I__3110 (
            .O(N__19744),
            .I(N__19741));
    LocalMux I__3109 (
            .O(N__19741),
            .I(N__19738));
    Span4Mux_h I__3108 (
            .O(N__19738),
            .I(N__19735));
    Odrv4 I__3107 (
            .O(N__19735),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_3 ));
    InMux I__3106 (
            .O(N__19732),
            .I(N__19729));
    LocalMux I__3105 (
            .O(N__19729),
            .I(N__19725));
    CascadeMux I__3104 (
            .O(N__19728),
            .I(N__19722));
    Sp12to4 I__3103 (
            .O(N__19725),
            .I(N__19719));
    InMux I__3102 (
            .O(N__19722),
            .I(N__19716));
    Odrv12 I__3101 (
            .O(N__19719),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_3 ));
    LocalMux I__3100 (
            .O(N__19716),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_3 ));
    InMux I__3099 (
            .O(N__19711),
            .I(N__19708));
    LocalMux I__3098 (
            .O(N__19708),
            .I(N__19704));
    InMux I__3097 (
            .O(N__19707),
            .I(N__19701));
    Span4Mux_s3_h I__3096 (
            .O(N__19704),
            .I(N__19696));
    LocalMux I__3095 (
            .O(N__19701),
            .I(N__19696));
    Span4Mux_v I__3094 (
            .O(N__19696),
            .I(N__19693));
    Odrv4 I__3093 (
            .O(N__19693),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__3092 (
            .O(N__19690),
            .I(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ));
    CascadeMux I__3091 (
            .O(N__19687),
            .I(N__19684));
    InMux I__3090 (
            .O(N__19684),
            .I(N__19681));
    LocalMux I__3089 (
            .O(N__19681),
            .I(N__19678));
    Span4Mux_v I__3088 (
            .O(N__19678),
            .I(N__19675));
    Odrv4 I__3087 (
            .O(N__19675),
            .I(\POWERLED.dutycycle_RNIZ0Z_4 ));
    InMux I__3086 (
            .O(N__19672),
            .I(N__19668));
    InMux I__3085 (
            .O(N__19671),
            .I(N__19665));
    LocalMux I__3084 (
            .O(N__19668),
            .I(N__19662));
    LocalMux I__3083 (
            .O(N__19665),
            .I(N__19659));
    Span12Mux_s5_h I__3082 (
            .O(N__19662),
            .I(N__19656));
    Span4Mux_v I__3081 (
            .O(N__19659),
            .I(N__19653));
    Odrv12 I__3080 (
            .O(N__19656),
            .I(\POWERLED.mult1_un110_sum ));
    Odrv4 I__3079 (
            .O(N__19653),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__3078 (
            .O(N__19648),
            .I(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ));
    InMux I__3077 (
            .O(N__19645),
            .I(N__19642));
    LocalMux I__3076 (
            .O(N__19642),
            .I(N__19639));
    Span4Mux_h I__3075 (
            .O(N__19639),
            .I(N__19636));
    Odrv4 I__3074 (
            .O(N__19636),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_9 ));
    InMux I__3073 (
            .O(N__19633),
            .I(N__19629));
    InMux I__3072 (
            .O(N__19632),
            .I(N__19626));
    LocalMux I__3071 (
            .O(N__19629),
            .I(N__19623));
    LocalMux I__3070 (
            .O(N__19626),
            .I(N__19620));
    Span12Mux_s5_h I__3069 (
            .O(N__19623),
            .I(N__19617));
    Span4Mux_v I__3068 (
            .O(N__19620),
            .I(N__19614));
    Odrv12 I__3067 (
            .O(N__19617),
            .I(\POWERLED.mult1_un103_sum ));
    Odrv4 I__3066 (
            .O(N__19614),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__3065 (
            .O(N__19609),
            .I(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ));
    CascadeMux I__3064 (
            .O(N__19606),
            .I(N__19603));
    InMux I__3063 (
            .O(N__19603),
            .I(N__19600));
    LocalMux I__3062 (
            .O(N__19600),
            .I(N__19597));
    Span4Mux_v I__3061 (
            .O(N__19597),
            .I(N__19594));
    Odrv4 I__3060 (
            .O(N__19594),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_10 ));
    InMux I__3059 (
            .O(N__19591),
            .I(\POWERLED.un1_dutycycle_53_cry_6 ));
    InMux I__3058 (
            .O(N__19588),
            .I(N__19585));
    LocalMux I__3057 (
            .O(N__19585),
            .I(N__19582));
    Span4Mux_v I__3056 (
            .O(N__19582),
            .I(N__19579));
    Odrv4 I__3055 (
            .O(N__19579),
            .I(\POWERLED.dutycycle_RNIZ0Z_11 ));
    InMux I__3054 (
            .O(N__19576),
            .I(bfn_6_10_0_));
    CascadeMux I__3053 (
            .O(N__19573),
            .I(N__19570));
    InMux I__3052 (
            .O(N__19570),
            .I(N__19567));
    LocalMux I__3051 (
            .O(N__19567),
            .I(N__19564));
    Span4Mux_h I__3050 (
            .O(N__19564),
            .I(N__19561));
    Odrv4 I__3049 (
            .O(N__19561),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_12 ));
    InMux I__3048 (
            .O(N__19558),
            .I(N__19555));
    LocalMux I__3047 (
            .O(N__19555),
            .I(N__19551));
    InMux I__3046 (
            .O(N__19554),
            .I(N__19548));
    Span4Mux_s2_v I__3045 (
            .O(N__19551),
            .I(N__19543));
    LocalMux I__3044 (
            .O(N__19548),
            .I(N__19543));
    Span4Mux_v I__3043 (
            .O(N__19543),
            .I(N__19540));
    Odrv4 I__3042 (
            .O(N__19540),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__3041 (
            .O(N__19537),
            .I(\POWERLED.un1_dutycycle_53_cry_8 ));
    InMux I__3040 (
            .O(N__19534),
            .I(N__19531));
    LocalMux I__3039 (
            .O(N__19531),
            .I(N__19528));
    Span4Mux_v I__3038 (
            .O(N__19528),
            .I(N__19525));
    Odrv4 I__3037 (
            .O(N__19525),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_13 ));
    InMux I__3036 (
            .O(N__19522),
            .I(\POWERLED.un1_dutycycle_53_cry_9 ));
    CascadeMux I__3035 (
            .O(N__19519),
            .I(N__19516));
    InMux I__3034 (
            .O(N__19516),
            .I(N__19513));
    LocalMux I__3033 (
            .O(N__19513),
            .I(N__19510));
    Odrv12 I__3032 (
            .O(N__19510),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_14 ));
    InMux I__3031 (
            .O(N__19507),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    CascadeMux I__3030 (
            .O(N__19504),
            .I(N__19501));
    InMux I__3029 (
            .O(N__19501),
            .I(N__19495));
    InMux I__3028 (
            .O(N__19500),
            .I(N__19495));
    LocalMux I__3027 (
            .O(N__19495),
            .I(N__19492));
    Odrv4 I__3026 (
            .O(N__19492),
            .I(\POWERLED.dutycycle_en_10 ));
    CascadeMux I__3025 (
            .O(N__19489),
            .I(N__19486));
    InMux I__3024 (
            .O(N__19486),
            .I(N__19480));
    InMux I__3023 (
            .O(N__19485),
            .I(N__19480));
    LocalMux I__3022 (
            .O(N__19480),
            .I(\POWERLED.dutycycleZ1Z_13 ));
    InMux I__3021 (
            .O(N__19477),
            .I(N__19471));
    InMux I__3020 (
            .O(N__19476),
            .I(N__19471));
    LocalMux I__3019 (
            .O(N__19471),
            .I(N__19468));
    Span4Mux_h I__3018 (
            .O(N__19468),
            .I(N__19465));
    Odrv4 I__3017 (
            .O(N__19465),
            .I(\POWERLED.un1_dutycycle_53_50_0 ));
    CascadeMux I__3016 (
            .O(N__19462),
            .I(\POWERLED.dutycycle_RNI_12Z0Z_9_cascade_ ));
    InMux I__3015 (
            .O(N__19459),
            .I(N__19456));
    LocalMux I__3014 (
            .O(N__19456),
            .I(\POWERLED.dutycycle_RNI_15Z0Z_9 ));
    InMux I__3013 (
            .O(N__19453),
            .I(N__19448));
    InMux I__3012 (
            .O(N__19452),
            .I(N__19443));
    InMux I__3011 (
            .O(N__19451),
            .I(N__19443));
    LocalMux I__3010 (
            .O(N__19448),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_9 ));
    LocalMux I__3009 (
            .O(N__19443),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_9 ));
    InMux I__3008 (
            .O(N__19438),
            .I(N__19435));
    LocalMux I__3007 (
            .O(N__19435),
            .I(N__19432));
    Span4Mux_h I__3006 (
            .O(N__19432),
            .I(N__19429));
    Span4Mux_h I__3005 (
            .O(N__19429),
            .I(N__19426));
    Odrv4 I__3004 (
            .O(N__19426),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_0 ));
    InMux I__3003 (
            .O(N__19423),
            .I(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ));
    CascadeMux I__3002 (
            .O(N__19420),
            .I(N__19417));
    InMux I__3001 (
            .O(N__19417),
            .I(N__19414));
    LocalMux I__3000 (
            .O(N__19414),
            .I(N__19411));
    Span4Mux_h I__2999 (
            .O(N__19411),
            .I(N__19408));
    Odrv4 I__2998 (
            .O(N__19408),
            .I(\POWERLED.dutycycle_RNIZ0Z_2 ));
    InMux I__2997 (
            .O(N__19405),
            .I(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ));
    InMux I__2996 (
            .O(N__19402),
            .I(N__19399));
    LocalMux I__2995 (
            .O(N__19399),
            .I(N__19396));
    Span4Mux_h I__2994 (
            .O(N__19396),
            .I(N__19393));
    Odrv4 I__2993 (
            .O(N__19393),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_2 ));
    InMux I__2992 (
            .O(N__19390),
            .I(N__19386));
    InMux I__2991 (
            .O(N__19389),
            .I(N__19383));
    LocalMux I__2990 (
            .O(N__19386),
            .I(N__19380));
    LocalMux I__2989 (
            .O(N__19383),
            .I(N__19377));
    Span4Mux_v I__2988 (
            .O(N__19380),
            .I(N__19374));
    Span12Mux_s5_h I__2987 (
            .O(N__19377),
            .I(N__19371));
    Odrv4 I__2986 (
            .O(N__19374),
            .I(\POWERLED.mult1_un124_sum ));
    Odrv12 I__2985 (
            .O(N__19371),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__2984 (
            .O(N__19366),
            .I(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ));
    InMux I__2983 (
            .O(N__19363),
            .I(N__19360));
    LocalMux I__2982 (
            .O(N__19360),
            .I(\POWERLED.un1_clk_100khz_39_and_i_0_0 ));
    CascadeMux I__2981 (
            .O(N__19357),
            .I(\POWERLED.un1_clk_100khz_30_and_i_0_0_cascade_ ));
    InMux I__2980 (
            .O(N__19354),
            .I(N__19351));
    LocalMux I__2979 (
            .O(N__19351),
            .I(\POWERLED.dutycycle_RNI4J2O7Z0Z_9 ));
    CascadeMux I__2978 (
            .O(N__19348),
            .I(N__19345));
    InMux I__2977 (
            .O(N__19345),
            .I(N__19339));
    InMux I__2976 (
            .O(N__19344),
            .I(N__19339));
    LocalMux I__2975 (
            .O(N__19339),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__2974 (
            .O(N__19336),
            .I(\POWERLED.dutycycle_RNI4J2O7Z0Z_9_cascade_ ));
    InMux I__2973 (
            .O(N__19333),
            .I(N__19327));
    InMux I__2972 (
            .O(N__19332),
            .I(N__19327));
    LocalMux I__2971 (
            .O(N__19327),
            .I(\POWERLED.dutycycleZ1Z_11 ));
    CascadeMux I__2970 (
            .O(N__19324),
            .I(N__19321));
    InMux I__2969 (
            .O(N__19321),
            .I(N__19318));
    LocalMux I__2968 (
            .O(N__19318),
            .I(\POWERLED.dutycycle_en_7 ));
    InMux I__2967 (
            .O(N__19315),
            .I(N__19310));
    InMux I__2966 (
            .O(N__19314),
            .I(N__19307));
    InMux I__2965 (
            .O(N__19313),
            .I(N__19304));
    LocalMux I__2964 (
            .O(N__19310),
            .I(N__19301));
    LocalMux I__2963 (
            .O(N__19307),
            .I(N__19298));
    LocalMux I__2962 (
            .O(N__19304),
            .I(N__19294));
    Span4Mux_v I__2961 (
            .O(N__19301),
            .I(N__19289));
    Span4Mux_s3_h I__2960 (
            .O(N__19298),
            .I(N__19289));
    InMux I__2959 (
            .O(N__19297),
            .I(N__19286));
    Span4Mux_h I__2958 (
            .O(N__19294),
            .I(N__19283));
    Odrv4 I__2957 (
            .O(N__19289),
            .I(\POWERLED.un1_dutycycle_53_20_1 ));
    LocalMux I__2956 (
            .O(N__19286),
            .I(\POWERLED.un1_dutycycle_53_20_1 ));
    Odrv4 I__2955 (
            .O(N__19283),
            .I(\POWERLED.un1_dutycycle_53_20_1 ));
    CascadeMux I__2954 (
            .O(N__19276),
            .I(\POWERLED.un1_dutycycle_53_3_2_1_cascade_ ));
    CascadeMux I__2953 (
            .O(N__19273),
            .I(\POWERLED.un1_dutycycle_53_3_2_cascade_ ));
    CascadeMux I__2952 (
            .O(N__19270),
            .I(N__19267));
    InMux I__2951 (
            .O(N__19267),
            .I(N__19261));
    InMux I__2950 (
            .O(N__19266),
            .I(N__19261));
    LocalMux I__2949 (
            .O(N__19261),
            .I(\POWERLED.dutycycleZ1Z_14 ));
    CascadeMux I__2948 (
            .O(N__19258),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    InMux I__2947 (
            .O(N__19255),
            .I(N__19252));
    LocalMux I__2946 (
            .O(N__19252),
            .I(\POWERLED.dutycycle_RNI_13Z0Z_9 ));
    InMux I__2945 (
            .O(N__19249),
            .I(N__19246));
    LocalMux I__2944 (
            .O(N__19246),
            .I(\POWERLED.un1_dutycycle_53_2_0 ));
    CascadeMux I__2943 (
            .O(N__19243),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_11_cascade_ ));
    CascadeMux I__2942 (
            .O(N__19240),
            .I(\POWERLED.un1_dutycycle_53_axb_11_cascade_ ));
    InMux I__2941 (
            .O(N__19237),
            .I(N__19233));
    InMux I__2940 (
            .O(N__19236),
            .I(N__19230));
    LocalMux I__2939 (
            .O(N__19233),
            .I(N__19227));
    LocalMux I__2938 (
            .O(N__19230),
            .I(N__19222));
    Span4Mux_v I__2937 (
            .O(N__19227),
            .I(N__19222));
    Odrv4 I__2936 (
            .O(N__19222),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_4 ));
    CascadeMux I__2935 (
            .O(N__19219),
            .I(\POWERLED.dutycycle_en_7_cascade_ ));
    CascadeMux I__2934 (
            .O(N__19216),
            .I(N__19212));
    InMux I__2933 (
            .O(N__19215),
            .I(N__19209));
    InMux I__2932 (
            .O(N__19212),
            .I(N__19206));
    LocalMux I__2931 (
            .O(N__19209),
            .I(\POWERLED.count_offZ0Z_10 ));
    LocalMux I__2930 (
            .O(N__19206),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__2929 (
            .O(N__19201),
            .I(N__19195));
    InMux I__2928 (
            .O(N__19200),
            .I(N__19195));
    LocalMux I__2927 (
            .O(N__19195),
            .I(\POWERLED.count_off_1_10 ));
    InMux I__2926 (
            .O(N__19192),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    InMux I__2925 (
            .O(N__19189),
            .I(N__19185));
    InMux I__2924 (
            .O(N__19188),
            .I(N__19182));
    LocalMux I__2923 (
            .O(N__19185),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__2922 (
            .O(N__19182),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__2921 (
            .O(N__19177),
            .I(N__19171));
    InMux I__2920 (
            .O(N__19176),
            .I(N__19171));
    LocalMux I__2919 (
            .O(N__19171),
            .I(\POWERLED.count_off_1_11 ));
    InMux I__2918 (
            .O(N__19168),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    InMux I__2917 (
            .O(N__19165),
            .I(N__19161));
    InMux I__2916 (
            .O(N__19164),
            .I(N__19158));
    LocalMux I__2915 (
            .O(N__19161),
            .I(\POWERLED.count_offZ0Z_12 ));
    LocalMux I__2914 (
            .O(N__19158),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__2913 (
            .O(N__19153),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__2912 (
            .O(N__19150),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__2911 (
            .O(N__19147),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__2910 (
            .O(N__19144),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__2909 (
            .O(N__19141),
            .I(N__19137));
    InMux I__2908 (
            .O(N__19140),
            .I(N__19134));
    LocalMux I__2907 (
            .O(N__19137),
            .I(\POWERLED.count_off_1_12 ));
    LocalMux I__2906 (
            .O(N__19134),
            .I(\POWERLED.count_off_1_12 ));
    InMux I__2905 (
            .O(N__19129),
            .I(N__19126));
    LocalMux I__2904 (
            .O(N__19126),
            .I(\POWERLED.count_off_0_12 ));
    InMux I__2903 (
            .O(N__19123),
            .I(\POWERLED.un3_count_off_1_cry_1 ));
    InMux I__2902 (
            .O(N__19120),
            .I(N__19116));
    InMux I__2901 (
            .O(N__19119),
            .I(N__19113));
    LocalMux I__2900 (
            .O(N__19116),
            .I(N__19110));
    LocalMux I__2899 (
            .O(N__19113),
            .I(\POWERLED.count_offZ0Z_3 ));
    Odrv4 I__2898 (
            .O(N__19110),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__2897 (
            .O(N__19105),
            .I(N__19099));
    InMux I__2896 (
            .O(N__19104),
            .I(N__19099));
    LocalMux I__2895 (
            .O(N__19099),
            .I(N__19096));
    Odrv4 I__2894 (
            .O(N__19096),
            .I(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ));
    InMux I__2893 (
            .O(N__19093),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    InMux I__2892 (
            .O(N__19090),
            .I(N__19086));
    InMux I__2891 (
            .O(N__19089),
            .I(N__19083));
    LocalMux I__2890 (
            .O(N__19086),
            .I(N__19078));
    LocalMux I__2889 (
            .O(N__19083),
            .I(N__19078));
    Odrv4 I__2888 (
            .O(N__19078),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__2887 (
            .O(N__19075),
            .I(N__19069));
    InMux I__2886 (
            .O(N__19074),
            .I(N__19069));
    LocalMux I__2885 (
            .O(N__19069),
            .I(N__19066));
    Odrv4 I__2884 (
            .O(N__19066),
            .I(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ));
    InMux I__2883 (
            .O(N__19063),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    InMux I__2882 (
            .O(N__19060),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    InMux I__2881 (
            .O(N__19057),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    InMux I__2880 (
            .O(N__19054),
            .I(N__19050));
    InMux I__2879 (
            .O(N__19053),
            .I(N__19047));
    LocalMux I__2878 (
            .O(N__19050),
            .I(N__19044));
    LocalMux I__2877 (
            .O(N__19047),
            .I(\POWERLED.count_offZ0Z_7 ));
    Odrv12 I__2876 (
            .O(N__19044),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__2875 (
            .O(N__19039),
            .I(N__19033));
    InMux I__2874 (
            .O(N__19038),
            .I(N__19033));
    LocalMux I__2873 (
            .O(N__19033),
            .I(N__19030));
    Odrv4 I__2872 (
            .O(N__19030),
            .I(\POWERLED.count_off_1_7 ));
    InMux I__2871 (
            .O(N__19027),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__2870 (
            .O(N__19024),
            .I(N__19021));
    LocalMux I__2869 (
            .O(N__19021),
            .I(N__19018));
    Odrv4 I__2868 (
            .O(N__19018),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__2867 (
            .O(N__19015),
            .I(N__19012));
    LocalMux I__2866 (
            .O(N__19012),
            .I(N__19008));
    InMux I__2865 (
            .O(N__19011),
            .I(N__19005));
    Span4Mux_s3_h I__2864 (
            .O(N__19008),
            .I(N__19000));
    LocalMux I__2863 (
            .O(N__19005),
            .I(N__19000));
    Odrv4 I__2862 (
            .O(N__19000),
            .I(\POWERLED.count_off_1_8 ));
    InMux I__2861 (
            .O(N__18997),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__2860 (
            .O(N__18994),
            .I(N__18991));
    LocalMux I__2859 (
            .O(N__18991),
            .I(\POWERLED.count_offZ0Z_9 ));
    InMux I__2858 (
            .O(N__18988),
            .I(N__18982));
    InMux I__2857 (
            .O(N__18987),
            .I(N__18982));
    LocalMux I__2856 (
            .O(N__18982),
            .I(\POWERLED.count_off_1_9 ));
    InMux I__2855 (
            .O(N__18979),
            .I(bfn_6_5_0_));
    CascadeMux I__2854 (
            .O(N__18976),
            .I(N__18973));
    InMux I__2853 (
            .O(N__18973),
            .I(N__18970));
    LocalMux I__2852 (
            .O(N__18970),
            .I(N__18967));
    Odrv4 I__2851 (
            .O(N__18967),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__2850 (
            .O(N__18964),
            .I(bfn_6_3_0_));
    InMux I__2849 (
            .O(N__18961),
            .I(N__18957));
    InMux I__2848 (
            .O(N__18960),
            .I(N__18954));
    LocalMux I__2847 (
            .O(N__18957),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__2846 (
            .O(N__18954),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__2845 (
            .O(N__18949),
            .I(N__18945));
    InMux I__2844 (
            .O(N__18948),
            .I(N__18942));
    LocalMux I__2843 (
            .O(N__18945),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__2842 (
            .O(N__18942),
            .I(\COUNTER.counterZ0Z_22 ));
    CascadeMux I__2841 (
            .O(N__18937),
            .I(N__18933));
    InMux I__2840 (
            .O(N__18936),
            .I(N__18930));
    InMux I__2839 (
            .O(N__18933),
            .I(N__18927));
    LocalMux I__2838 (
            .O(N__18930),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__2837 (
            .O(N__18927),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__2836 (
            .O(N__18922),
            .I(N__18918));
    InMux I__2835 (
            .O(N__18921),
            .I(N__18915));
    LocalMux I__2834 (
            .O(N__18918),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__2833 (
            .O(N__18915),
            .I(\COUNTER.counterZ0Z_20 ));
    CascadeMux I__2832 (
            .O(N__18910),
            .I(N__18907));
    InMux I__2831 (
            .O(N__18907),
            .I(N__18904));
    LocalMux I__2830 (
            .O(N__18904),
            .I(\COUNTER.un4_counter_5_and ));
    InMux I__2829 (
            .O(N__18901),
            .I(N__18897));
    InMux I__2828 (
            .O(N__18900),
            .I(N__18894));
    LocalMux I__2827 (
            .O(N__18897),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__2826 (
            .O(N__18894),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__2825 (
            .O(N__18889),
            .I(N__18885));
    InMux I__2824 (
            .O(N__18888),
            .I(N__18882));
    LocalMux I__2823 (
            .O(N__18885),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__2822 (
            .O(N__18882),
            .I(\COUNTER.counterZ0Z_27 ));
    CascadeMux I__2821 (
            .O(N__18877),
            .I(N__18873));
    InMux I__2820 (
            .O(N__18876),
            .I(N__18870));
    InMux I__2819 (
            .O(N__18873),
            .I(N__18867));
    LocalMux I__2818 (
            .O(N__18870),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__2817 (
            .O(N__18867),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__2816 (
            .O(N__18862),
            .I(N__18858));
    InMux I__2815 (
            .O(N__18861),
            .I(N__18855));
    LocalMux I__2814 (
            .O(N__18858),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__2813 (
            .O(N__18855),
            .I(\COUNTER.counterZ0Z_25 ));
    CascadeMux I__2812 (
            .O(N__18850),
            .I(N__18847));
    InMux I__2811 (
            .O(N__18847),
            .I(N__18844));
    LocalMux I__2810 (
            .O(N__18844),
            .I(\COUNTER.un4_counter_6_and ));
    InMux I__2809 (
            .O(N__18841),
            .I(N__18837));
    InMux I__2808 (
            .O(N__18840),
            .I(N__18834));
    LocalMux I__2807 (
            .O(N__18837),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__2806 (
            .O(N__18834),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__2805 (
            .O(N__18829),
            .I(N__18825));
    InMux I__2804 (
            .O(N__18828),
            .I(N__18822));
    LocalMux I__2803 (
            .O(N__18825),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__2802 (
            .O(N__18822),
            .I(\COUNTER.counterZ0Z_18 ));
    CascadeMux I__2801 (
            .O(N__18817),
            .I(N__18813));
    InMux I__2800 (
            .O(N__18816),
            .I(N__18810));
    InMux I__2799 (
            .O(N__18813),
            .I(N__18807));
    LocalMux I__2798 (
            .O(N__18810),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__2797 (
            .O(N__18807),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__2796 (
            .O(N__18802),
            .I(N__18798));
    InMux I__2795 (
            .O(N__18801),
            .I(N__18795));
    LocalMux I__2794 (
            .O(N__18798),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__2793 (
            .O(N__18795),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__2792 (
            .O(N__18790),
            .I(N__18787));
    InMux I__2791 (
            .O(N__18787),
            .I(N__18784));
    LocalMux I__2790 (
            .O(N__18784),
            .I(\COUNTER.un4_counter_4_and ));
    IoInMux I__2789 (
            .O(N__18781),
            .I(N__18778));
    LocalMux I__2788 (
            .O(N__18778),
            .I(N__18775));
    Span4Mux_s1_h I__2787 (
            .O(N__18775),
            .I(N__18772));
    Span4Mux_h I__2786 (
            .O(N__18772),
            .I(N__18768));
    IoInMux I__2785 (
            .O(N__18771),
            .I(N__18765));
    Span4Mux_v I__2784 (
            .O(N__18768),
            .I(N__18761));
    LocalMux I__2783 (
            .O(N__18765),
            .I(N__18758));
    InMux I__2782 (
            .O(N__18764),
            .I(N__18754));
    Span4Mux_v I__2781 (
            .O(N__18761),
            .I(N__18750));
    IoSpan4Mux I__2780 (
            .O(N__18758),
            .I(N__18747));
    InMux I__2779 (
            .O(N__18757),
            .I(N__18744));
    LocalMux I__2778 (
            .O(N__18754),
            .I(N__18741));
    InMux I__2777 (
            .O(N__18753),
            .I(N__18738));
    Span4Mux_v I__2776 (
            .O(N__18750),
            .I(N__18731));
    Span4Mux_s2_v I__2775 (
            .O(N__18747),
            .I(N__18731));
    LocalMux I__2774 (
            .O(N__18744),
            .I(N__18731));
    Span4Mux_s2_v I__2773 (
            .O(N__18741),
            .I(N__18726));
    LocalMux I__2772 (
            .O(N__18738),
            .I(N__18726));
    Odrv4 I__2771 (
            .O(N__18731),
            .I(pch_pwrok));
    Odrv4 I__2770 (
            .O(N__18726),
            .I(pch_pwrok));
    IoInMux I__2769 (
            .O(N__18721),
            .I(N__18718));
    LocalMux I__2768 (
            .O(N__18718),
            .I(N__18715));
    Odrv12 I__2767 (
            .O(N__18715),
            .I(vccst_pwrgd));
    CascadeMux I__2766 (
            .O(N__18712),
            .I(\POWERLED.mult1_un138_sum_s_8_cascade_ ));
    InMux I__2765 (
            .O(N__18709),
            .I(N__18706));
    LocalMux I__2764 (
            .O(N__18706),
            .I(N__18703));
    Span4Mux_v I__2763 (
            .O(N__18703),
            .I(N__18700));
    Odrv4 I__2762 (
            .O(N__18700),
            .I(\POWERLED.un85_clk_100khz_4 ));
    InMux I__2761 (
            .O(N__18697),
            .I(N__18693));
    InMux I__2760 (
            .O(N__18696),
            .I(N__18690));
    LocalMux I__2759 (
            .O(N__18693),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__2758 (
            .O(N__18690),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__2757 (
            .O(N__18685),
            .I(N__18681));
    InMux I__2756 (
            .O(N__18684),
            .I(N__18678));
    LocalMux I__2755 (
            .O(N__18681),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__2754 (
            .O(N__18678),
            .I(\COUNTER.counterZ0Z_10 ));
    CascadeMux I__2753 (
            .O(N__18673),
            .I(N__18669));
    InMux I__2752 (
            .O(N__18672),
            .I(N__18666));
    InMux I__2751 (
            .O(N__18669),
            .I(N__18663));
    LocalMux I__2750 (
            .O(N__18666),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__2749 (
            .O(N__18663),
            .I(\COUNTER.counterZ0Z_9 ));
    InMux I__2748 (
            .O(N__18658),
            .I(N__18654));
    InMux I__2747 (
            .O(N__18657),
            .I(N__18651));
    LocalMux I__2746 (
            .O(N__18654),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__2745 (
            .O(N__18651),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__2744 (
            .O(N__18646),
            .I(N__18642));
    InMux I__2743 (
            .O(N__18645),
            .I(N__18639));
    LocalMux I__2742 (
            .O(N__18642),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__2741 (
            .O(N__18639),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__2740 (
            .O(N__18634),
            .I(N__18630));
    InMux I__2739 (
            .O(N__18633),
            .I(N__18627));
    LocalMux I__2738 (
            .O(N__18630),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__2737 (
            .O(N__18627),
            .I(\COUNTER.counterZ0Z_13 ));
    CascadeMux I__2736 (
            .O(N__18622),
            .I(N__18618));
    InMux I__2735 (
            .O(N__18621),
            .I(N__18615));
    InMux I__2734 (
            .O(N__18618),
            .I(N__18612));
    LocalMux I__2733 (
            .O(N__18615),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__2732 (
            .O(N__18612),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__2731 (
            .O(N__18607),
            .I(N__18603));
    InMux I__2730 (
            .O(N__18606),
            .I(N__18600));
    LocalMux I__2729 (
            .O(N__18603),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__2728 (
            .O(N__18600),
            .I(\COUNTER.counterZ0Z_15 ));
    CascadeMux I__2727 (
            .O(N__18595),
            .I(N__18592));
    InMux I__2726 (
            .O(N__18592),
            .I(N__18589));
    LocalMux I__2725 (
            .O(N__18589),
            .I(N__18586));
    Odrv4 I__2724 (
            .O(N__18586),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__2723 (
            .O(N__18583),
            .I(N__18580));
    InMux I__2722 (
            .O(N__18580),
            .I(N__18577));
    LocalMux I__2721 (
            .O(N__18577),
            .I(N__18574));
    Odrv4 I__2720 (
            .O(N__18574),
            .I(\COUNTER.un4_counter_1_and ));
    CascadeMux I__2719 (
            .O(N__18571),
            .I(N__18568));
    InMux I__2718 (
            .O(N__18568),
            .I(N__18565));
    LocalMux I__2717 (
            .O(N__18565),
            .I(\COUNTER.un4_counter_2_and ));
    CascadeMux I__2716 (
            .O(N__18562),
            .I(N__18559));
    InMux I__2715 (
            .O(N__18559),
            .I(N__18556));
    LocalMux I__2714 (
            .O(N__18556),
            .I(\COUNTER.un4_counter_3_and ));
    InMux I__2713 (
            .O(N__18553),
            .I(N__18549));
    CascadeMux I__2712 (
            .O(N__18552),
            .I(N__18546));
    LocalMux I__2711 (
            .O(N__18549),
            .I(N__18540));
    InMux I__2710 (
            .O(N__18546),
            .I(N__18533));
    InMux I__2709 (
            .O(N__18545),
            .I(N__18533));
    InMux I__2708 (
            .O(N__18544),
            .I(N__18533));
    InMux I__2707 (
            .O(N__18543),
            .I(N__18530));
    Odrv4 I__2706 (
            .O(N__18540),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__2705 (
            .O(N__18533),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__2704 (
            .O(N__18530),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    CascadeMux I__2703 (
            .O(N__18523),
            .I(N__18519));
    InMux I__2702 (
            .O(N__18522),
            .I(N__18511));
    InMux I__2701 (
            .O(N__18519),
            .I(N__18511));
    InMux I__2700 (
            .O(N__18518),
            .I(N__18511));
    LocalMux I__2699 (
            .O(N__18511),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    InMux I__2698 (
            .O(N__18508),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    InMux I__2697 (
            .O(N__18505),
            .I(N__18502));
    LocalMux I__2696 (
            .O(N__18502),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__2695 (
            .O(N__18499),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    CascadeMux I__2694 (
            .O(N__18496),
            .I(N__18493));
    InMux I__2693 (
            .O(N__18493),
            .I(N__18490));
    LocalMux I__2692 (
            .O(N__18490),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__2691 (
            .O(N__18487),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    InMux I__2690 (
            .O(N__18484),
            .I(N__18481));
    LocalMux I__2689 (
            .O(N__18481),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__2688 (
            .O(N__18478),
            .I(N__18475));
    LocalMux I__2687 (
            .O(N__18475),
            .I(N__18471));
    CascadeMux I__2686 (
            .O(N__18474),
            .I(N__18468));
    Span4Mux_s2_v I__2685 (
            .O(N__18471),
            .I(N__18462));
    InMux I__2684 (
            .O(N__18468),
            .I(N__18457));
    InMux I__2683 (
            .O(N__18467),
            .I(N__18457));
    InMux I__2682 (
            .O(N__18466),
            .I(N__18454));
    InMux I__2681 (
            .O(N__18465),
            .I(N__18451));
    Odrv4 I__2680 (
            .O(N__18462),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2679 (
            .O(N__18457),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2678 (
            .O(N__18454),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__2677 (
            .O(N__18451),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    InMux I__2676 (
            .O(N__18442),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    CascadeMux I__2675 (
            .O(N__18439),
            .I(N__18435));
    InMux I__2674 (
            .O(N__18438),
            .I(N__18427));
    InMux I__2673 (
            .O(N__18435),
            .I(N__18427));
    InMux I__2672 (
            .O(N__18434),
            .I(N__18427));
    LocalMux I__2671 (
            .O(N__18427),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    CascadeMux I__2670 (
            .O(N__18424),
            .I(N__18421));
    InMux I__2669 (
            .O(N__18421),
            .I(N__18418));
    LocalMux I__2668 (
            .O(N__18418),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__2667 (
            .O(N__18415),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__2666 (
            .O(N__18412),
            .I(N__18409));
    LocalMux I__2665 (
            .O(N__18409),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__2664 (
            .O(N__18406),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    InMux I__2663 (
            .O(N__18403),
            .I(N__18400));
    LocalMux I__2662 (
            .O(N__18400),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__2661 (
            .O(N__18397),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    CascadeMux I__2660 (
            .O(N__18394),
            .I(N__18390));
    InMux I__2659 (
            .O(N__18393),
            .I(N__18382));
    InMux I__2658 (
            .O(N__18390),
            .I(N__18382));
    InMux I__2657 (
            .O(N__18389),
            .I(N__18382));
    LocalMux I__2656 (
            .O(N__18382),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__2655 (
            .O(N__18379),
            .I(N__18376));
    InMux I__2654 (
            .O(N__18376),
            .I(N__18373));
    LocalMux I__2653 (
            .O(N__18373),
            .I(N__18370));
    Odrv4 I__2652 (
            .O(N__18370),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__2651 (
            .O(N__18367),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    InMux I__2650 (
            .O(N__18364),
            .I(N__18361));
    LocalMux I__2649 (
            .O(N__18361),
            .I(N__18358));
    Odrv4 I__2648 (
            .O(N__18358),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__2647 (
            .O(N__18355),
            .I(N__18352));
    LocalMux I__2646 (
            .O(N__18352),
            .I(N__18349));
    Odrv4 I__2645 (
            .O(N__18349),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__2644 (
            .O(N__18346),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    CascadeMux I__2643 (
            .O(N__18343),
            .I(N__18340));
    InMux I__2642 (
            .O(N__18340),
            .I(N__18337));
    LocalMux I__2641 (
            .O(N__18337),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    CascadeMux I__2640 (
            .O(N__18334),
            .I(N__18331));
    InMux I__2639 (
            .O(N__18331),
            .I(N__18328));
    LocalMux I__2638 (
            .O(N__18328),
            .I(N__18325));
    Odrv4 I__2637 (
            .O(N__18325),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__2636 (
            .O(N__18322),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__2635 (
            .O(N__18319),
            .I(N__18316));
    LocalMux I__2634 (
            .O(N__18316),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    CascadeMux I__2633 (
            .O(N__18313),
            .I(N__18310));
    InMux I__2632 (
            .O(N__18310),
            .I(N__18307));
    LocalMux I__2631 (
            .O(N__18307),
            .I(N__18304));
    Odrv4 I__2630 (
            .O(N__18304),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__2629 (
            .O(N__18301),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    CascadeMux I__2628 (
            .O(N__18298),
            .I(N__18295));
    InMux I__2627 (
            .O(N__18295),
            .I(N__18292));
    LocalMux I__2626 (
            .O(N__18292),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__2625 (
            .O(N__18289),
            .I(N__18286));
    LocalMux I__2624 (
            .O(N__18286),
            .I(N__18283));
    Odrv4 I__2623 (
            .O(N__18283),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__2622 (
            .O(N__18280),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__2621 (
            .O(N__18277),
            .I(N__18274));
    LocalMux I__2620 (
            .O(N__18274),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__2619 (
            .O(N__18271),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    InMux I__2618 (
            .O(N__18268),
            .I(N__18264));
    CascadeMux I__2617 (
            .O(N__18267),
            .I(N__18260));
    LocalMux I__2616 (
            .O(N__18264),
            .I(N__18257));
    InMux I__2615 (
            .O(N__18263),
            .I(N__18252));
    InMux I__2614 (
            .O(N__18260),
            .I(N__18252));
    Span4Mux_s2_v I__2613 (
            .O(N__18257),
            .I(N__18247));
    LocalMux I__2612 (
            .O(N__18252),
            .I(N__18244));
    InMux I__2611 (
            .O(N__18251),
            .I(N__18241));
    InMux I__2610 (
            .O(N__18250),
            .I(N__18238));
    Odrv4 I__2609 (
            .O(N__18247),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    Odrv4 I__2608 (
            .O(N__18244),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2607 (
            .O(N__18241),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__2606 (
            .O(N__18238),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    InMux I__2605 (
            .O(N__18229),
            .I(N__18226));
    LocalMux I__2604 (
            .O(N__18226),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__2603 (
            .O(N__18223),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__2602 (
            .O(N__18220),
            .I(N__18215));
    InMux I__2601 (
            .O(N__18219),
            .I(N__18211));
    InMux I__2600 (
            .O(N__18218),
            .I(N__18206));
    InMux I__2599 (
            .O(N__18215),
            .I(N__18206));
    InMux I__2598 (
            .O(N__18214),
            .I(N__18203));
    LocalMux I__2597 (
            .O(N__18211),
            .I(N__18200));
    LocalMux I__2596 (
            .O(N__18206),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__2595 (
            .O(N__18203),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    Odrv4 I__2594 (
            .O(N__18200),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__2593 (
            .O(N__18193),
            .I(N__18189));
    CascadeMux I__2592 (
            .O(N__18192),
            .I(N__18185));
    InMux I__2591 (
            .O(N__18189),
            .I(N__18178));
    InMux I__2590 (
            .O(N__18188),
            .I(N__18178));
    InMux I__2589 (
            .O(N__18185),
            .I(N__18178));
    LocalMux I__2588 (
            .O(N__18178),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    InMux I__2587 (
            .O(N__18175),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    InMux I__2586 (
            .O(N__18172),
            .I(N__18169));
    LocalMux I__2585 (
            .O(N__18169),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__2584 (
            .O(N__18166),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__2583 (
            .O(N__18163),
            .I(N__18160));
    LocalMux I__2582 (
            .O(N__18160),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__2581 (
            .O(N__18157),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__2580 (
            .O(N__18154),
            .I(N__18151));
    LocalMux I__2579 (
            .O(N__18151),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__2578 (
            .O(N__18148),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    CascadeMux I__2577 (
            .O(N__18145),
            .I(N__18142));
    InMux I__2576 (
            .O(N__18142),
            .I(N__18139));
    LocalMux I__2575 (
            .O(N__18139),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__2574 (
            .O(N__18136),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__2573 (
            .O(N__18133),
            .I(N__18130));
    LocalMux I__2572 (
            .O(N__18130),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    InMux I__2571 (
            .O(N__18127),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__2570 (
            .O(N__18124),
            .I(N__18121));
    InMux I__2569 (
            .O(N__18121),
            .I(N__18118));
    LocalMux I__2568 (
            .O(N__18118),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__2567 (
            .O(N__18115),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__2566 (
            .O(N__18112),
            .I(\POWERLED.mult1_un61_sum_s_8_cascade_ ));
    InMux I__2565 (
            .O(N__18109),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    CascadeMux I__2564 (
            .O(N__18106),
            .I(N__18103));
    InMux I__2563 (
            .O(N__18103),
            .I(N__18100));
    LocalMux I__2562 (
            .O(N__18100),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__2561 (
            .O(N__18097),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    InMux I__2560 (
            .O(N__18094),
            .I(N__18091));
    LocalMux I__2559 (
            .O(N__18091),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__2558 (
            .O(N__18088),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__2557 (
            .O(N__18085),
            .I(N__18082));
    LocalMux I__2556 (
            .O(N__18082),
            .I(N__18079));
    Span4Mux_s2_v I__2555 (
            .O(N__18079),
            .I(N__18075));
    CascadeMux I__2554 (
            .O(N__18078),
            .I(N__18071));
    Span4Mux_h I__2553 (
            .O(N__18075),
            .I(N__18067));
    InMux I__2552 (
            .O(N__18074),
            .I(N__18062));
    InMux I__2551 (
            .O(N__18071),
            .I(N__18062));
    InMux I__2550 (
            .O(N__18070),
            .I(N__18059));
    Odrv4 I__2549 (
            .O(N__18067),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__2548 (
            .O(N__18062),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__2547 (
            .O(N__18059),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__2546 (
            .O(N__18052),
            .I(N__18049));
    InMux I__2545 (
            .O(N__18049),
            .I(N__18046));
    LocalMux I__2544 (
            .O(N__18046),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__2543 (
            .O(N__18043),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    InMux I__2542 (
            .O(N__18040),
            .I(N__18037));
    LocalMux I__2541 (
            .O(N__18037),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    CascadeMux I__2540 (
            .O(N__18034),
            .I(N__18030));
    CascadeMux I__2539 (
            .O(N__18033),
            .I(N__18026));
    InMux I__2538 (
            .O(N__18030),
            .I(N__18019));
    InMux I__2537 (
            .O(N__18029),
            .I(N__18019));
    InMux I__2536 (
            .O(N__18026),
            .I(N__18019));
    LocalMux I__2535 (
            .O(N__18019),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__2534 (
            .O(N__18016),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    CascadeMux I__2533 (
            .O(N__18013),
            .I(N__18010));
    InMux I__2532 (
            .O(N__18010),
            .I(N__18007));
    LocalMux I__2531 (
            .O(N__18007),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    InMux I__2530 (
            .O(N__18004),
            .I(N__17999));
    InMux I__2529 (
            .O(N__18003),
            .I(N__17996));
    InMux I__2528 (
            .O(N__18002),
            .I(N__17993));
    LocalMux I__2527 (
            .O(N__17999),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__2526 (
            .O(N__17996),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__2525 (
            .O(N__17993),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    CascadeMux I__2524 (
            .O(N__17986),
            .I(N__17983));
    InMux I__2523 (
            .O(N__17983),
            .I(N__17980));
    LocalMux I__2522 (
            .O(N__17980),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    CascadeMux I__2521 (
            .O(N__17977),
            .I(N__17974));
    InMux I__2520 (
            .O(N__17974),
            .I(N__17971));
    LocalMux I__2519 (
            .O(N__17971),
            .I(\POWERLED.mult1_un47_sum_s_4_sf ));
    CascadeMux I__2518 (
            .O(N__17968),
            .I(N__17965));
    InMux I__2517 (
            .O(N__17965),
            .I(N__17962));
    LocalMux I__2516 (
            .O(N__17962),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    InMux I__2515 (
            .O(N__17959),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__2514 (
            .O(N__17956),
            .I(N__17953));
    InMux I__2513 (
            .O(N__17953),
            .I(N__17950));
    LocalMux I__2512 (
            .O(N__17950),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__2511 (
            .O(N__17947),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__2510 (
            .O(N__17944),
            .I(N__17941));
    LocalMux I__2509 (
            .O(N__17941),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__2508 (
            .O(N__17938),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__2507 (
            .O(N__17935),
            .I(N__17932));
    InMux I__2506 (
            .O(N__17932),
            .I(N__17929));
    LocalMux I__2505 (
            .O(N__17929),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__2504 (
            .O(N__17926),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    CascadeMux I__2503 (
            .O(N__17923),
            .I(N__17920));
    InMux I__2502 (
            .O(N__17920),
            .I(N__17917));
    LocalMux I__2501 (
            .O(N__17917),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__2500 (
            .O(N__17914),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__2499 (
            .O(N__17911),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    InMux I__2498 (
            .O(N__17908),
            .I(N__17904));
    InMux I__2497 (
            .O(N__17907),
            .I(N__17901));
    LocalMux I__2496 (
            .O(N__17904),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    LocalMux I__2495 (
            .O(N__17901),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    CascadeMux I__2494 (
            .O(N__17896),
            .I(N__17893));
    InMux I__2493 (
            .O(N__17893),
            .I(N__17890));
    LocalMux I__2492 (
            .O(N__17890),
            .I(\POWERLED.un1_dutycycle_53_4_3 ));
    InMux I__2491 (
            .O(N__17887),
            .I(N__17884));
    LocalMux I__2490 (
            .O(N__17884),
            .I(N__17879));
    CascadeMux I__2489 (
            .O(N__17883),
            .I(N__17876));
    CascadeMux I__2488 (
            .O(N__17882),
            .I(N__17873));
    Span4Mux_v I__2487 (
            .O(N__17879),
            .I(N__17869));
    InMux I__2486 (
            .O(N__17876),
            .I(N__17862));
    InMux I__2485 (
            .O(N__17873),
            .I(N__17862));
    InMux I__2484 (
            .O(N__17872),
            .I(N__17862));
    Span4Mux_h I__2483 (
            .O(N__17869),
            .I(N__17857));
    LocalMux I__2482 (
            .O(N__17862),
            .I(N__17857));
    Span4Mux_s1_h I__2481 (
            .O(N__17857),
            .I(N__17854));
    Odrv4 I__2480 (
            .O(N__17854),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    CascadeMux I__2479 (
            .O(N__17851),
            .I(N__17848));
    InMux I__2478 (
            .O(N__17848),
            .I(N__17845));
    LocalMux I__2477 (
            .O(N__17845),
            .I(N__17840));
    InMux I__2476 (
            .O(N__17844),
            .I(N__17836));
    InMux I__2475 (
            .O(N__17843),
            .I(N__17833));
    Span4Mux_h I__2474 (
            .O(N__17840),
            .I(N__17830));
    InMux I__2473 (
            .O(N__17839),
            .I(N__17827));
    LocalMux I__2472 (
            .O(N__17836),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    LocalMux I__2471 (
            .O(N__17833),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    Odrv4 I__2470 (
            .O(N__17830),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    LocalMux I__2469 (
            .O(N__17827),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    InMux I__2468 (
            .O(N__17818),
            .I(N__17815));
    LocalMux I__2467 (
            .O(N__17815),
            .I(N__17808));
    InMux I__2466 (
            .O(N__17814),
            .I(N__17803));
    InMux I__2465 (
            .O(N__17813),
            .I(N__17803));
    InMux I__2464 (
            .O(N__17812),
            .I(N__17798));
    InMux I__2463 (
            .O(N__17811),
            .I(N__17798));
    Span4Mux_h I__2462 (
            .O(N__17808),
            .I(N__17795));
    LocalMux I__2461 (
            .O(N__17803),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__2460 (
            .O(N__17798),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__2459 (
            .O(N__17795),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    InMux I__2458 (
            .O(N__17788),
            .I(N__17785));
    LocalMux I__2457 (
            .O(N__17785),
            .I(N__17782));
    Span12Mux_s6_v I__2456 (
            .O(N__17782),
            .I(N__17779));
    Odrv12 I__2455 (
            .O(N__17779),
            .I(\POWERLED.curr_state_1_0 ));
    InMux I__2454 (
            .O(N__17776),
            .I(N__17773));
    LocalMux I__2453 (
            .O(N__17773),
            .I(N__17770));
    Odrv4 I__2452 (
            .O(N__17770),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_10 ));
    InMux I__2451 (
            .O(N__17767),
            .I(N__17764));
    LocalMux I__2450 (
            .O(N__17764),
            .I(N__17761));
    Odrv4 I__2449 (
            .O(N__17761),
            .I(\POWERLED.dutycycle_RNI_9Z0Z_9 ));
    CascadeMux I__2448 (
            .O(N__17758),
            .I(N__17755));
    InMux I__2447 (
            .O(N__17755),
            .I(N__17751));
    InMux I__2446 (
            .O(N__17754),
            .I(N__17748));
    LocalMux I__2445 (
            .O(N__17751),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    LocalMux I__2444 (
            .O(N__17748),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    CascadeMux I__2443 (
            .O(N__17743),
            .I(\POWERLED.dutycycle_en_12_cascade_ ));
    InMux I__2442 (
            .O(N__17740),
            .I(N__17737));
    LocalMux I__2441 (
            .O(N__17737),
            .I(\POWERLED.un1_clk_100khz_48_and_i_i_a3_0_0 ));
    InMux I__2440 (
            .O(N__17734),
            .I(N__17731));
    LocalMux I__2439 (
            .O(N__17731),
            .I(\POWERLED.dutycycle_en_12 ));
    CascadeMux I__2438 (
            .O(N__17728),
            .I(N__17724));
    InMux I__2437 (
            .O(N__17727),
            .I(N__17719));
    InMux I__2436 (
            .O(N__17724),
            .I(N__17719));
    LocalMux I__2435 (
            .O(N__17719),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    CascadeMux I__2434 (
            .O(N__17716),
            .I(\POWERLED.dutycycleZ0Z_13_cascade_ ));
    CascadeMux I__2433 (
            .O(N__17713),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_15_cascade_ ));
    CascadeMux I__2432 (
            .O(N__17710),
            .I(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ));
    CascadeMux I__2431 (
            .O(N__17707),
            .I(N__17704));
    InMux I__2430 (
            .O(N__17704),
            .I(N__17697));
    InMux I__2429 (
            .O(N__17703),
            .I(N__17697));
    InMux I__2428 (
            .O(N__17702),
            .I(N__17694));
    LocalMux I__2427 (
            .O(N__17697),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__2426 (
            .O(N__17694),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    InMux I__2425 (
            .O(N__17689),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__2424 (
            .O(N__17686),
            .I(N__17683));
    InMux I__2423 (
            .O(N__17683),
            .I(N__17680));
    LocalMux I__2422 (
            .O(N__17680),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__2421 (
            .O(N__17677),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__2420 (
            .O(N__17674),
            .I(\POWERLED.dutycycle_eena_5_cascade_ ));
    CascadeMux I__2419 (
            .O(N__17671),
            .I(\POWERLED.dutycycleZ1Z_5_cascade_ ));
    InMux I__2418 (
            .O(N__17668),
            .I(N__17665));
    LocalMux I__2417 (
            .O(N__17665),
            .I(\POWERLED.dutycycle_eena_5_1 ));
    CascadeMux I__2416 (
            .O(N__17662),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    CascadeMux I__2415 (
            .O(N__17659),
            .I(\POWERLED.dutycycle_eena_6_1_cascade_ ));
    InMux I__2414 (
            .O(N__17656),
            .I(N__17653));
    LocalMux I__2413 (
            .O(N__17653),
            .I(\POWERLED.dutycycle_eena_6 ));
    CascadeMux I__2412 (
            .O(N__17650),
            .I(\POWERLED.dutycycle_eena_6_cascade_ ));
    InMux I__2411 (
            .O(N__17647),
            .I(N__17643));
    InMux I__2410 (
            .O(N__17646),
            .I(N__17640));
    LocalMux I__2409 (
            .O(N__17643),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    LocalMux I__2408 (
            .O(N__17640),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    InMux I__2407 (
            .O(N__17635),
            .I(N__17632));
    LocalMux I__2406 (
            .O(N__17632),
            .I(\POWERLED.dutycycle_eena_5 ));
    InMux I__2405 (
            .O(N__17629),
            .I(N__17623));
    InMux I__2404 (
            .O(N__17628),
            .I(N__17623));
    LocalMux I__2403 (
            .O(N__17623),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    CascadeMux I__2402 (
            .O(N__17620),
            .I(\POWERLED.N_4_0_cascade_ ));
    CascadeMux I__2401 (
            .O(N__17617),
            .I(\POWERLED.dutycycle_eena_8_1_cascade_ ));
    CascadeMux I__2400 (
            .O(N__17614),
            .I(\POWERLED.dutycycle_eena_8_cascade_ ));
    InMux I__2399 (
            .O(N__17611),
            .I(N__17608));
    LocalMux I__2398 (
            .O(N__17608),
            .I(\POWERLED.dutycycle_eena_8 ));
    InMux I__2397 (
            .O(N__17605),
            .I(N__17599));
    InMux I__2396 (
            .O(N__17604),
            .I(N__17599));
    LocalMux I__2395 (
            .O(N__17599),
            .I(\POWERLED.dutycycleZ1Z_3 ));
    CascadeMux I__2394 (
            .O(N__17596),
            .I(\POWERLED.dutycycleZ0Z_6_cascade_ ));
    CascadeMux I__2393 (
            .O(N__17593),
            .I(\POWERLED.dutycycle_eena_4_1_cascade_ ));
    CascadeMux I__2392 (
            .O(N__17590),
            .I(N__17587));
    InMux I__2391 (
            .O(N__17587),
            .I(N__17584));
    LocalMux I__2390 (
            .O(N__17584),
            .I(\POWERLED.dutycycle_eena_4 ));
    CascadeMux I__2389 (
            .O(N__17581),
            .I(\POWERLED.dutycycle_eena_4_cascade_ ));
    InMux I__2388 (
            .O(N__17578),
            .I(N__17572));
    InMux I__2387 (
            .O(N__17577),
            .I(N__17572));
    LocalMux I__2386 (
            .O(N__17572),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    InMux I__2385 (
            .O(N__17569),
            .I(\COUNTER.counter_1_cry_30 ));
    CascadeMux I__2384 (
            .O(N__17566),
            .I(N__17563));
    InMux I__2383 (
            .O(N__17563),
            .I(N__17557));
    InMux I__2382 (
            .O(N__17562),
            .I(N__17557));
    LocalMux I__2381 (
            .O(N__17557),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__2380 (
            .O(N__17554),
            .I(N__17548));
    InMux I__2379 (
            .O(N__17553),
            .I(N__17548));
    LocalMux I__2378 (
            .O(N__17548),
            .I(\COUNTER.counterZ0Z_31 ));
    CascadeMux I__2377 (
            .O(N__17545),
            .I(N__17541));
    CascadeMux I__2376 (
            .O(N__17544),
            .I(N__17538));
    InMux I__2375 (
            .O(N__17541),
            .I(N__17533));
    InMux I__2374 (
            .O(N__17538),
            .I(N__17533));
    LocalMux I__2373 (
            .O(N__17533),
            .I(\COUNTER.counterZ0Z_30 ));
    CascadeMux I__2372 (
            .O(N__17530),
            .I(N__17527));
    InMux I__2371 (
            .O(N__17527),
            .I(N__17521));
    InMux I__2370 (
            .O(N__17526),
            .I(N__17521));
    LocalMux I__2369 (
            .O(N__17521),
            .I(\COUNTER.counterZ0Z_29 ));
    InMux I__2368 (
            .O(N__17518),
            .I(N__17515));
    LocalMux I__2367 (
            .O(N__17515),
            .I(\POWERLED.count_off_0_9 ));
    CascadeMux I__2366 (
            .O(N__17512),
            .I(\POWERLED.count_offZ0Z_9_cascade_ ));
    InMux I__2365 (
            .O(N__17509),
            .I(N__17506));
    LocalMux I__2364 (
            .O(N__17506),
            .I(\POWERLED.count_off_0_10 ));
    InMux I__2363 (
            .O(N__17503),
            .I(N__17500));
    LocalMux I__2362 (
            .O(N__17500),
            .I(\POWERLED.count_off_0_11 ));
    InMux I__2361 (
            .O(N__17497),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__2360 (
            .O(N__17494),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__2359 (
            .O(N__17491),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__2358 (
            .O(N__17488),
            .I(bfn_5_4_0_));
    InMux I__2357 (
            .O(N__17485),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__2356 (
            .O(N__17482),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__2355 (
            .O(N__17479),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__2354 (
            .O(N__17476),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__2353 (
            .O(N__17473),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__2352 (
            .O(N__17470),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__2351 (
            .O(N__17467),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__2350 (
            .O(N__17464),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__2349 (
            .O(N__17461),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__2348 (
            .O(N__17458),
            .I(bfn_5_3_0_));
    InMux I__2347 (
            .O(N__17455),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__2346 (
            .O(N__17452),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__2345 (
            .O(N__17449),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__2344 (
            .O(N__17446),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__2343 (
            .O(N__17443),
            .I(\COUNTER.counter_1_cry_3 ));
    CascadeMux I__2342 (
            .O(N__17440),
            .I(N__17435));
    InMux I__2341 (
            .O(N__17439),
            .I(N__17432));
    InMux I__2340 (
            .O(N__17438),
            .I(N__17429));
    InMux I__2339 (
            .O(N__17435),
            .I(N__17426));
    LocalMux I__2338 (
            .O(N__17432),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__2337 (
            .O(N__17429),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__2336 (
            .O(N__17426),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__2335 (
            .O(N__17419),
            .I(N__17416));
    LocalMux I__2334 (
            .O(N__17416),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__2333 (
            .O(N__17413),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__2332 (
            .O(N__17410),
            .I(N__17405));
    InMux I__2331 (
            .O(N__17409),
            .I(N__17400));
    InMux I__2330 (
            .O(N__17408),
            .I(N__17400));
    LocalMux I__2329 (
            .O(N__17405),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__2328 (
            .O(N__17400),
            .I(\COUNTER.counterZ0Z_6 ));
    CascadeMux I__2327 (
            .O(N__17395),
            .I(N__17392));
    InMux I__2326 (
            .O(N__17392),
            .I(N__17389));
    LocalMux I__2325 (
            .O(N__17389),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__2324 (
            .O(N__17386),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__2323 (
            .O(N__17383),
            .I(N__17379));
    InMux I__2322 (
            .O(N__17382),
            .I(N__17376));
    LocalMux I__2321 (
            .O(N__17379),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__2320 (
            .O(N__17376),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__2319 (
            .O(N__17371),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__2318 (
            .O(N__17368),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__2317 (
            .O(N__17365),
            .I(bfn_5_2_0_));
    InMux I__2316 (
            .O(N__17362),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__2315 (
            .O(N__17359),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__2314 (
            .O(N__17356),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__2313 (
            .O(N__17353),
            .I(N__17350));
    LocalMux I__2312 (
            .O(N__17350),
            .I(N__17347));
    Odrv4 I__2311 (
            .O(N__17347),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__2310 (
            .O(N__17344),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    CascadeMux I__2309 (
            .O(N__17341),
            .I(N__17338));
    InMux I__2308 (
            .O(N__17338),
            .I(N__17335));
    LocalMux I__2307 (
            .O(N__17335),
            .I(N__17332));
    Odrv4 I__2306 (
            .O(N__17332),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__2305 (
            .O(N__17329),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    CascadeMux I__2304 (
            .O(N__17326),
            .I(N__17323));
    InMux I__2303 (
            .O(N__17323),
            .I(N__17320));
    LocalMux I__2302 (
            .O(N__17320),
            .I(N__17317));
    Odrv4 I__2301 (
            .O(N__17317),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__2300 (
            .O(N__17314),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__2299 (
            .O(N__17311),
            .I(N__17306));
    InMux I__2298 (
            .O(N__17310),
            .I(N__17301));
    InMux I__2297 (
            .O(N__17309),
            .I(N__17301));
    LocalMux I__2296 (
            .O(N__17306),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    LocalMux I__2295 (
            .O(N__17301),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__2294 (
            .O(N__17296),
            .I(N__17293));
    LocalMux I__2293 (
            .O(N__17293),
            .I(N__17290));
    Odrv4 I__2292 (
            .O(N__17290),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__2291 (
            .O(N__17287),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__2290 (
            .O(N__17284),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    InMux I__2289 (
            .O(N__17281),
            .I(N__17276));
    CascadeMux I__2288 (
            .O(N__17280),
            .I(N__17272));
    InMux I__2287 (
            .O(N__17279),
            .I(N__17269));
    LocalMux I__2286 (
            .O(N__17276),
            .I(N__17266));
    InMux I__2285 (
            .O(N__17275),
            .I(N__17261));
    InMux I__2284 (
            .O(N__17272),
            .I(N__17261));
    LocalMux I__2283 (
            .O(N__17269),
            .I(N__17257));
    Span4Mux_v I__2282 (
            .O(N__17266),
            .I(N__17252));
    LocalMux I__2281 (
            .O(N__17261),
            .I(N__17252));
    InMux I__2280 (
            .O(N__17260),
            .I(N__17249));
    Odrv4 I__2279 (
            .O(N__17257),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    Odrv4 I__2278 (
            .O(N__17252),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__2277 (
            .O(N__17249),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    InMux I__2276 (
            .O(N__17242),
            .I(N__17237));
    InMux I__2275 (
            .O(N__17241),
            .I(N__17232));
    InMux I__2274 (
            .O(N__17240),
            .I(N__17232));
    LocalMux I__2273 (
            .O(N__17237),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__2272 (
            .O(N__17232),
            .I(\COUNTER.counterZ0Z_1 ));
    CascadeMux I__2271 (
            .O(N__17227),
            .I(N__17224));
    InMux I__2270 (
            .O(N__17224),
            .I(N__17220));
    InMux I__2269 (
            .O(N__17223),
            .I(N__17216));
    LocalMux I__2268 (
            .O(N__17220),
            .I(N__17213));
    InMux I__2267 (
            .O(N__17219),
            .I(N__17209));
    LocalMux I__2266 (
            .O(N__17216),
            .I(N__17204));
    Span4Mux_s0_v I__2265 (
            .O(N__17213),
            .I(N__17204));
    InMux I__2264 (
            .O(N__17212),
            .I(N__17201));
    LocalMux I__2263 (
            .O(N__17209),
            .I(\COUNTER.counterZ0Z_0 ));
    Odrv4 I__2262 (
            .O(N__17204),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__2261 (
            .O(N__17201),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__2260 (
            .O(N__17194),
            .I(N__17189));
    InMux I__2259 (
            .O(N__17193),
            .I(N__17184));
    InMux I__2258 (
            .O(N__17192),
            .I(N__17184));
    LocalMux I__2257 (
            .O(N__17189),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__2256 (
            .O(N__17184),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__2255 (
            .O(N__17179),
            .I(N__17176));
    LocalMux I__2254 (
            .O(N__17176),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__2253 (
            .O(N__17173),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__2252 (
            .O(N__17170),
            .I(N__17165));
    InMux I__2251 (
            .O(N__17169),
            .I(N__17160));
    InMux I__2250 (
            .O(N__17168),
            .I(N__17160));
    LocalMux I__2249 (
            .O(N__17165),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__2248 (
            .O(N__17160),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__2247 (
            .O(N__17155),
            .I(N__17152));
    LocalMux I__2246 (
            .O(N__17152),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__2245 (
            .O(N__17149),
            .I(\COUNTER.counter_1_cry_2 ));
    CascadeMux I__2244 (
            .O(N__17146),
            .I(N__17141));
    InMux I__2243 (
            .O(N__17145),
            .I(N__17138));
    InMux I__2242 (
            .O(N__17144),
            .I(N__17135));
    InMux I__2241 (
            .O(N__17141),
            .I(N__17132));
    LocalMux I__2240 (
            .O(N__17138),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__2239 (
            .O(N__17135),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__2238 (
            .O(N__17132),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__2237 (
            .O(N__17125),
            .I(N__17122));
    LocalMux I__2236 (
            .O(N__17122),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__2235 (
            .O(N__17119),
            .I(N__17116));
    LocalMux I__2234 (
            .O(N__17116),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__2233 (
            .O(N__17113),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__2232 (
            .O(N__17110),
            .I(N__17107));
    InMux I__2231 (
            .O(N__17107),
            .I(N__17094));
    InMux I__2230 (
            .O(N__17106),
            .I(N__17094));
    InMux I__2229 (
            .O(N__17105),
            .I(N__17094));
    InMux I__2228 (
            .O(N__17104),
            .I(N__17087));
    InMux I__2227 (
            .O(N__17103),
            .I(N__17087));
    InMux I__2226 (
            .O(N__17102),
            .I(N__17087));
    InMux I__2225 (
            .O(N__17101),
            .I(N__17084));
    LocalMux I__2224 (
            .O(N__17094),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2223 (
            .O(N__17087),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__2222 (
            .O(N__17084),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    InMux I__2221 (
            .O(N__17077),
            .I(N__17074));
    LocalMux I__2220 (
            .O(N__17074),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__2219 (
            .O(N__17071),
            .I(N__17068));
    LocalMux I__2218 (
            .O(N__17068),
            .I(N__17065));
    Span4Mux_s3_v I__2217 (
            .O(N__17065),
            .I(N__17062));
    Odrv4 I__2216 (
            .O(N__17062),
            .I(vpp_ok));
    IoInMux I__2215 (
            .O(N__17059),
            .I(N__17056));
    LocalMux I__2214 (
            .O(N__17056),
            .I(N__17053));
    IoSpan4Mux I__2213 (
            .O(N__17053),
            .I(N__17050));
    Odrv4 I__2212 (
            .O(N__17050),
            .I(vddq_en));
    InMux I__2211 (
            .O(N__17047),
            .I(N__17044));
    LocalMux I__2210 (
            .O(N__17044),
            .I(N__17041));
    Span4Mux_s3_h I__2209 (
            .O(N__17041),
            .I(N__17038));
    Odrv4 I__2208 (
            .O(N__17038),
            .I(\POWERLED.mult1_un75_sum_i_8 ));
    CascadeMux I__2207 (
            .O(N__17035),
            .I(N__17032));
    InMux I__2206 (
            .O(N__17032),
            .I(N__17029));
    LocalMux I__2205 (
            .O(N__17029),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__2204 (
            .O(N__17026),
            .I(N__17023));
    LocalMux I__2203 (
            .O(N__17023),
            .I(N__17020));
    Odrv4 I__2202 (
            .O(N__17020),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__2201 (
            .O(N__17017),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__2200 (
            .O(N__17014),
            .I(N__17011));
    LocalMux I__2199 (
            .O(N__17011),
            .I(N__17008));
    Odrv12 I__2198 (
            .O(N__17008),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__2197 (
            .O(N__17005),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    CascadeMux I__2196 (
            .O(N__17002),
            .I(N__16998));
    InMux I__2195 (
            .O(N__17001),
            .I(N__16990));
    InMux I__2194 (
            .O(N__16998),
            .I(N__16990));
    InMux I__2193 (
            .O(N__16997),
            .I(N__16990));
    LocalMux I__2192 (
            .O(N__16990),
            .I(N__16986));
    InMux I__2191 (
            .O(N__16989),
            .I(N__16983));
    Odrv4 I__2190 (
            .O(N__16986),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__2189 (
            .O(N__16983),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    CascadeMux I__2188 (
            .O(N__16978),
            .I(N__16974));
    InMux I__2187 (
            .O(N__16977),
            .I(N__16966));
    InMux I__2186 (
            .O(N__16974),
            .I(N__16966));
    InMux I__2185 (
            .O(N__16973),
            .I(N__16966));
    LocalMux I__2184 (
            .O(N__16966),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    CascadeMux I__2183 (
            .O(N__16963),
            .I(N__16960));
    InMux I__2182 (
            .O(N__16960),
            .I(N__16957));
    LocalMux I__2181 (
            .O(N__16957),
            .I(N__16954));
    Odrv4 I__2180 (
            .O(N__16954),
            .I(\POWERLED.mult1_un124_sum_i ));
    InMux I__2179 (
            .O(N__16951),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__2178 (
            .O(N__16948),
            .I(N__16945));
    LocalMux I__2177 (
            .O(N__16945),
            .I(N__16942));
    Odrv4 I__2176 (
            .O(N__16942),
            .I(\POWERLED.mult1_un131_sum_axb_4_l_fx ));
    CascadeMux I__2175 (
            .O(N__16939),
            .I(N__16936));
    InMux I__2174 (
            .O(N__16936),
            .I(N__16932));
    InMux I__2173 (
            .O(N__16935),
            .I(N__16929));
    LocalMux I__2172 (
            .O(N__16932),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    LocalMux I__2171 (
            .O(N__16929),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__2170 (
            .O(N__16924),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    CascadeMux I__2169 (
            .O(N__16921),
            .I(N__16918));
    InMux I__2168 (
            .O(N__16918),
            .I(N__16915));
    LocalMux I__2167 (
            .O(N__16915),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__2166 (
            .O(N__16912),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__2165 (
            .O(N__16909),
            .I(N__16906));
    LocalMux I__2164 (
            .O(N__16906),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__2163 (
            .O(N__16903),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__2162 (
            .O(N__16900),
            .I(N__16897));
    LocalMux I__2161 (
            .O(N__16897),
            .I(N__16894));
    Odrv12 I__2160 (
            .O(N__16894),
            .I(\POWERLED.mult1_un131_sum_axb_7_l_fx ));
    CascadeMux I__2159 (
            .O(N__16891),
            .I(N__16888));
    InMux I__2158 (
            .O(N__16888),
            .I(N__16884));
    InMux I__2157 (
            .O(N__16887),
            .I(N__16881));
    LocalMux I__2156 (
            .O(N__16884),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    LocalMux I__2155 (
            .O(N__16881),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__2154 (
            .O(N__16876),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__2153 (
            .O(N__16873),
            .I(N__16870));
    LocalMux I__2152 (
            .O(N__16870),
            .I(N__16867));
    Span4Mux_v I__2151 (
            .O(N__16867),
            .I(N__16864));
    Odrv4 I__2150 (
            .O(N__16864),
            .I(\POWERLED.mult1_un110_sum_i ));
    CascadeMux I__2149 (
            .O(N__16861),
            .I(N__16858));
    InMux I__2148 (
            .O(N__16858),
            .I(N__16855));
    LocalMux I__2147 (
            .O(N__16855),
            .I(\POWERLED.mult1_un117_sum_i ));
    InMux I__2146 (
            .O(N__16852),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    InMux I__2145 (
            .O(N__16849),
            .I(N__16846));
    LocalMux I__2144 (
            .O(N__16846),
            .I(N__16843));
    Odrv4 I__2143 (
            .O(N__16843),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__2142 (
            .O(N__16840),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__2141 (
            .O(N__16837),
            .I(N__16834));
    LocalMux I__2140 (
            .O(N__16834),
            .I(N__16831));
    Odrv4 I__2139 (
            .O(N__16831),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__2138 (
            .O(N__16828),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    CascadeMux I__2137 (
            .O(N__16825),
            .I(N__16822));
    InMux I__2136 (
            .O(N__16822),
            .I(N__16819));
    LocalMux I__2135 (
            .O(N__16819),
            .I(N__16816));
    Odrv4 I__2134 (
            .O(N__16816),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__2133 (
            .O(N__16813),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    CascadeMux I__2132 (
            .O(N__16810),
            .I(N__16807));
    InMux I__2131 (
            .O(N__16807),
            .I(N__16804));
    LocalMux I__2130 (
            .O(N__16804),
            .I(N__16801));
    Odrv12 I__2129 (
            .O(N__16801),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__2128 (
            .O(N__16798),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    IoInMux I__2127 (
            .O(N__16795),
            .I(N__16792));
    LocalMux I__2126 (
            .O(N__16792),
            .I(N__16788));
    IoInMux I__2125 (
            .O(N__16791),
            .I(N__16785));
    Span4Mux_s3_h I__2124 (
            .O(N__16788),
            .I(N__16782));
    LocalMux I__2123 (
            .O(N__16785),
            .I(N__16779));
    Odrv4 I__2122 (
            .O(N__16782),
            .I(v5s_enn));
    Odrv12 I__2121 (
            .O(N__16779),
            .I(v5s_enn));
    CascadeMux I__2120 (
            .O(N__16774),
            .I(N__16771));
    InMux I__2119 (
            .O(N__16771),
            .I(N__16768));
    LocalMux I__2118 (
            .O(N__16768),
            .I(\POWERLED.mult1_un47_sum_i ));
    InMux I__2117 (
            .O(N__16765),
            .I(N__16762));
    LocalMux I__2116 (
            .O(N__16762),
            .I(N__16759));
    Span4Mux_v I__2115 (
            .O(N__16759),
            .I(N__16756));
    Odrv4 I__2114 (
            .O(N__16756),
            .I(\POWERLED.mult1_un103_sum_i ));
    IoInMux I__2113 (
            .O(N__16753),
            .I(N__16750));
    LocalMux I__2112 (
            .O(N__16750),
            .I(N__16747));
    Span4Mux_s3_h I__2111 (
            .O(N__16747),
            .I(N__16744));
    Odrv4 I__2110 (
            .O(N__16744),
            .I(v33a_enn));
    InMux I__2109 (
            .O(N__16741),
            .I(N__16738));
    LocalMux I__2108 (
            .O(N__16738),
            .I(N__16735));
    Span4Mux_s3_h I__2107 (
            .O(N__16735),
            .I(N__16732));
    Odrv4 I__2106 (
            .O(N__16732),
            .I(\POWERLED.un85_clk_100khz_6 ));
    CascadeMux I__2105 (
            .O(N__16729),
            .I(\POWERLED.un2_count_clk_17_0_a2_1_cascade_ ));
    CascadeMux I__2104 (
            .O(N__16726),
            .I(\POWERLED.un2_count_clk_17_0_a2_5_cascade_ ));
    InMux I__2103 (
            .O(N__16723),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__2102 (
            .O(N__16720),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__2101 (
            .O(N__16717),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__2100 (
            .O(N__16714),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__2099 (
            .O(N__16711),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__2098 (
            .O(N__16708),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    InMux I__2097 (
            .O(N__16705),
            .I(N__16702));
    LocalMux I__2096 (
            .O(N__16702),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    CascadeMux I__2095 (
            .O(N__16699),
            .I(\POWERLED.dutycycle_eena_3_1_cascade_ ));
    InMux I__2094 (
            .O(N__16696),
            .I(N__16693));
    LocalMux I__2093 (
            .O(N__16693),
            .I(\POWERLED.dutycycle_eena_3 ));
    InMux I__2092 (
            .O(N__16690),
            .I(N__16684));
    InMux I__2091 (
            .O(N__16689),
            .I(N__16684));
    LocalMux I__2090 (
            .O(N__16684),
            .I(N__16681));
    Odrv4 I__2089 (
            .O(N__16681),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    CascadeMux I__2088 (
            .O(N__16678),
            .I(\POWERLED.dutycycle_eena_3_cascade_ ));
    CascadeMux I__2087 (
            .O(N__16675),
            .I(\POWERLED.dutycycleZ0Z_2_cascade_ ));
    CascadeMux I__2086 (
            .O(N__16672),
            .I(\POWERLED.un1_dutycycle_53_4_0_cascade_ ));
    InMux I__2085 (
            .O(N__16669),
            .I(N__16666));
    LocalMux I__2084 (
            .O(N__16666),
            .I(\POWERLED.un1_dutycycle_53_4_3_1 ));
    CascadeMux I__2083 (
            .O(N__16663),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_12_cascade_ ));
    InMux I__2082 (
            .O(N__16660),
            .I(N__16657));
    LocalMux I__2081 (
            .O(N__16657),
            .I(\POWERLED.un1_dutycycle_53_8_3 ));
    CascadeMux I__2080 (
            .O(N__16654),
            .I(N__16650));
    InMux I__2079 (
            .O(N__16653),
            .I(N__16647));
    InMux I__2078 (
            .O(N__16650),
            .I(N__16644));
    LocalMux I__2077 (
            .O(N__16647),
            .I(N__16641));
    LocalMux I__2076 (
            .O(N__16644),
            .I(N__16636));
    Span4Mux_h I__2075 (
            .O(N__16641),
            .I(N__16633));
    InMux I__2074 (
            .O(N__16640),
            .I(N__16628));
    InMux I__2073 (
            .O(N__16639),
            .I(N__16628));
    Span12Mux_s3_h I__2072 (
            .O(N__16636),
            .I(N__16625));
    Odrv4 I__2071 (
            .O(N__16633),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3 ));
    LocalMux I__2070 (
            .O(N__16628),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3 ));
    Odrv12 I__2069 (
            .O(N__16625),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3 ));
    InMux I__2068 (
            .O(N__16618),
            .I(N__16615));
    LocalMux I__2067 (
            .O(N__16615),
            .I(\POWERLED.un1_dutycycle_53_56_a0_1 ));
    InMux I__2066 (
            .O(N__16612),
            .I(N__16609));
    LocalMux I__2065 (
            .O(N__16609),
            .I(\POWERLED.un1_dutycycle_53_56_a1_1 ));
    CascadeMux I__2064 (
            .O(N__16606),
            .I(\POWERLED.un1_clk_100khz_45_and_i_i_a3_0_0_cascade_ ));
    CascadeMux I__2063 (
            .O(N__16603),
            .I(\POWERLED.N_4_cascade_ ));
    CascadeMux I__2062 (
            .O(N__16600),
            .I(\POWERLED.un1_dutycycle_53_axb_7_cascade_ ));
    CascadeMux I__2061 (
            .O(N__16597),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3_cascade_ ));
    InMux I__2060 (
            .O(N__16594),
            .I(N__16591));
    LocalMux I__2059 (
            .O(N__16591),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_10 ));
    CascadeMux I__2058 (
            .O(N__16588),
            .I(\POWERLED.un1_dutycycle_53_axb_4_1_cascade_ ));
    InMux I__2057 (
            .O(N__16585),
            .I(N__16582));
    LocalMux I__2056 (
            .O(N__16582),
            .I(\POWERLED.un1_dutycycle_53_8_2_0 ));
    CascadeMux I__2055 (
            .O(N__16579),
            .I(\POWERLED.un1_dutycycle_53_8_2_cascade_ ));
    CascadeMux I__2054 (
            .O(N__16576),
            .I(\POWERLED.un1_dutycycle_53_8_5_cascade_ ));
    InMux I__2053 (
            .O(N__16573),
            .I(N__16570));
    LocalMux I__2052 (
            .O(N__16570),
            .I(\POWERLED.count_off_0_7 ));
    InMux I__2051 (
            .O(N__16567),
            .I(N__16563));
    InMux I__2050 (
            .O(N__16566),
            .I(N__16560));
    LocalMux I__2049 (
            .O(N__16563),
            .I(N__16557));
    LocalMux I__2048 (
            .O(N__16560),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    Odrv4 I__2047 (
            .O(N__16557),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    InMux I__2046 (
            .O(N__16552),
            .I(N__16548));
    InMux I__2045 (
            .O(N__16551),
            .I(N__16545));
    LocalMux I__2044 (
            .O(N__16548),
            .I(N__16542));
    LocalMux I__2043 (
            .O(N__16545),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    Odrv12 I__2042 (
            .O(N__16542),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    CascadeMux I__2041 (
            .O(N__16537),
            .I(N__16534));
    InMux I__2040 (
            .O(N__16534),
            .I(N__16531));
    LocalMux I__2039 (
            .O(N__16531),
            .I(N__16527));
    InMux I__2038 (
            .O(N__16530),
            .I(N__16524));
    Span4Mux_v I__2037 (
            .O(N__16527),
            .I(N__16521));
    LocalMux I__2036 (
            .O(N__16524),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    Odrv4 I__2035 (
            .O(N__16521),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    InMux I__2034 (
            .O(N__16516),
            .I(N__16512));
    InMux I__2033 (
            .O(N__16515),
            .I(N__16509));
    LocalMux I__2032 (
            .O(N__16512),
            .I(N__16506));
    LocalMux I__2031 (
            .O(N__16509),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    Odrv4 I__2030 (
            .O(N__16506),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    InMux I__2029 (
            .O(N__16501),
            .I(N__16498));
    LocalMux I__2028 (
            .O(N__16498),
            .I(N__16495));
    Odrv4 I__2027 (
            .O(N__16495),
            .I(\DSW_PWRGD.un4_count_8 ));
    CascadeMux I__2026 (
            .O(N__16492),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_3_cascade_ ));
    InMux I__2025 (
            .O(N__16489),
            .I(N__16486));
    LocalMux I__2024 (
            .O(N__16486),
            .I(N__16483));
    Span4Mux_h I__2023 (
            .O(N__16483),
            .I(N__16479));
    InMux I__2022 (
            .O(N__16482),
            .I(N__16476));
    Odrv4 I__2021 (
            .O(N__16479),
            .I(\POWERLED.un1_dutycycle_53_20_0_0 ));
    LocalMux I__2020 (
            .O(N__16476),
            .I(\POWERLED.un1_dutycycle_53_20_0_0 ));
    CascadeMux I__2019 (
            .O(N__16471),
            .I(\POWERLED.o2_cascade_ ));
    CascadeMux I__2018 (
            .O(N__16468),
            .I(N__16465));
    InMux I__2017 (
            .O(N__16465),
            .I(N__16462));
    LocalMux I__2016 (
            .O(N__16462),
            .I(\POWERLED.un1_dutycycle_53_axb_7_1 ));
    InMux I__2015 (
            .O(N__16459),
            .I(N__16456));
    LocalMux I__2014 (
            .O(N__16456),
            .I(\POWERLED.count_off_0_4 ));
    InMux I__2013 (
            .O(N__16453),
            .I(N__16450));
    LocalMux I__2012 (
            .O(N__16450),
            .I(N__16447));
    Odrv4 I__2011 (
            .O(N__16447),
            .I(\POWERLED.count_off_0_8 ));
    CascadeMux I__2010 (
            .O(N__16444),
            .I(\POWERLED.count_offZ0Z_8_cascade_ ));
    CascadeMux I__2009 (
            .O(N__16441),
            .I(N__16438));
    InMux I__2008 (
            .O(N__16438),
            .I(N__16435));
    LocalMux I__2007 (
            .O(N__16435),
            .I(\POWERLED.count_off_0_3 ));
    InMux I__2006 (
            .O(N__16432),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__2005 (
            .O(N__16429),
            .I(N__16425));
    InMux I__2004 (
            .O(N__16428),
            .I(N__16420));
    InMux I__2003 (
            .O(N__16425),
            .I(N__16415));
    InMux I__2002 (
            .O(N__16424),
            .I(N__16415));
    InMux I__2001 (
            .O(N__16423),
            .I(N__16412));
    LocalMux I__2000 (
            .O(N__16420),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__1999 (
            .O(N__16415),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__1998 (
            .O(N__16412),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    CascadeMux I__1997 (
            .O(N__16405),
            .I(\POWERLED.mult1_un96_sum_s_8_cascade_ ));
    CascadeMux I__1996 (
            .O(N__16402),
            .I(N__16398));
    InMux I__1995 (
            .O(N__16401),
            .I(N__16390));
    InMux I__1994 (
            .O(N__16398),
            .I(N__16390));
    InMux I__1993 (
            .O(N__16397),
            .I(N__16390));
    LocalMux I__1992 (
            .O(N__16390),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__1991 (
            .O(N__16387),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    CascadeMux I__1990 (
            .O(N__16384),
            .I(N__16380));
    CascadeMux I__1989 (
            .O(N__16383),
            .I(N__16377));
    InMux I__1988 (
            .O(N__16380),
            .I(N__16372));
    InMux I__1987 (
            .O(N__16377),
            .I(N__16369));
    InMux I__1986 (
            .O(N__16376),
            .I(N__16366));
    InMux I__1985 (
            .O(N__16375),
            .I(N__16363));
    LocalMux I__1984 (
            .O(N__16372),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1983 (
            .O(N__16369),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1982 (
            .O(N__16366),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__1981 (
            .O(N__16363),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__1980 (
            .O(N__16354),
            .I(\POWERLED.mult1_un103_sum_s_8_cascade_ ));
    CascadeMux I__1979 (
            .O(N__16351),
            .I(N__16347));
    CascadeMux I__1978 (
            .O(N__16350),
            .I(N__16343));
    InMux I__1977 (
            .O(N__16347),
            .I(N__16336));
    InMux I__1976 (
            .O(N__16346),
            .I(N__16336));
    InMux I__1975 (
            .O(N__16343),
            .I(N__16336));
    LocalMux I__1974 (
            .O(N__16336),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    InMux I__1973 (
            .O(N__16333),
            .I(N__16330));
    LocalMux I__1972 (
            .O(N__16330),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__1971 (
            .O(N__16327),
            .I(\POWERLED.mult1_un96_sum_cry_2_c ));
    CascadeMux I__1970 (
            .O(N__16324),
            .I(N__16321));
    InMux I__1969 (
            .O(N__16321),
            .I(N__16318));
    LocalMux I__1968 (
            .O(N__16318),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__1967 (
            .O(N__16315),
            .I(\POWERLED.mult1_un96_sum_cry_3_c ));
    InMux I__1966 (
            .O(N__16312),
            .I(N__16309));
    LocalMux I__1965 (
            .O(N__16309),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__1964 (
            .O(N__16306),
            .I(\POWERLED.mult1_un96_sum_cry_4_c ));
    CascadeMux I__1963 (
            .O(N__16303),
            .I(N__16300));
    InMux I__1962 (
            .O(N__16300),
            .I(N__16297));
    LocalMux I__1961 (
            .O(N__16297),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    InMux I__1960 (
            .O(N__16294),
            .I(\POWERLED.mult1_un96_sum_cry_5_c ));
    CascadeMux I__1959 (
            .O(N__16291),
            .I(N__16288));
    InMux I__1958 (
            .O(N__16288),
            .I(N__16279));
    InMux I__1957 (
            .O(N__16287),
            .I(N__16279));
    InMux I__1956 (
            .O(N__16286),
            .I(N__16279));
    LocalMux I__1955 (
            .O(N__16279),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__1954 (
            .O(N__16276),
            .I(N__16273));
    LocalMux I__1953 (
            .O(N__16273),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__1952 (
            .O(N__16270),
            .I(\POWERLED.mult1_un96_sum_cry_6_c ));
    InMux I__1951 (
            .O(N__16267),
            .I(N__16264));
    LocalMux I__1950 (
            .O(N__16264),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__1949 (
            .O(N__16261),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__1948 (
            .O(N__16258),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    InMux I__1947 (
            .O(N__16255),
            .I(N__16250));
    CascadeMux I__1946 (
            .O(N__16254),
            .I(N__16247));
    CascadeMux I__1945 (
            .O(N__16253),
            .I(N__16244));
    LocalMux I__1944 (
            .O(N__16250),
            .I(N__16239));
    InMux I__1943 (
            .O(N__16247),
            .I(N__16236));
    InMux I__1942 (
            .O(N__16244),
            .I(N__16233));
    InMux I__1941 (
            .O(N__16243),
            .I(N__16230));
    InMux I__1940 (
            .O(N__16242),
            .I(N__16227));
    Odrv4 I__1939 (
            .O(N__16239),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1938 (
            .O(N__16236),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1937 (
            .O(N__16233),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1936 (
            .O(N__16230),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__1935 (
            .O(N__16227),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__1934 (
            .O(N__16216),
            .I(N__16211));
    CascadeMux I__1933 (
            .O(N__16215),
            .I(N__16208));
    CascadeMux I__1932 (
            .O(N__16214),
            .I(N__16205));
    InMux I__1931 (
            .O(N__16211),
            .I(N__16202));
    InMux I__1930 (
            .O(N__16208),
            .I(N__16197));
    InMux I__1929 (
            .O(N__16205),
            .I(N__16197));
    LocalMux I__1928 (
            .O(N__16202),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    LocalMux I__1927 (
            .O(N__16197),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    CascadeMux I__1926 (
            .O(N__16192),
            .I(N__16189));
    InMux I__1925 (
            .O(N__16189),
            .I(N__16186));
    LocalMux I__1924 (
            .O(N__16186),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__1923 (
            .O(N__16183),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    InMux I__1922 (
            .O(N__16180),
            .I(N__16177));
    LocalMux I__1921 (
            .O(N__16177),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__1920 (
            .O(N__16174),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__1919 (
            .O(N__16171),
            .I(N__16168));
    LocalMux I__1918 (
            .O(N__16168),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__1917 (
            .O(N__16165),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    InMux I__1916 (
            .O(N__16162),
            .I(N__16159));
    LocalMux I__1915 (
            .O(N__16159),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__1914 (
            .O(N__16156),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__1913 (
            .O(N__16153),
            .I(N__16150));
    LocalMux I__1912 (
            .O(N__16150),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__1911 (
            .O(N__16147),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    InMux I__1910 (
            .O(N__16144),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__1909 (
            .O(N__16141),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__1908 (
            .O(N__16138),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__1907 (
            .O(N__16135),
            .I(\POWERLED.mult1_un117_sum_s_8_cascade_ ));
    InMux I__1906 (
            .O(N__16132),
            .I(N__16129));
    LocalMux I__1905 (
            .O(N__16129),
            .I(\POWERLED.un85_clk_100khz_7 ));
    InMux I__1904 (
            .O(N__16126),
            .I(N__16123));
    LocalMux I__1903 (
            .O(N__16123),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__1902 (
            .O(N__16120),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    InMux I__1901 (
            .O(N__16117),
            .I(N__16114));
    LocalMux I__1900 (
            .O(N__16114),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__1899 (
            .O(N__16111),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    InMux I__1898 (
            .O(N__16108),
            .I(N__16105));
    LocalMux I__1897 (
            .O(N__16105),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__1896 (
            .O(N__16102),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__1895 (
            .O(N__16099),
            .I(N__16096));
    LocalMux I__1894 (
            .O(N__16096),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__1893 (
            .O(N__16093),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    CascadeMux I__1892 (
            .O(N__16090),
            .I(N__16087));
    InMux I__1891 (
            .O(N__16087),
            .I(N__16081));
    InMux I__1890 (
            .O(N__16086),
            .I(N__16081));
    LocalMux I__1889 (
            .O(N__16081),
            .I(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ));
    InMux I__1888 (
            .O(N__16078),
            .I(N__16075));
    LocalMux I__1887 (
            .O(N__16075),
            .I(\POWERLED.count_0_15 ));
    InMux I__1886 (
            .O(N__16072),
            .I(N__16068));
    InMux I__1885 (
            .O(N__16071),
            .I(N__16064));
    LocalMux I__1884 (
            .O(N__16068),
            .I(N__16061));
    InMux I__1883 (
            .O(N__16067),
            .I(N__16058));
    LocalMux I__1882 (
            .O(N__16064),
            .I(\POWERLED.countZ0Z_7 ));
    Odrv4 I__1881 (
            .O(N__16061),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__1880 (
            .O(N__16058),
            .I(\POWERLED.countZ0Z_7 ));
    CascadeMux I__1879 (
            .O(N__16051),
            .I(N__16048));
    InMux I__1878 (
            .O(N__16048),
            .I(N__16042));
    InMux I__1877 (
            .O(N__16047),
            .I(N__16042));
    LocalMux I__1876 (
            .O(N__16042),
            .I(N__16039));
    Odrv4 I__1875 (
            .O(N__16039),
            .I(\POWERLED.count_1_7 ));
    InMux I__1874 (
            .O(N__16036),
            .I(N__16033));
    LocalMux I__1873 (
            .O(N__16033),
            .I(\POWERLED.count_0_7 ));
    InMux I__1872 (
            .O(N__16030),
            .I(N__16027));
    LocalMux I__1871 (
            .O(N__16027),
            .I(N__16023));
    InMux I__1870 (
            .O(N__16026),
            .I(N__16020));
    Span4Mux_s3_v I__1869 (
            .O(N__16023),
            .I(N__16014));
    LocalMux I__1868 (
            .O(N__16020),
            .I(N__16014));
    InMux I__1867 (
            .O(N__16019),
            .I(N__16011));
    Odrv4 I__1866 (
            .O(N__16014),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__1865 (
            .O(N__16011),
            .I(\POWERLED.countZ0Z_8 ));
    CascadeMux I__1864 (
            .O(N__16006),
            .I(N__16002));
    InMux I__1863 (
            .O(N__16005),
            .I(N__15997));
    InMux I__1862 (
            .O(N__16002),
            .I(N__15997));
    LocalMux I__1861 (
            .O(N__15997),
            .I(N__15994));
    Odrv4 I__1860 (
            .O(N__15994),
            .I(\POWERLED.count_1_8 ));
    InMux I__1859 (
            .O(N__15991),
            .I(N__15988));
    LocalMux I__1858 (
            .O(N__15988),
            .I(\POWERLED.count_0_8 ));
    InMux I__1857 (
            .O(N__15985),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__1856 (
            .O(N__15982),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__1855 (
            .O(N__15979),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__1854 (
            .O(N__15976),
            .I(N__15971));
    InMux I__1853 (
            .O(N__15975),
            .I(N__15968));
    InMux I__1852 (
            .O(N__15974),
            .I(N__15965));
    LocalMux I__1851 (
            .O(N__15971),
            .I(N__15960));
    LocalMux I__1850 (
            .O(N__15968),
            .I(N__15960));
    LocalMux I__1849 (
            .O(N__15965),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv12 I__1848 (
            .O(N__15960),
            .I(\POWERLED.countZ0Z_12 ));
    InMux I__1847 (
            .O(N__15955),
            .I(N__15949));
    InMux I__1846 (
            .O(N__15954),
            .I(N__15949));
    LocalMux I__1845 (
            .O(N__15949),
            .I(\POWERLED.count_1_12 ));
    InMux I__1844 (
            .O(N__15946),
            .I(\POWERLED.un1_count_cry_11_cZ0 ));
    InMux I__1843 (
            .O(N__15943),
            .I(N__15938));
    CascadeMux I__1842 (
            .O(N__15942),
            .I(N__15935));
    InMux I__1841 (
            .O(N__15941),
            .I(N__15932));
    LocalMux I__1840 (
            .O(N__15938),
            .I(N__15929));
    InMux I__1839 (
            .O(N__15935),
            .I(N__15926));
    LocalMux I__1838 (
            .O(N__15932),
            .I(N__15923));
    Sp12to4 I__1837 (
            .O(N__15929),
            .I(N__15918));
    LocalMux I__1836 (
            .O(N__15926),
            .I(N__15918));
    Odrv4 I__1835 (
            .O(N__15923),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv12 I__1834 (
            .O(N__15918),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__1833 (
            .O(N__15913),
            .I(N__15907));
    InMux I__1832 (
            .O(N__15912),
            .I(N__15907));
    LocalMux I__1831 (
            .O(N__15907),
            .I(N__15904));
    Odrv4 I__1830 (
            .O(N__15904),
            .I(\POWERLED.count_1_13 ));
    InMux I__1829 (
            .O(N__15901),
            .I(\POWERLED.un1_count_cry_12 ));
    InMux I__1828 (
            .O(N__15898),
            .I(N__15894));
    InMux I__1827 (
            .O(N__15897),
            .I(N__15890));
    LocalMux I__1826 (
            .O(N__15894),
            .I(N__15887));
    InMux I__1825 (
            .O(N__15893),
            .I(N__15884));
    LocalMux I__1824 (
            .O(N__15890),
            .I(N__15881));
    Span4Mux_v I__1823 (
            .O(N__15887),
            .I(N__15876));
    LocalMux I__1822 (
            .O(N__15884),
            .I(N__15876));
    Odrv4 I__1821 (
            .O(N__15881),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__1820 (
            .O(N__15876),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__1819 (
            .O(N__15871),
            .I(N__15865));
    InMux I__1818 (
            .O(N__15870),
            .I(N__15865));
    LocalMux I__1817 (
            .O(N__15865),
            .I(N__15862));
    Odrv4 I__1816 (
            .O(N__15862),
            .I(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ));
    InMux I__1815 (
            .O(N__15859),
            .I(\POWERLED.un1_count_cry_13_cZ0 ));
    CascadeMux I__1814 (
            .O(N__15856),
            .I(N__15852));
    InMux I__1813 (
            .O(N__15855),
            .I(N__15830));
    InMux I__1812 (
            .O(N__15852),
            .I(N__15830));
    InMux I__1811 (
            .O(N__15851),
            .I(N__15830));
    InMux I__1810 (
            .O(N__15850),
            .I(N__15821));
    InMux I__1809 (
            .O(N__15849),
            .I(N__15821));
    InMux I__1808 (
            .O(N__15848),
            .I(N__15821));
    InMux I__1807 (
            .O(N__15847),
            .I(N__15821));
    InMux I__1806 (
            .O(N__15846),
            .I(N__15814));
    InMux I__1805 (
            .O(N__15845),
            .I(N__15814));
    InMux I__1804 (
            .O(N__15844),
            .I(N__15814));
    InMux I__1803 (
            .O(N__15843),
            .I(N__15807));
    InMux I__1802 (
            .O(N__15842),
            .I(N__15807));
    InMux I__1801 (
            .O(N__15841),
            .I(N__15807));
    InMux I__1800 (
            .O(N__15840),
            .I(N__15798));
    InMux I__1799 (
            .O(N__15839),
            .I(N__15798));
    InMux I__1798 (
            .O(N__15838),
            .I(N__15798));
    InMux I__1797 (
            .O(N__15837),
            .I(N__15798));
    LocalMux I__1796 (
            .O(N__15830),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__1795 (
            .O(N__15821),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__1794 (
            .O(N__15814),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__1793 (
            .O(N__15807),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__1792 (
            .O(N__15798),
            .I(\POWERLED.count_0_sqmuxa_i ));
    InMux I__1791 (
            .O(N__15787),
            .I(\POWERLED.un1_count_cry_14 ));
    InMux I__1790 (
            .O(N__15784),
            .I(N__15781));
    LocalMux I__1789 (
            .O(N__15781),
            .I(N__15778));
    Span4Mux_v I__1788 (
            .O(N__15778),
            .I(N__15775));
    Odrv4 I__1787 (
            .O(N__15775),
            .I(\POWERLED.count_0_9 ));
    InMux I__1786 (
            .O(N__15772),
            .I(N__15769));
    LocalMux I__1785 (
            .O(N__15769),
            .I(N__15765));
    InMux I__1784 (
            .O(N__15768),
            .I(N__15762));
    Odrv4 I__1783 (
            .O(N__15765),
            .I(\POWERLED.count_1_9 ));
    LocalMux I__1782 (
            .O(N__15762),
            .I(\POWERLED.count_1_9 ));
    InMux I__1781 (
            .O(N__15757),
            .I(N__15754));
    LocalMux I__1780 (
            .O(N__15754),
            .I(N__15749));
    InMux I__1779 (
            .O(N__15753),
            .I(N__15746));
    InMux I__1778 (
            .O(N__15752),
            .I(N__15743));
    Odrv4 I__1777 (
            .O(N__15749),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__1776 (
            .O(N__15746),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__1775 (
            .O(N__15743),
            .I(\POWERLED.countZ0Z_9 ));
    InMux I__1774 (
            .O(N__15736),
            .I(N__15732));
    InMux I__1773 (
            .O(N__15735),
            .I(N__15728));
    LocalMux I__1772 (
            .O(N__15732),
            .I(N__15725));
    InMux I__1771 (
            .O(N__15731),
            .I(N__15722));
    LocalMux I__1770 (
            .O(N__15728),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__1769 (
            .O(N__15725),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__1768 (
            .O(N__15722),
            .I(\POWERLED.countZ0Z_6 ));
    CascadeMux I__1767 (
            .O(N__15715),
            .I(N__15712));
    InMux I__1766 (
            .O(N__15712),
            .I(N__15706));
    InMux I__1765 (
            .O(N__15711),
            .I(N__15706));
    LocalMux I__1764 (
            .O(N__15706),
            .I(N__15703));
    Odrv4 I__1763 (
            .O(N__15703),
            .I(\POWERLED.count_1_6 ));
    InMux I__1762 (
            .O(N__15700),
            .I(N__15697));
    LocalMux I__1761 (
            .O(N__15697),
            .I(\POWERLED.count_0_6 ));
    InMux I__1760 (
            .O(N__15694),
            .I(N__15691));
    LocalMux I__1759 (
            .O(N__15691),
            .I(N__15688));
    Span12Mux_s1_h I__1758 (
            .O(N__15688),
            .I(N__15683));
    InMux I__1757 (
            .O(N__15687),
            .I(N__15680));
    InMux I__1756 (
            .O(N__15686),
            .I(N__15677));
    Odrv12 I__1755 (
            .O(N__15683),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__1754 (
            .O(N__15680),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__1753 (
            .O(N__15677),
            .I(\POWERLED.countZ0Z_15 ));
    InMux I__1752 (
            .O(N__15670),
            .I(N__15665));
    InMux I__1751 (
            .O(N__15669),
            .I(N__15662));
    InMux I__1750 (
            .O(N__15668),
            .I(N__15659));
    LocalMux I__1749 (
            .O(N__15665),
            .I(N__15654));
    LocalMux I__1748 (
            .O(N__15662),
            .I(N__15654));
    LocalMux I__1747 (
            .O(N__15659),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv12 I__1746 (
            .O(N__15654),
            .I(\POWERLED.countZ0Z_4 ));
    CascadeMux I__1745 (
            .O(N__15649),
            .I(N__15646));
    InMux I__1744 (
            .O(N__15646),
            .I(N__15640));
    InMux I__1743 (
            .O(N__15645),
            .I(N__15640));
    LocalMux I__1742 (
            .O(N__15640),
            .I(\POWERLED.count_1_4 ));
    InMux I__1741 (
            .O(N__15637),
            .I(\POWERLED.un1_count_cry_3 ));
    InMux I__1740 (
            .O(N__15634),
            .I(N__15631));
    LocalMux I__1739 (
            .O(N__15631),
            .I(N__15626));
    InMux I__1738 (
            .O(N__15630),
            .I(N__15623));
    InMux I__1737 (
            .O(N__15629),
            .I(N__15620));
    Span4Mux_v I__1736 (
            .O(N__15626),
            .I(N__15615));
    LocalMux I__1735 (
            .O(N__15623),
            .I(N__15615));
    LocalMux I__1734 (
            .O(N__15620),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__1733 (
            .O(N__15615),
            .I(\POWERLED.countZ0Z_5 ));
    CascadeMux I__1732 (
            .O(N__15610),
            .I(N__15607));
    InMux I__1731 (
            .O(N__15607),
            .I(N__15601));
    InMux I__1730 (
            .O(N__15606),
            .I(N__15601));
    LocalMux I__1729 (
            .O(N__15601),
            .I(\POWERLED.count_1_5 ));
    InMux I__1728 (
            .O(N__15598),
            .I(\POWERLED.un1_count_cry_4 ));
    InMux I__1727 (
            .O(N__15595),
            .I(\POWERLED.un1_count_cry_5 ));
    InMux I__1726 (
            .O(N__15592),
            .I(\POWERLED.un1_count_cry_6 ));
    InMux I__1725 (
            .O(N__15589),
            .I(\POWERLED.un1_count_cry_7 ));
    InMux I__1724 (
            .O(N__15586),
            .I(bfn_2_11_0_));
    InMux I__1723 (
            .O(N__15583),
            .I(N__15580));
    LocalMux I__1722 (
            .O(N__15580),
            .I(N__15575));
    InMux I__1721 (
            .O(N__15579),
            .I(N__15572));
    InMux I__1720 (
            .O(N__15578),
            .I(N__15569));
    Span4Mux_v I__1719 (
            .O(N__15575),
            .I(N__15562));
    LocalMux I__1718 (
            .O(N__15572),
            .I(N__15562));
    LocalMux I__1717 (
            .O(N__15569),
            .I(N__15562));
    Odrv4 I__1716 (
            .O(N__15562),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__1715 (
            .O(N__15559),
            .I(N__15553));
    InMux I__1714 (
            .O(N__15558),
            .I(N__15553));
    LocalMux I__1713 (
            .O(N__15553),
            .I(N__15550));
    Odrv4 I__1712 (
            .O(N__15550),
            .I(\POWERLED.count_1_10 ));
    InMux I__1711 (
            .O(N__15547),
            .I(\POWERLED.un1_count_cry_9 ));
    InMux I__1710 (
            .O(N__15544),
            .I(N__15540));
    InMux I__1709 (
            .O(N__15543),
            .I(N__15537));
    LocalMux I__1708 (
            .O(N__15540),
            .I(N__15533));
    LocalMux I__1707 (
            .O(N__15537),
            .I(N__15530));
    InMux I__1706 (
            .O(N__15536),
            .I(N__15527));
    Span4Mux_v I__1705 (
            .O(N__15533),
            .I(N__15520));
    Span4Mux_v I__1704 (
            .O(N__15530),
            .I(N__15520));
    LocalMux I__1703 (
            .O(N__15527),
            .I(N__15520));
    Odrv4 I__1702 (
            .O(N__15520),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__1701 (
            .O(N__15517),
            .I(N__15511));
    InMux I__1700 (
            .O(N__15516),
            .I(N__15511));
    LocalMux I__1699 (
            .O(N__15511),
            .I(N__15508));
    Odrv4 I__1698 (
            .O(N__15508),
            .I(\POWERLED.count_1_11 ));
    InMux I__1697 (
            .O(N__15505),
            .I(\POWERLED.un1_count_cry_10 ));
    InMux I__1696 (
            .O(N__15502),
            .I(N__15499));
    LocalMux I__1695 (
            .O(N__15499),
            .I(\POWERLED.count_0_10 ));
    InMux I__1694 (
            .O(N__15496),
            .I(N__15493));
    LocalMux I__1693 (
            .O(N__15493),
            .I(\POWERLED.count_0_2 ));
    InMux I__1692 (
            .O(N__15490),
            .I(N__15487));
    LocalMux I__1691 (
            .O(N__15487),
            .I(\POWERLED.count_0_11 ));
    InMux I__1690 (
            .O(N__15484),
            .I(N__15481));
    LocalMux I__1689 (
            .O(N__15481),
            .I(N__15476));
    InMux I__1688 (
            .O(N__15480),
            .I(N__15473));
    InMux I__1687 (
            .O(N__15479),
            .I(N__15470));
    Odrv12 I__1686 (
            .O(N__15476),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__1685 (
            .O(N__15473),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__1684 (
            .O(N__15470),
            .I(\POWERLED.countZ0Z_1 ));
    InMux I__1683 (
            .O(N__15463),
            .I(N__15459));
    CascadeMux I__1682 (
            .O(N__15462),
            .I(N__15452));
    LocalMux I__1681 (
            .O(N__15459),
            .I(N__15449));
    InMux I__1680 (
            .O(N__15458),
            .I(N__15446));
    InMux I__1679 (
            .O(N__15457),
            .I(N__15439));
    InMux I__1678 (
            .O(N__15456),
            .I(N__15439));
    InMux I__1677 (
            .O(N__15455),
            .I(N__15439));
    InMux I__1676 (
            .O(N__15452),
            .I(N__15436));
    Odrv4 I__1675 (
            .O(N__15449),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__1674 (
            .O(N__15446),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__1673 (
            .O(N__15439),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__1672 (
            .O(N__15436),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__1671 (
            .O(N__15427),
            .I(N__15424));
    LocalMux I__1670 (
            .O(N__15424),
            .I(N__15419));
    InMux I__1669 (
            .O(N__15423),
            .I(N__15416));
    InMux I__1668 (
            .O(N__15422),
            .I(N__15413));
    Span4Mux_v I__1667 (
            .O(N__15419),
            .I(N__15408));
    LocalMux I__1666 (
            .O(N__15416),
            .I(N__15408));
    LocalMux I__1665 (
            .O(N__15413),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__1664 (
            .O(N__15408),
            .I(\POWERLED.countZ0Z_2 ));
    CascadeMux I__1663 (
            .O(N__15403),
            .I(N__15399));
    InMux I__1662 (
            .O(N__15402),
            .I(N__15394));
    InMux I__1661 (
            .O(N__15399),
            .I(N__15394));
    LocalMux I__1660 (
            .O(N__15394),
            .I(\POWERLED.count_1_2 ));
    InMux I__1659 (
            .O(N__15391),
            .I(\POWERLED.un1_count_cry_1 ));
    CascadeMux I__1658 (
            .O(N__15388),
            .I(N__15384));
    InMux I__1657 (
            .O(N__15387),
            .I(N__15380));
    InMux I__1656 (
            .O(N__15384),
            .I(N__15377));
    InMux I__1655 (
            .O(N__15383),
            .I(N__15374));
    LocalMux I__1654 (
            .O(N__15380),
            .I(N__15369));
    LocalMux I__1653 (
            .O(N__15377),
            .I(N__15369));
    LocalMux I__1652 (
            .O(N__15374),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__1651 (
            .O(N__15369),
            .I(\POWERLED.countZ0Z_3 ));
    CascadeMux I__1650 (
            .O(N__15364),
            .I(N__15361));
    InMux I__1649 (
            .O(N__15361),
            .I(N__15355));
    InMux I__1648 (
            .O(N__15360),
            .I(N__15355));
    LocalMux I__1647 (
            .O(N__15355),
            .I(\POWERLED.count_1_3 ));
    InMux I__1646 (
            .O(N__15352),
            .I(\POWERLED.un1_count_cry_2 ));
    CascadeMux I__1645 (
            .O(N__15349),
            .I(\POWERLED.dutycycle_RNIZ0Z_1_cascade_ ));
    CascadeMux I__1644 (
            .O(N__15346),
            .I(N__15343));
    InMux I__1643 (
            .O(N__15343),
            .I(N__15340));
    LocalMux I__1642 (
            .O(N__15340),
            .I(\POWERLED.un1_dutycycle_53_axb_3_1 ));
    CascadeMux I__1641 (
            .O(N__15337),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_9_cascade_ ));
    CascadeMux I__1640 (
            .O(N__15334),
            .I(DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_));
    SRMux I__1639 (
            .O(N__15331),
            .I(N__15327));
    SRMux I__1638 (
            .O(N__15330),
            .I(N__15323));
    LocalMux I__1637 (
            .O(N__15327),
            .I(N__15320));
    SRMux I__1636 (
            .O(N__15326),
            .I(N__15317));
    LocalMux I__1635 (
            .O(N__15323),
            .I(N__15314));
    Span4Mux_v I__1634 (
            .O(N__15320),
            .I(N__15311));
    LocalMux I__1633 (
            .O(N__15317),
            .I(N__15308));
    Span4Mux_s2_h I__1632 (
            .O(N__15314),
            .I(N__15305));
    Span4Mux_s1_h I__1631 (
            .O(N__15311),
            .I(N__15300));
    Span4Mux_s1_h I__1630 (
            .O(N__15308),
            .I(N__15300));
    Odrv4 I__1629 (
            .O(N__15305),
            .I(G_27));
    Odrv4 I__1628 (
            .O(N__15300),
            .I(G_27));
    CascadeMux I__1627 (
            .O(N__15295),
            .I(G_27_cascade_));
    CEMux I__1626 (
            .O(N__15292),
            .I(N__15289));
    LocalMux I__1625 (
            .O(N__15289),
            .I(N__15286));
    Odrv4 I__1624 (
            .O(N__15286),
            .I(\DSW_PWRGD.N_29_1 ));
    CascadeMux I__1623 (
            .O(N__15283),
            .I(\POWERLED.d_i1_mux_cascade_ ));
    CascadeMux I__1622 (
            .O(N__15280),
            .I(\POWERLED.dutycycle_RNI_16Z0Z_9_cascade_ ));
    CascadeMux I__1621 (
            .O(N__15277),
            .I(\POWERLED.d_i3_mux_cascade_ ));
    InMux I__1620 (
            .O(N__15274),
            .I(N__15268));
    InMux I__1619 (
            .O(N__15273),
            .I(N__15268));
    LocalMux I__1618 (
            .O(N__15268),
            .I(\POWERLED.un1_i3_mux ));
    InMux I__1617 (
            .O(N__15265),
            .I(N__15261));
    InMux I__1616 (
            .O(N__15264),
            .I(N__15258));
    LocalMux I__1615 (
            .O(N__15261),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    LocalMux I__1614 (
            .O(N__15258),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    InMux I__1613 (
            .O(N__15253),
            .I(N__15249));
    InMux I__1612 (
            .O(N__15252),
            .I(N__15246));
    LocalMux I__1611 (
            .O(N__15249),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    LocalMux I__1610 (
            .O(N__15246),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    CascadeMux I__1609 (
            .O(N__15241),
            .I(N__15237));
    InMux I__1608 (
            .O(N__15240),
            .I(N__15234));
    InMux I__1607 (
            .O(N__15237),
            .I(N__15231));
    LocalMux I__1606 (
            .O(N__15234),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    LocalMux I__1605 (
            .O(N__15231),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    InMux I__1604 (
            .O(N__15226),
            .I(N__15222));
    InMux I__1603 (
            .O(N__15225),
            .I(N__15219));
    LocalMux I__1602 (
            .O(N__15222),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    LocalMux I__1601 (
            .O(N__15219),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    InMux I__1600 (
            .O(N__15214),
            .I(N__15211));
    LocalMux I__1599 (
            .O(N__15211),
            .I(\DSW_PWRGD.un4_count_10 ));
    InMux I__1598 (
            .O(N__15208),
            .I(N__15204));
    InMux I__1597 (
            .O(N__15207),
            .I(N__15201));
    LocalMux I__1596 (
            .O(N__15204),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    LocalMux I__1595 (
            .O(N__15201),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    InMux I__1594 (
            .O(N__15196),
            .I(N__15192));
    InMux I__1593 (
            .O(N__15195),
            .I(N__15189));
    LocalMux I__1592 (
            .O(N__15192),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    LocalMux I__1591 (
            .O(N__15189),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    CascadeMux I__1590 (
            .O(N__15184),
            .I(N__15180));
    InMux I__1589 (
            .O(N__15183),
            .I(N__15177));
    InMux I__1588 (
            .O(N__15180),
            .I(N__15174));
    LocalMux I__1587 (
            .O(N__15177),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    LocalMux I__1586 (
            .O(N__15174),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    InMux I__1585 (
            .O(N__15169),
            .I(N__15165));
    InMux I__1584 (
            .O(N__15168),
            .I(N__15162));
    LocalMux I__1583 (
            .O(N__15165),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    LocalMux I__1582 (
            .O(N__15162),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    InMux I__1581 (
            .O(N__15157),
            .I(N__15154));
    LocalMux I__1580 (
            .O(N__15154),
            .I(\DSW_PWRGD.un4_count_11 ));
    CascadeMux I__1579 (
            .O(N__15151),
            .I(N__15147));
    InMux I__1578 (
            .O(N__15150),
            .I(N__15144));
    InMux I__1577 (
            .O(N__15147),
            .I(N__15141));
    LocalMux I__1576 (
            .O(N__15144),
            .I(\DSW_PWRGD.un1_curr_state10_0 ));
    LocalMux I__1575 (
            .O(N__15141),
            .I(\DSW_PWRGD.un1_curr_state10_0 ));
    InMux I__1574 (
            .O(N__15136),
            .I(N__15121));
    InMux I__1573 (
            .O(N__15135),
            .I(N__15121));
    InMux I__1572 (
            .O(N__15134),
            .I(N__15121));
    InMux I__1571 (
            .O(N__15133),
            .I(N__15121));
    InMux I__1570 (
            .O(N__15132),
            .I(N__15121));
    LocalMux I__1569 (
            .O(N__15121),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__1568 (
            .O(N__15118),
            .I(N__15113));
    InMux I__1567 (
            .O(N__15117),
            .I(N__15100));
    InMux I__1566 (
            .O(N__15116),
            .I(N__15100));
    InMux I__1565 (
            .O(N__15113),
            .I(N__15100));
    InMux I__1564 (
            .O(N__15112),
            .I(N__15100));
    InMux I__1563 (
            .O(N__15111),
            .I(N__15100));
    LocalMux I__1562 (
            .O(N__15100),
            .I(N__15097));
    Span4Mux_v I__1561 (
            .O(N__15097),
            .I(N__15094));
    Span4Mux_v I__1560 (
            .O(N__15094),
            .I(N__15091));
    Odrv4 I__1559 (
            .O(N__15091),
            .I(v33dsw_ok));
    CascadeMux I__1558 (
            .O(N__15088),
            .I(N__15082));
    CascadeMux I__1557 (
            .O(N__15087),
            .I(N__15079));
    CascadeMux I__1556 (
            .O(N__15086),
            .I(N__15076));
    InMux I__1555 (
            .O(N__15085),
            .I(N__15072));
    InMux I__1554 (
            .O(N__15082),
            .I(N__15063));
    InMux I__1553 (
            .O(N__15079),
            .I(N__15063));
    InMux I__1552 (
            .O(N__15076),
            .I(N__15063));
    InMux I__1551 (
            .O(N__15075),
            .I(N__15063));
    LocalMux I__1550 (
            .O(N__15072),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__1549 (
            .O(N__15063),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    InMux I__1548 (
            .O(N__15058),
            .I(N__15055));
    LocalMux I__1547 (
            .O(N__15055),
            .I(N__15050));
    InMux I__1546 (
            .O(N__15054),
            .I(N__15045));
    InMux I__1545 (
            .O(N__15053),
            .I(N__15045));
    Odrv4 I__1544 (
            .O(N__15050),
            .I(\DSW_PWRGD.N_1_i ));
    LocalMux I__1543 (
            .O(N__15045),
            .I(\DSW_PWRGD.N_1_i ));
    InMux I__1542 (
            .O(N__15040),
            .I(N__15037));
    LocalMux I__1541 (
            .O(N__15037),
            .I(N__15034));
    Span12Mux_s8_h I__1540 (
            .O(N__15034),
            .I(N__15031));
    Odrv12 I__1539 (
            .O(N__15031),
            .I(gpio_fpga_soc_1));
    CascadeMux I__1538 (
            .O(N__15028),
            .I(N__15024));
    InMux I__1537 (
            .O(N__15027),
            .I(N__15007));
    InMux I__1536 (
            .O(N__15024),
            .I(N__15007));
    InMux I__1535 (
            .O(N__15023),
            .I(N__15007));
    InMux I__1534 (
            .O(N__15022),
            .I(N__15003));
    InMux I__1533 (
            .O(N__15021),
            .I(N__14992));
    InMux I__1532 (
            .O(N__15020),
            .I(N__14992));
    InMux I__1531 (
            .O(N__15019),
            .I(N__14992));
    InMux I__1530 (
            .O(N__15018),
            .I(N__14992));
    InMux I__1529 (
            .O(N__15017),
            .I(N__14992));
    InMux I__1528 (
            .O(N__15016),
            .I(N__14989));
    InMux I__1527 (
            .O(N__15015),
            .I(N__14986));
    InMux I__1526 (
            .O(N__15014),
            .I(N__14983));
    LocalMux I__1525 (
            .O(N__15007),
            .I(N__14980));
    InMux I__1524 (
            .O(N__15006),
            .I(N__14977));
    LocalMux I__1523 (
            .O(N__15003),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__1522 (
            .O(N__14992),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__1521 (
            .O(N__14989),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__1520 (
            .O(N__14986),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__1519 (
            .O(N__14983),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    Odrv4 I__1518 (
            .O(N__14980),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    LocalMux I__1517 (
            .O(N__14977),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    CascadeMux I__1516 (
            .O(N__14962),
            .I(\HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_ ));
    InMux I__1515 (
            .O(N__14959),
            .I(N__14956));
    LocalMux I__1514 (
            .O(N__14956),
            .I(\HDA_STRAP.curr_state_RNO_0Z0Z_0 ));
    CascadeMux I__1513 (
            .O(N__14953),
            .I(N__14945));
    CascadeMux I__1512 (
            .O(N__14952),
            .I(N__14942));
    CascadeMux I__1511 (
            .O(N__14951),
            .I(N__14938));
    CascadeMux I__1510 (
            .O(N__14950),
            .I(N__14933));
    CascadeMux I__1509 (
            .O(N__14949),
            .I(N__14930));
    CascadeMux I__1508 (
            .O(N__14948),
            .I(N__14925));
    InMux I__1507 (
            .O(N__14945),
            .I(N__14918));
    InMux I__1506 (
            .O(N__14942),
            .I(N__14918));
    InMux I__1505 (
            .O(N__14941),
            .I(N__14915));
    InMux I__1504 (
            .O(N__14938),
            .I(N__14908));
    InMux I__1503 (
            .O(N__14937),
            .I(N__14908));
    InMux I__1502 (
            .O(N__14936),
            .I(N__14908));
    InMux I__1501 (
            .O(N__14933),
            .I(N__14900));
    InMux I__1500 (
            .O(N__14930),
            .I(N__14900));
    InMux I__1499 (
            .O(N__14929),
            .I(N__14900));
    InMux I__1498 (
            .O(N__14928),
            .I(N__14891));
    InMux I__1497 (
            .O(N__14925),
            .I(N__14891));
    InMux I__1496 (
            .O(N__14924),
            .I(N__14891));
    InMux I__1495 (
            .O(N__14923),
            .I(N__14891));
    LocalMux I__1494 (
            .O(N__14918),
            .I(N__14884));
    LocalMux I__1493 (
            .O(N__14915),
            .I(N__14884));
    LocalMux I__1492 (
            .O(N__14908),
            .I(N__14884));
    InMux I__1491 (
            .O(N__14907),
            .I(N__14881));
    LocalMux I__1490 (
            .O(N__14900),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__1489 (
            .O(N__14891),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    Odrv12 I__1488 (
            .O(N__14884),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__1487 (
            .O(N__14881),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    InMux I__1486 (
            .O(N__14872),
            .I(N__14869));
    LocalMux I__1485 (
            .O(N__14869),
            .I(\HDA_STRAP.N_5_0 ));
    InMux I__1484 (
            .O(N__14866),
            .I(N__14862));
    InMux I__1483 (
            .O(N__14865),
            .I(N__14859));
    LocalMux I__1482 (
            .O(N__14862),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    LocalMux I__1481 (
            .O(N__14859),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    InMux I__1480 (
            .O(N__14854),
            .I(N__14850));
    InMux I__1479 (
            .O(N__14853),
            .I(N__14847));
    LocalMux I__1478 (
            .O(N__14850),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    LocalMux I__1477 (
            .O(N__14847),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    CascadeMux I__1476 (
            .O(N__14842),
            .I(N__14839));
    InMux I__1475 (
            .O(N__14839),
            .I(N__14835));
    InMux I__1474 (
            .O(N__14838),
            .I(N__14832));
    LocalMux I__1473 (
            .O(N__14835),
            .I(N__14829));
    LocalMux I__1472 (
            .O(N__14832),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    Odrv4 I__1471 (
            .O(N__14829),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    InMux I__1470 (
            .O(N__14824),
            .I(N__14820));
    InMux I__1469 (
            .O(N__14823),
            .I(N__14817));
    LocalMux I__1468 (
            .O(N__14820),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    LocalMux I__1467 (
            .O(N__14817),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    CascadeMux I__1466 (
            .O(N__14812),
            .I(\DSW_PWRGD.un4_count_9_cascade_ ));
    InMux I__1465 (
            .O(N__14809),
            .I(N__14805));
    InMux I__1464 (
            .O(N__14808),
            .I(N__14802));
    LocalMux I__1463 (
            .O(N__14805),
            .I(\HDA_STRAP.countZ0Z_15 ));
    LocalMux I__1462 (
            .O(N__14802),
            .I(\HDA_STRAP.countZ0Z_15 ));
    CascadeMux I__1461 (
            .O(N__14797),
            .I(N__14793));
    InMux I__1460 (
            .O(N__14796),
            .I(N__14790));
    InMux I__1459 (
            .O(N__14793),
            .I(N__14787));
    LocalMux I__1458 (
            .O(N__14790),
            .I(\HDA_STRAP.countZ0Z_14 ));
    LocalMux I__1457 (
            .O(N__14787),
            .I(\HDA_STRAP.countZ0Z_14 ));
    InMux I__1456 (
            .O(N__14782),
            .I(N__14779));
    LocalMux I__1455 (
            .O(N__14779),
            .I(N__14776));
    Odrv4 I__1454 (
            .O(N__14776),
            .I(\HDA_STRAP.un4_count_12 ));
    InMux I__1453 (
            .O(N__14773),
            .I(N__14770));
    LocalMux I__1452 (
            .O(N__14770),
            .I(\HDA_STRAP.count_RNO_0Z0Z_6 ));
    InMux I__1451 (
            .O(N__14767),
            .I(N__14763));
    InMux I__1450 (
            .O(N__14766),
            .I(N__14760));
    LocalMux I__1449 (
            .O(N__14763),
            .I(\HDA_STRAP.countZ0Z_6 ));
    LocalMux I__1448 (
            .O(N__14760),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__1447 (
            .O(N__14755),
            .I(N__14752));
    LocalMux I__1446 (
            .O(N__14752),
            .I(\HDA_STRAP.count_RNO_0Z0Z_8 ));
    InMux I__1445 (
            .O(N__14749),
            .I(N__14745));
    InMux I__1444 (
            .O(N__14748),
            .I(N__14742));
    LocalMux I__1443 (
            .O(N__14745),
            .I(\HDA_STRAP.countZ0Z_8 ));
    LocalMux I__1442 (
            .O(N__14742),
            .I(\HDA_STRAP.countZ0Z_8 ));
    InMux I__1441 (
            .O(N__14737),
            .I(N__14734));
    LocalMux I__1440 (
            .O(N__14734),
            .I(\HDA_STRAP.count_RNO_0Z0Z_11 ));
    InMux I__1439 (
            .O(N__14731),
            .I(N__14727));
    InMux I__1438 (
            .O(N__14730),
            .I(N__14724));
    LocalMux I__1437 (
            .O(N__14727),
            .I(\HDA_STRAP.countZ0Z_11 ));
    LocalMux I__1436 (
            .O(N__14724),
            .I(\HDA_STRAP.countZ0Z_11 ));
    CascadeMux I__1435 (
            .O(N__14719),
            .I(\HDA_STRAP.N_14_cascade_ ));
    InMux I__1434 (
            .O(N__14716),
            .I(N__14705));
    InMux I__1433 (
            .O(N__14715),
            .I(N__14694));
    InMux I__1432 (
            .O(N__14714),
            .I(N__14694));
    InMux I__1431 (
            .O(N__14713),
            .I(N__14694));
    InMux I__1430 (
            .O(N__14712),
            .I(N__14694));
    InMux I__1429 (
            .O(N__14711),
            .I(N__14694));
    InMux I__1428 (
            .O(N__14710),
            .I(N__14687));
    InMux I__1427 (
            .O(N__14709),
            .I(N__14687));
    InMux I__1426 (
            .O(N__14708),
            .I(N__14687));
    LocalMux I__1425 (
            .O(N__14705),
            .I(N__14684));
    LocalMux I__1424 (
            .O(N__14694),
            .I(\HDA_STRAP.un4_count ));
    LocalMux I__1423 (
            .O(N__14687),
            .I(\HDA_STRAP.un4_count ));
    Odrv4 I__1422 (
            .O(N__14684),
            .I(\HDA_STRAP.un4_count ));
    InMux I__1421 (
            .O(N__14677),
            .I(N__14673));
    InMux I__1420 (
            .O(N__14676),
            .I(N__14670));
    LocalMux I__1419 (
            .O(N__14673),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    LocalMux I__1418 (
            .O(N__14670),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    IoInMux I__1417 (
            .O(N__14665),
            .I(N__14662));
    LocalMux I__1416 (
            .O(N__14662),
            .I(N__14659));
    IoSpan4Mux I__1415 (
            .O(N__14659),
            .I(N__14656));
    Span4Mux_s1_h I__1414 (
            .O(N__14656),
            .I(N__14653));
    Odrv4 I__1413 (
            .O(N__14653),
            .I(hda_sdo_atp));
    InMux I__1412 (
            .O(N__14650),
            .I(N__14647));
    LocalMux I__1411 (
            .O(N__14647),
            .I(\HDA_STRAP.count_RNO_0Z0Z_0 ));
    CascadeMux I__1410 (
            .O(N__14644),
            .I(\HDA_STRAP.un4_count_cascade_ ));
    InMux I__1409 (
            .O(N__14641),
            .I(N__14637));
    InMux I__1408 (
            .O(N__14640),
            .I(N__14634));
    LocalMux I__1407 (
            .O(N__14637),
            .I(\HDA_STRAP.countZ0Z_2 ));
    LocalMux I__1406 (
            .O(N__14634),
            .I(\HDA_STRAP.countZ0Z_2 ));
    InMux I__1405 (
            .O(N__14629),
            .I(N__14625));
    InMux I__1404 (
            .O(N__14628),
            .I(N__14622));
    LocalMux I__1403 (
            .O(N__14625),
            .I(\HDA_STRAP.countZ0Z_4 ));
    LocalMux I__1402 (
            .O(N__14622),
            .I(\HDA_STRAP.countZ0Z_4 ));
    CascadeMux I__1401 (
            .O(N__14617),
            .I(N__14614));
    InMux I__1400 (
            .O(N__14614),
            .I(N__14610));
    InMux I__1399 (
            .O(N__14613),
            .I(N__14607));
    LocalMux I__1398 (
            .O(N__14610),
            .I(\HDA_STRAP.countZ0Z_3 ));
    LocalMux I__1397 (
            .O(N__14607),
            .I(\HDA_STRAP.countZ0Z_3 ));
    InMux I__1396 (
            .O(N__14602),
            .I(N__14598));
    InMux I__1395 (
            .O(N__14601),
            .I(N__14595));
    LocalMux I__1394 (
            .O(N__14598),
            .I(\HDA_STRAP.countZ0Z_5 ));
    LocalMux I__1393 (
            .O(N__14595),
            .I(\HDA_STRAP.countZ0Z_5 ));
    InMux I__1392 (
            .O(N__14590),
            .I(N__14587));
    LocalMux I__1391 (
            .O(N__14587),
            .I(\HDA_STRAP.un4_count_10 ));
    InMux I__1390 (
            .O(N__14584),
            .I(N__14581));
    LocalMux I__1389 (
            .O(N__14581),
            .I(N__14578));
    Odrv4 I__1388 (
            .O(N__14578),
            .I(\HDA_STRAP.count_RNO_0Z0Z_17 ));
    InMux I__1387 (
            .O(N__14575),
            .I(N__14571));
    InMux I__1386 (
            .O(N__14574),
            .I(N__14568));
    LocalMux I__1385 (
            .O(N__14571),
            .I(\HDA_STRAP.countZ0Z_1 ));
    LocalMux I__1384 (
            .O(N__14568),
            .I(\HDA_STRAP.countZ0Z_1 ));
    CascadeMux I__1383 (
            .O(N__14563),
            .I(N__14560));
    InMux I__1382 (
            .O(N__14560),
            .I(N__14557));
    LocalMux I__1381 (
            .O(N__14557),
            .I(N__14554));
    Span4Mux_s2_h I__1380 (
            .O(N__14554),
            .I(N__14550));
    InMux I__1379 (
            .O(N__14553),
            .I(N__14547));
    Odrv4 I__1378 (
            .O(N__14550),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__1377 (
            .O(N__14547),
            .I(\HDA_STRAP.countZ0Z_0 ));
    InMux I__1376 (
            .O(N__14542),
            .I(N__14539));
    LocalMux I__1375 (
            .O(N__14539),
            .I(N__14535));
    InMux I__1374 (
            .O(N__14538),
            .I(N__14532));
    Odrv4 I__1373 (
            .O(N__14535),
            .I(\HDA_STRAP.countZ0Z_17 ));
    LocalMux I__1372 (
            .O(N__14532),
            .I(\HDA_STRAP.countZ0Z_17 ));
    CascadeMux I__1371 (
            .O(N__14527),
            .I(\HDA_STRAP.un4_count_9_cascade_ ));
    InMux I__1370 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__1369 (
            .O(N__14521),
            .I(\HDA_STRAP.un4_count_13 ));
    CascadeMux I__1368 (
            .O(N__14518),
            .I(N__14515));
    InMux I__1367 (
            .O(N__14515),
            .I(N__14512));
    LocalMux I__1366 (
            .O(N__14512),
            .I(N__14509));
    Odrv4 I__1365 (
            .O(N__14509),
            .I(\HDA_STRAP.count_RNO_0Z0Z_16 ));
    InMux I__1364 (
            .O(N__14506),
            .I(N__14503));
    LocalMux I__1363 (
            .O(N__14503),
            .I(N__14499));
    InMux I__1362 (
            .O(N__14502),
            .I(N__14496));
    Odrv4 I__1361 (
            .O(N__14499),
            .I(\HDA_STRAP.countZ0Z_16 ));
    LocalMux I__1360 (
            .O(N__14496),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__1359 (
            .O(N__14491),
            .I(N__14488));
    LocalMux I__1358 (
            .O(N__14488),
            .I(\HDA_STRAP.count_RNO_0Z0Z_10 ));
    InMux I__1357 (
            .O(N__14485),
            .I(N__14481));
    InMux I__1356 (
            .O(N__14484),
            .I(N__14478));
    LocalMux I__1355 (
            .O(N__14481),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__1354 (
            .O(N__14478),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__1353 (
            .O(N__14473),
            .I(N__14469));
    InMux I__1352 (
            .O(N__14472),
            .I(N__14466));
    LocalMux I__1351 (
            .O(N__14469),
            .I(\HDA_STRAP.countZ0Z_12 ));
    LocalMux I__1350 (
            .O(N__14466),
            .I(\HDA_STRAP.countZ0Z_12 ));
    InMux I__1349 (
            .O(N__14461),
            .I(N__14457));
    InMux I__1348 (
            .O(N__14460),
            .I(N__14454));
    LocalMux I__1347 (
            .O(N__14457),
            .I(\HDA_STRAP.countZ0Z_9 ));
    LocalMux I__1346 (
            .O(N__14454),
            .I(\HDA_STRAP.countZ0Z_9 ));
    CascadeMux I__1345 (
            .O(N__14449),
            .I(N__14445));
    InMux I__1344 (
            .O(N__14448),
            .I(N__14442));
    InMux I__1343 (
            .O(N__14445),
            .I(N__14439));
    LocalMux I__1342 (
            .O(N__14442),
            .I(\HDA_STRAP.countZ0Z_13 ));
    LocalMux I__1341 (
            .O(N__14439),
            .I(\HDA_STRAP.countZ0Z_13 ));
    InMux I__1340 (
            .O(N__14434),
            .I(N__14430));
    InMux I__1339 (
            .O(N__14433),
            .I(N__14427));
    LocalMux I__1338 (
            .O(N__14430),
            .I(\HDA_STRAP.countZ0Z_7 ));
    LocalMux I__1337 (
            .O(N__14427),
            .I(\HDA_STRAP.countZ0Z_7 ));
    CascadeMux I__1336 (
            .O(N__14422),
            .I(N__14419));
    InMux I__1335 (
            .O(N__14419),
            .I(N__14416));
    LocalMux I__1334 (
            .O(N__14416),
            .I(\HDA_STRAP.un4_count_11 ));
    InMux I__1333 (
            .O(N__14413),
            .I(N__14410));
    LocalMux I__1332 (
            .O(N__14410),
            .I(N__14407));
    Odrv12 I__1331 (
            .O(N__14407),
            .I(\POWERLED.un85_clk_100khz_5 ));
    CascadeMux I__1330 (
            .O(N__14404),
            .I(N__14401));
    InMux I__1329 (
            .O(N__14401),
            .I(N__14398));
    LocalMux I__1328 (
            .O(N__14398),
            .I(\POWERLED.un85_clk_100khz_9 ));
    InMux I__1327 (
            .O(N__14395),
            .I(N__14392));
    LocalMux I__1326 (
            .O(N__14392),
            .I(N__14389));
    Odrv4 I__1325 (
            .O(N__14389),
            .I(\POWERLED.un85_clk_100khz_8 ));
    CascadeMux I__1324 (
            .O(N__14386),
            .I(N__14383));
    InMux I__1323 (
            .O(N__14383),
            .I(N__14380));
    LocalMux I__1322 (
            .O(N__14380),
            .I(N__14377));
    Odrv4 I__1321 (
            .O(N__14377),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    CascadeMux I__1320 (
            .O(N__14374),
            .I(N__14371));
    InMux I__1319 (
            .O(N__14371),
            .I(N__14368));
    LocalMux I__1318 (
            .O(N__14368),
            .I(N__14365));
    Odrv4 I__1317 (
            .O(N__14365),
            .I(\POWERLED.un85_clk_100khz_10 ));
    CascadeMux I__1316 (
            .O(N__14362),
            .I(N__14359));
    InMux I__1315 (
            .O(N__14359),
            .I(N__14356));
    LocalMux I__1314 (
            .O(N__14356),
            .I(N__14353));
    Odrv12 I__1313 (
            .O(N__14353),
            .I(\POWERLED.mult1_un89_sum_i_8 ));
    InMux I__1312 (
            .O(N__14350),
            .I(N__14347));
    LocalMux I__1311 (
            .O(N__14347),
            .I(N__14344));
    Odrv12 I__1310 (
            .O(N__14344),
            .I(\POWERLED.un85_clk_100khz_3 ));
    InMux I__1309 (
            .O(N__14341),
            .I(N__14338));
    LocalMux I__1308 (
            .O(N__14338),
            .I(\POWERLED.N_5118_i ));
    InMux I__1307 (
            .O(N__14335),
            .I(N__14332));
    LocalMux I__1306 (
            .O(N__14332),
            .I(\POWERLED.N_5119_i ));
    InMux I__1305 (
            .O(N__14329),
            .I(N__14326));
    LocalMux I__1304 (
            .O(N__14326),
            .I(\POWERLED.N_5120_i ));
    InMux I__1303 (
            .O(N__14323),
            .I(N__14320));
    LocalMux I__1302 (
            .O(N__14320),
            .I(\POWERLED.N_5121_i ));
    CascadeMux I__1301 (
            .O(N__14317),
            .I(N__14314));
    InMux I__1300 (
            .O(N__14314),
            .I(N__14311));
    LocalMux I__1299 (
            .O(N__14311),
            .I(N__14308));
    Odrv4 I__1298 (
            .O(N__14308),
            .I(\POWERLED.N_5122_i ));
    InMux I__1297 (
            .O(N__14305),
            .I(N__14302));
    LocalMux I__1296 (
            .O(N__14302),
            .I(\POWERLED.N_5123_i ));
    InMux I__1295 (
            .O(N__14299),
            .I(N__14296));
    LocalMux I__1294 (
            .O(N__14296),
            .I(\POWERLED.N_5124_i ));
    InMux I__1293 (
            .O(N__14293),
            .I(bfn_1_15_0_));
    CascadeMux I__1292 (
            .O(N__14290),
            .I(N__14287));
    InMux I__1291 (
            .O(N__14287),
            .I(N__14284));
    LocalMux I__1290 (
            .O(N__14284),
            .I(N__14281));
    Odrv12 I__1289 (
            .O(N__14281),
            .I(\POWERLED.mult1_un82_sum_i_8 ));
    CascadeMux I__1288 (
            .O(N__14278),
            .I(N__14275));
    InMux I__1287 (
            .O(N__14275),
            .I(N__14272));
    LocalMux I__1286 (
            .O(N__14272),
            .I(\POWERLED.N_5110_i ));
    CascadeMux I__1285 (
            .O(N__14269),
            .I(N__14266));
    InMux I__1284 (
            .O(N__14266),
            .I(N__14263));
    LocalMux I__1283 (
            .O(N__14263),
            .I(N__14260));
    Odrv4 I__1282 (
            .O(N__14260),
            .I(\POWERLED.N_5111_i ));
    CascadeMux I__1281 (
            .O(N__14257),
            .I(N__14254));
    InMux I__1280 (
            .O(N__14254),
            .I(N__14251));
    LocalMux I__1279 (
            .O(N__14251),
            .I(N__14248));
    Odrv4 I__1278 (
            .O(N__14248),
            .I(\POWERLED.N_5112_i ));
    CascadeMux I__1277 (
            .O(N__14245),
            .I(N__14242));
    InMux I__1276 (
            .O(N__14242),
            .I(N__14239));
    LocalMux I__1275 (
            .O(N__14239),
            .I(\POWERLED.N_5113_i ));
    CascadeMux I__1274 (
            .O(N__14236),
            .I(N__14233));
    InMux I__1273 (
            .O(N__14233),
            .I(N__14230));
    LocalMux I__1272 (
            .O(N__14230),
            .I(\POWERLED.N_5114_i ));
    CascadeMux I__1271 (
            .O(N__14227),
            .I(N__14224));
    InMux I__1270 (
            .O(N__14224),
            .I(N__14221));
    LocalMux I__1269 (
            .O(N__14221),
            .I(\POWERLED.N_5115_i ));
    CascadeMux I__1268 (
            .O(N__14218),
            .I(N__14215));
    InMux I__1267 (
            .O(N__14215),
            .I(N__14212));
    LocalMux I__1266 (
            .O(N__14212),
            .I(N__14209));
    Odrv4 I__1265 (
            .O(N__14209),
            .I(\POWERLED.N_5116_i ));
    CascadeMux I__1264 (
            .O(N__14206),
            .I(N__14203));
    InMux I__1263 (
            .O(N__14203),
            .I(N__14200));
    LocalMux I__1262 (
            .O(N__14200),
            .I(\POWERLED.N_5117_i ));
    InMux I__1261 (
            .O(N__14197),
            .I(N__14191));
    InMux I__1260 (
            .O(N__14196),
            .I(N__14191));
    LocalMux I__1259 (
            .O(N__14191),
            .I(\POWERLED.g0_i_o3_0 ));
    CascadeMux I__1258 (
            .O(N__14188),
            .I(\POWERLED.un79_clk_100khzlt6_cascade_ ));
    CascadeMux I__1257 (
            .O(N__14185),
            .I(\POWERLED.un79_clk_100khzlto15_5_cascade_ ));
    CascadeMux I__1256 (
            .O(N__14182),
            .I(\POWERLED.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__1255 (
            .O(N__14179),
            .I(N__14176));
    LocalMux I__1254 (
            .O(N__14176),
            .I(\POWERLED.un79_clk_100khzlto15_3 ));
    CascadeMux I__1253 (
            .O(N__14173),
            .I(\POWERLED.count_RNIZ0Z_8_cascade_ ));
    SRMux I__1252 (
            .O(N__14170),
            .I(N__14167));
    LocalMux I__1251 (
            .O(N__14167),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    InMux I__1250 (
            .O(N__14164),
            .I(N__14158));
    InMux I__1249 (
            .O(N__14163),
            .I(N__14158));
    LocalMux I__1248 (
            .O(N__14158),
            .I(\POWERLED.N_8 ));
    CascadeMux I__1247 (
            .O(N__14155),
            .I(N__14152));
    InMux I__1246 (
            .O(N__14152),
            .I(N__14149));
    LocalMux I__1245 (
            .O(N__14149),
            .I(\POWERLED.un1_count_cry_0_i ));
    InMux I__1244 (
            .O(N__14146),
            .I(N__14143));
    LocalMux I__1243 (
            .O(N__14143),
            .I(\POWERLED.count_0_12 ));
    IoInMux I__1242 (
            .O(N__14140),
            .I(N__14137));
    LocalMux I__1241 (
            .O(N__14137),
            .I(N__14134));
    Span4Mux_s0_v I__1240 (
            .O(N__14134),
            .I(N__14131));
    Span4Mux_v I__1239 (
            .O(N__14131),
            .I(N__14128));
    Odrv4 I__1238 (
            .O(N__14128),
            .I(pwrbtn_led));
    CascadeMux I__1237 (
            .O(N__14125),
            .I(\POWERLED.curr_state_3_0_cascade_ ));
    CascadeMux I__1236 (
            .O(N__14122),
            .I(\POWERLED.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__1235 (
            .O(N__14119),
            .I(\POWERLED.count_0_sqmuxa_i_cascade_ ));
    CascadeMux I__1234 (
            .O(N__14116),
            .I(\POWERLED.count_1_0_cascade_ ));
    InMux I__1233 (
            .O(N__14113),
            .I(N__14110));
    LocalMux I__1232 (
            .O(N__14110),
            .I(\POWERLED.count_0_0 ));
    InMux I__1231 (
            .O(N__14107),
            .I(N__14101));
    InMux I__1230 (
            .O(N__14106),
            .I(N__14101));
    LocalMux I__1229 (
            .O(N__14101),
            .I(\POWERLED.pwm_outZ0 ));
    InMux I__1228 (
            .O(N__14098),
            .I(N__14095));
    LocalMux I__1227 (
            .O(N__14095),
            .I(\POWERLED.count_0_5 ));
    InMux I__1226 (
            .O(N__14092),
            .I(N__14089));
    LocalMux I__1225 (
            .O(N__14089),
            .I(\POWERLED.count_0_14 ));
    CascadeMux I__1224 (
            .O(N__14086),
            .I(\POWERLED.count_1_1_cascade_ ));
    CascadeMux I__1223 (
            .O(N__14083),
            .I(\POWERLED.countZ0Z_1_cascade_ ));
    InMux I__1222 (
            .O(N__14080),
            .I(N__14077));
    LocalMux I__1221 (
            .O(N__14077),
            .I(\POWERLED.count_0_1 ));
    InMux I__1220 (
            .O(N__14074),
            .I(N__14071));
    LocalMux I__1219 (
            .O(N__14071),
            .I(\POWERLED.count_0_3 ));
    InMux I__1218 (
            .O(N__14068),
            .I(\DSW_PWRGD.un1_count_1_cry_11 ));
    InMux I__1217 (
            .O(N__14065),
            .I(\DSW_PWRGD.un1_count_1_cry_12 ));
    InMux I__1216 (
            .O(N__14062),
            .I(\DSW_PWRGD.un1_count_1_cry_13 ));
    InMux I__1215 (
            .O(N__14059),
            .I(bfn_1_7_0_));
    InMux I__1214 (
            .O(N__14056),
            .I(N__14053));
    LocalMux I__1213 (
            .O(N__14053),
            .I(\POWERLED.count_0_4 ));
    InMux I__1212 (
            .O(N__14050),
            .I(N__14047));
    LocalMux I__1211 (
            .O(N__14047),
            .I(\POWERLED.count_0_13 ));
    InMux I__1210 (
            .O(N__14044),
            .I(\DSW_PWRGD.un1_count_1_cry_2 ));
    InMux I__1209 (
            .O(N__14041),
            .I(\DSW_PWRGD.un1_count_1_cry_3 ));
    InMux I__1208 (
            .O(N__14038),
            .I(\DSW_PWRGD.un1_count_1_cry_4 ));
    InMux I__1207 (
            .O(N__14035),
            .I(\DSW_PWRGD.un1_count_1_cry_5 ));
    InMux I__1206 (
            .O(N__14032),
            .I(\DSW_PWRGD.un1_count_1_cry_6 ));
    InMux I__1205 (
            .O(N__14029),
            .I(bfn_1_6_0_));
    InMux I__1204 (
            .O(N__14026),
            .I(\DSW_PWRGD.un1_count_1_cry_8 ));
    InMux I__1203 (
            .O(N__14023),
            .I(\DSW_PWRGD.un1_count_1_cry_9 ));
    InMux I__1202 (
            .O(N__14020),
            .I(\DSW_PWRGD.un1_count_1_cry_10 ));
    InMux I__1201 (
            .O(N__14017),
            .I(\HDA_STRAP.un1_count_1_cry_12 ));
    InMux I__1200 (
            .O(N__14014),
            .I(\HDA_STRAP.un1_count_1_cry_13 ));
    InMux I__1199 (
            .O(N__14011),
            .I(\HDA_STRAP.un1_count_1_cry_14 ));
    InMux I__1198 (
            .O(N__14008),
            .I(bfn_1_3_0_));
    InMux I__1197 (
            .O(N__14005),
            .I(\HDA_STRAP.un1_count_1_cry_16 ));
    CascadeMux I__1196 (
            .O(N__14002),
            .I(N__13998));
    InMux I__1195 (
            .O(N__14001),
            .I(N__13995));
    InMux I__1194 (
            .O(N__13998),
            .I(N__13992));
    LocalMux I__1193 (
            .O(N__13995),
            .I(N__13987));
    LocalMux I__1192 (
            .O(N__13992),
            .I(N__13987));
    Odrv4 I__1191 (
            .O(N__13987),
            .I(\HDA_STRAP.curr_state_RNIH91AZ0Z_1 ));
    InMux I__1190 (
            .O(N__13984),
            .I(\DSW_PWRGD.un1_count_1_cry_0 ));
    InMux I__1189 (
            .O(N__13981),
            .I(\DSW_PWRGD.un1_count_1_cry_1 ));
    InMux I__1188 (
            .O(N__13978),
            .I(\HDA_STRAP.un1_count_1_cry_3 ));
    InMux I__1187 (
            .O(N__13975),
            .I(\HDA_STRAP.un1_count_1_cry_4 ));
    InMux I__1186 (
            .O(N__13972),
            .I(\HDA_STRAP.un1_count_1_cry_5 ));
    InMux I__1185 (
            .O(N__13969),
            .I(\HDA_STRAP.un1_count_1_cry_6 ));
    InMux I__1184 (
            .O(N__13966),
            .I(bfn_1_2_0_));
    InMux I__1183 (
            .O(N__13963),
            .I(\HDA_STRAP.un1_count_1_cry_8 ));
    InMux I__1182 (
            .O(N__13960),
            .I(\HDA_STRAP.un1_count_1_cry_9 ));
    InMux I__1181 (
            .O(N__13957),
            .I(\HDA_STRAP.un1_count_1_cry_10 ));
    InMux I__1180 (
            .O(N__13954),
            .I(\HDA_STRAP.un1_count_1_cry_11 ));
    InMux I__1179 (
            .O(N__13951),
            .I(\HDA_STRAP.un1_count_1_cry_0 ));
    InMux I__1178 (
            .O(N__13948),
            .I(\HDA_STRAP.un1_count_1_cry_1 ));
    InMux I__1177 (
            .O(N__13945),
            .I(\HDA_STRAP.un1_count_1_cry_2 ));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_4_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_16_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(COUNTER_un4_counter_7),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_5_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_1_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7 ),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_1_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_1_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_7 ),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(\HDA_STRAP.un1_count_1_cry_15 ),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_1_7_0_));
    ICE_GB N_29_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__22537),
            .GLOBALBUFFEROUTPUT(N_29_g));
    ICE_GB N_570_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__29826),
            .GLOBALBUFFEROUTPUT(N_570_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_0_LC_1_1_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_0_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_0_LC_1_1_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_0_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(N__14553),
            .in2(N__14002),
            .in3(N__14001),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_1_1_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_1_1_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_1_LC_1_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_1_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_1_LC_1_1_1  (
            .in0(_gnd_net_),
            .in1(N__14574),
            .in2(_gnd_net_),
            .in3(N__13951),
            .lcout(\HDA_STRAP.countZ0Z_1 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_0 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_1 ),
            .clk(N__34372),
            .ce(N__34689),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_1_1_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_2_LC_1_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_1_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_2_LC_1_1_2  (
            .in0(_gnd_net_),
            .in1(N__14641),
            .in2(_gnd_net_),
            .in3(N__13948),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_2 ),
            .clk(N__34372),
            .ce(N__34689),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_1_1_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_3_LC_1_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_1_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_3_LC_1_1_3  (
            .in0(_gnd_net_),
            .in1(N__14613),
            .in2(_gnd_net_),
            .in3(N__13945),
            .lcout(\HDA_STRAP.countZ0Z_3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_3 ),
            .clk(N__34372),
            .ce(N__34689),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_1_1_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_4_LC_1_1_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_1_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_4_LC_1_1_4  (
            .in0(_gnd_net_),
            .in1(N__14629),
            .in2(_gnd_net_),
            .in3(N__13978),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_4 ),
            .clk(N__34372),
            .ce(N__34689),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_1_1_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_5_LC_1_1_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_1_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_5_LC_1_1_5  (
            .in0(_gnd_net_),
            .in1(N__14602),
            .in2(_gnd_net_),
            .in3(N__13975),
            .lcout(\HDA_STRAP.countZ0Z_5 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_5 ),
            .clk(N__34372),
            .ce(N__34689),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_6_LC_1_1_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_6_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_6_LC_1_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_6_LC_1_1_6  (
            .in0(_gnd_net_),
            .in1(N__14767),
            .in2(_gnd_net_),
            .in3(N__13972),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_5 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_1_1_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_7_LC_1_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_1_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_7_LC_1_1_7  (
            .in0(_gnd_net_),
            .in1(N__14434),
            .in2(_gnd_net_),
            .in3(N__13969),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_7 ),
            .clk(N__34372),
            .ce(N__34689),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_8_LC_1_2_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_8_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_8_LC_1_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_8_LC_1_2_0  (
            .in0(_gnd_net_),
            .in1(N__14749),
            .in2(_gnd_net_),
            .in3(N__13966),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_1_2_1 .C_ON=1'b1;
    defparam \HDA_STRAP.count_9_LC_1_2_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_1_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_9_LC_1_2_1  (
            .in0(_gnd_net_),
            .in1(N__14461),
            .in2(_gnd_net_),
            .in3(N__13963),
            .lcout(\HDA_STRAP.countZ0Z_9 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_8 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_9 ),
            .clk(N__34389),
            .ce(N__34711),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_10_LC_1_2_2 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_10_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_10_LC_1_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_10_LC_1_2_2  (
            .in0(_gnd_net_),
            .in1(N__14485),
            .in2(_gnd_net_),
            .in3(N__13960),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_11_LC_1_2_3 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_11_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_11_LC_1_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_11_LC_1_2_3  (
            .in0(_gnd_net_),
            .in1(N__14731),
            .in2(_gnd_net_),
            .in3(N__13957),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_1_2_4 .C_ON=1'b1;
    defparam \HDA_STRAP.count_12_LC_1_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_1_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_12_LC_1_2_4  (
            .in0(_gnd_net_),
            .in1(N__14473),
            .in2(_gnd_net_),
            .in3(N__13954),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_12 ),
            .clk(N__34389),
            .ce(N__34711),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_1_2_5 .C_ON=1'b1;
    defparam \HDA_STRAP.count_13_LC_1_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_1_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_13_LC_1_2_5  (
            .in0(_gnd_net_),
            .in1(N__14448),
            .in2(_gnd_net_),
            .in3(N__14017),
            .lcout(\HDA_STRAP.countZ0Z_13 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_13 ),
            .clk(N__34389),
            .ce(N__34711),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_1_2_6 .C_ON=1'b1;
    defparam \HDA_STRAP.count_14_LC_1_2_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_1_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_14_LC_1_2_6  (
            .in0(_gnd_net_),
            .in1(N__14796),
            .in2(_gnd_net_),
            .in3(N__14014),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_14 ),
            .clk(N__34389),
            .ce(N__34711),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_1_2_7 .C_ON=1'b1;
    defparam \HDA_STRAP.count_15_LC_1_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_1_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_15_LC_1_2_7  (
            .in0(_gnd_net_),
            .in1(N__14809),
            .in2(_gnd_net_),
            .in3(N__14011),
            .lcout(\HDA_STRAP.countZ0Z_15 ),
            .ltout(),
            .carryin(\HDA_STRAP.un1_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un1_count_1_cry_15 ),
            .clk(N__34389),
            .ce(N__34711),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_16_LC_1_3_0 .C_ON=1'b1;
    defparam \HDA_STRAP.count_RNO_0_16_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_16_LC_1_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNO_0_16_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__14506),
            .in2(_gnd_net_),
            .in3(N__14008),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\HDA_STRAP.un1_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNO_0_17_LC_1_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNO_0_17_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNO_0_17_LC_1_3_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \HDA_STRAP.count_RNO_0_17_LC_1_3_1  (
            .in0(_gnd_net_),
            .in1(N__14542),
            .in2(_gnd_net_),
            .in3(N__14005),
            .lcout(\HDA_STRAP.count_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIH91A_1_LC_1_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIH91A_1_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIH91A_1_LC_1_3_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \HDA_STRAP.curr_state_RNIH91A_1_LC_1_3_2  (
            .in0(N__14907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15006),
            .lcout(\HDA_STRAP.curr_state_RNIH91AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_0_LC_1_5_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_0_LC_1_5_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_0_LC_1_5_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_0_LC_1_5_0  (
            .in0(N__34866),
            .in1(N__15169),
            .in2(N__15151),
            .in3(N__15150),
            .lcout(\DSW_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_0 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_1_LC_1_5_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_1_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_1_LC_1_5_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_1_LC_1_5_1  (
            .in0(N__34862),
            .in1(N__16566),
            .in2(_gnd_net_),
            .in3(N__13984),
            .lcout(\DSW_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_0 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_1 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_2_LC_1_5_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_2_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_2_LC_1_5_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_2_LC_1_5_2  (
            .in0(N__34867),
            .in1(N__15265),
            .in2(_gnd_net_),
            .in3(N__13981),
            .lcout(\DSW_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_1 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_2 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_3_LC_1_5_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_3_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_3_LC_1_5_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_3_LC_1_5_3  (
            .in0(N__34863),
            .in1(N__15226),
            .in2(_gnd_net_),
            .in3(N__14044),
            .lcout(\DSW_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_2 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_3 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_4_LC_1_5_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_4_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_4_LC_1_5_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_4_LC_1_5_4  (
            .in0(N__34868),
            .in1(N__16515),
            .in2(_gnd_net_),
            .in3(N__14041),
            .lcout(\DSW_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_3 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_4 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_5_LC_1_5_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_5_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_5_LC_1_5_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_5_LC_1_5_5  (
            .in0(N__34864),
            .in1(N__15253),
            .in2(_gnd_net_),
            .in3(N__14038),
            .lcout(\DSW_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_4 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_5 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_6_LC_1_5_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_6_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_6_LC_1_5_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_6_LC_1_5_6  (
            .in0(N__34869),
            .in1(N__16551),
            .in2(_gnd_net_),
            .in3(N__14035),
            .lcout(\DSW_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_5 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_6 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_7_LC_1_5_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_7_LC_1_5_7 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_7_LC_1_5_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_7_LC_1_5_7  (
            .in0(N__34865),
            .in1(N__15240),
            .in2(_gnd_net_),
            .in3(N__14032),
            .lcout(\DSW_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_6 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_7 ),
            .clk(N__34373),
            .ce(),
            .sr(N__15326));
    defparam \DSW_PWRGD.count_8_LC_1_6_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_8_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_8_LC_1_6_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_8_LC_1_6_0  (
            .in0(N__34891),
            .in1(N__15183),
            .in2(_gnd_net_),
            .in3(N__14029),
            .lcout(\DSW_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_8 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.count_9_LC_1_6_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_9_LC_1_6_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_9_LC_1_6_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_9_LC_1_6_1  (
            .in0(N__34879),
            .in1(N__16530),
            .in2(_gnd_net_),
            .in3(N__14026),
            .lcout(\DSW_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_8 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_9 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.count_10_LC_1_6_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_10_LC_1_6_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_10_LC_1_6_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_10_LC_1_6_2  (
            .in0(N__34888),
            .in1(N__15196),
            .in2(_gnd_net_),
            .in3(N__14023),
            .lcout(\DSW_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_9 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_10 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.count_11_LC_1_6_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_11_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_11_LC_1_6_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_11_LC_1_6_3  (
            .in0(N__34877),
            .in1(N__15208),
            .in2(_gnd_net_),
            .in3(N__14020),
            .lcout(\DSW_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_10 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_11 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.count_12_LC_1_6_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_12_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_12_LC_1_6_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_12_LC_1_6_4  (
            .in0(N__34889),
            .in1(N__14824),
            .in2(_gnd_net_),
            .in3(N__14068),
            .lcout(\DSW_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_11 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_12 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.count_13_LC_1_6_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_13_LC_1_6_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_13_LC_1_6_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_13_LC_1_6_5  (
            .in0(N__34878),
            .in1(N__14854),
            .in2(_gnd_net_),
            .in3(N__14065),
            .lcout(\DSW_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_12 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_13 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.count_14_LC_1_6_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_14_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_14_LC_1_6_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_14_LC_1_6_6  (
            .in0(N__34890),
            .in1(N__14866),
            .in2(_gnd_net_),
            .in3(N__14062),
            .lcout(\DSW_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_13 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14 ),
            .clk(N__34440),
            .ce(),
            .sr(N__15331));
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_6_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(N__34500),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_14 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_15_LC_1_7_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_15_LC_1_7_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_esr_15_LC_1_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DSW_PWRGD.count_esr_15_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__14838),
            .in2(_gnd_net_),
            .in3(N__14059),
            .lcout(\DSW_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34444),
            .ce(N__15292),
            .sr(N__15330));
    defparam \POWERLED.count_RNI0LHN_4_LC_1_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI0LHN_4_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI0LHN_4_LC_1_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI0LHN_4_LC_1_9_0  (
            .in0(N__14056),
            .in1(N__30613),
            .in2(_gnd_net_),
            .in3(N__15645),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_4_LC_1_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_1_9_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_4_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15649),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34432),
            .ce(N__30781),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI0M6O_13_LC_1_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI0M6O_13_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI0M6O_13_LC_1_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNI0M6O_13_LC_1_9_2  (
            .in0(N__15913),
            .in1(N__14050),
            .in2(_gnd_net_),
            .in3(N__30615),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_13_LC_1_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_1_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_13_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15912),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34432),
            .ce(N__30781),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI2OIN_5_LC_1_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI2OIN_5_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI2OIN_5_LC_1_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI2OIN_5_LC_1_9_4  (
            .in0(N__14098),
            .in1(N__30614),
            .in2(_gnd_net_),
            .in3(N__15606),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_1_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_1_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_1_9_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_5_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15610),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34432),
            .ce(N__30781),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI2P7O_14_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI2P7O_14_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI2P7O_14_LC_1_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNI2P7O_14_LC_1_9_6  (
            .in0(N__15871),
            .in1(N__14092),
            .in2(_gnd_net_),
            .in3(N__30616),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_1_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_1_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_14_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15870),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34432),
            .ce(N__30781),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_1_LC_1_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_1_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_1_LC_1_10_0 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \POWERLED.count_RNI_1_LC_1_10_0  (
            .in0(N__15479),
            .in1(N__15455),
            .in2(_gnd_net_),
            .in3(N__15851),
            .lcout(),
            .ltout(\POWERLED.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGBFE_1_LC_1_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGBFE_1_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGBFE_1_LC_1_10_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \POWERLED.count_RNIGBFE_1_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__30620),
            .in2(N__14086),
            .in3(N__14080),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(\POWERLED.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_1_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_1_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_1_10_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_1_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__15457),
            .in2(N__14083),
            .in3(N__15855),
            .lcout(\POWERLED.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(N__30784),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_1_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_1_10_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_0_LC_1_10_3  (
            .in0(N__15456),
            .in1(_gnd_net_),
            .in2(N__15856),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(N__30784),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUHGN_3_LC_1_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUHGN_3_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUHGN_3_LC_1_10_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \POWERLED.count_RNIUHGN_3_LC_1_10_4  (
            .in0(N__14074),
            .in1(_gnd_net_),
            .in2(N__30631),
            .in3(N__15360),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_1_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_1_10_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_3_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15364),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(N__30784),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIUI5O_12_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIUI5O_12_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIUI5O_12_LC_1_10_6 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \POWERLED.count_RNIUI5O_12_LC_1_10_6  (
            .in0(N__15955),
            .in1(N__14146),
            .in2(N__30632),
            .in3(_gnd_net_),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_1_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_1_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_12_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15954),
            .lcout(\POWERLED.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34429),
            .ce(N__30784),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNIB7P12_LC_1_11_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIB7P12_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIB7P12_LC_1_11_0 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \POWERLED.pwm_out_RNIB7P12_LC_1_11_0  (
            .in0(N__14107),
            .in1(N__14197),
            .in2(N__17883),
            .in3(N__14164),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_1_11_1 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_1_11_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_1_11_1  (
            .in0(N__17844),
            .in1(N__17812),
            .in2(_gnd_net_),
            .in3(N__17872),
            .lcout(),
            .ltout(\POWERLED.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_1_11_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI2P6L_0_LC_1_11_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \POWERLED.curr_state_RNI2P6L_0_LC_1_11_2  (
            .in0(N__17788),
            .in1(_gnd_net_),
            .in2(N__14125),
            .in3(N__30577),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(\POWERLED.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_1_11_3 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIE5D5_0_LC_1_11_3 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \POWERLED.curr_state_RNIE5D5_0_LC_1_11_3  (
            .in0(N__30578),
            .in1(_gnd_net_),
            .in2(N__14122),
            .in3(N__17839),
            .lcout(\POWERLED.count_0_sqmuxa_i ),
            .ltout(\POWERLED.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_0_LC_1_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_0_LC_1_11_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.count_RNI_0_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14119),
            .in3(N__15458),
            .lcout(),
            .ltout(\POWERLED.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIFAFE_0_LC_1_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNIFAFE_0_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIFAFE_0_LC_1_11_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIFAFE_0_LC_1_11_5  (
            .in0(N__30579),
            .in1(_gnd_net_),
            .in2(N__14116),
            .in3(N__14113),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_1_11_6 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_1_11_6 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \POWERLED.pwm_out_LC_1_11_6  (
            .in0(N__14106),
            .in1(N__14196),
            .in2(N__17882),
            .in3(N__14163),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34460),
            .ce(),
            .sr(N__14170));
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_1_11_7 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI1KAM_0_LC_1_11_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.curr_state_RNI1KAM_0_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(N__30809),
            .in2(_gnd_net_),
            .in3(N__17811),
            .lcout(\POWERLED.g0_i_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_2_LC_1_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_2_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_2_LC_1_12_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.count_RNI_2_LC_1_12_0  (
            .in0(N__15423),
            .in1(_gnd_net_),
            .in2(N__15388),
            .in3(N__15669),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_5_LC_1_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_5_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_5_LC_1_12_1 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \POWERLED.count_RNI_5_LC_1_12_1  (
            .in0(N__15630),
            .in1(N__16067),
            .in2(N__14188),
            .in3(N__15731),
            .lcout(\POWERLED.un79_clk_100khzlto15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_1_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_1_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_10_LC_1_12_2  (
            .in0(N__15579),
            .in1(N__15543),
            .in2(N__15942),
            .in3(N__15975),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_15_LC_1_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_15_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_15_LC_1_12_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \POWERLED.count_RNI_15_LC_1_12_3  (
            .in0(N__15893),
            .in1(_gnd_net_),
            .in2(N__14185),
            .in3(N__15686),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_8_LC_1_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_8_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_8_LC_1_12_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNI_8_LC_1_12_4  (
            .in0(N__16019),
            .in1(N__15752),
            .in2(N__14182),
            .in3(N__14179),
            .lcout(\POWERLED.count_RNIZ0Z_8 ),
            .ltout(\POWERLED.count_RNIZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_1_12_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_1_12_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_1_12_5  (
            .in0(N__17814),
            .in1(_gnd_net_),
            .in2(N__14173),
            .in3(N__30630),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIFPNR_0_LC_1_12_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.curr_state_RNIFPNR_0_LC_1_12_6  (
            .in0(N__30810),
            .in1(N__17813),
            .in2(N__30636),
            .in3(N__17843),
            .lcout(\POWERLED.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_1_13_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_1_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__22552),
            .in2(N__14155),
            .in3(N__15463),
            .lcout(\POWERLED.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_1_13_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_1_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_1_13_1  (
            .in0(N__15484),
            .in1(N__22399),
            .in2(N__14278),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5110_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_1_13_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_1_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__20125),
            .in2(N__14269),
            .in3(N__15427),
            .lcout(\POWERLED.N_5111_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_1_13_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_1_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__14350),
            .in2(N__14257),
            .in3(N__15387),
            .lcout(\POWERLED.N_5112_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_1_13_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_1_13_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_1_13_4  (
            .in0(N__15670),
            .in1(N__18709),
            .in2(N__14245),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5113_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_1_13_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_1_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_1_13_5  (
            .in0(N__15634),
            .in1(N__14413),
            .in2(N__14236),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5114_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_1_13_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_1_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__16741),
            .in2(N__14227),
            .in3(N__15735),
            .lcout(\POWERLED.N_5115_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_1_13_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_1_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_1_13_7  (
            .in0(N__16071),
            .in1(N__16132),
            .in2(N__14218),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5116_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_1_14_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_1_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_1_14_0  (
            .in0(N__16030),
            .in1(N__14395),
            .in2(N__14206),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5117_i ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_1_14_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_1_14_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_1_14_1  (
            .in0(N__15757),
            .in1(N__14341),
            .in2(N__14404),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5118_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_1_14_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_1_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_1_14_2  (
            .in0(N__15583),
            .in1(N__14335),
            .in2(N__14374),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5119_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_1_14_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_1_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_1_14_3  (
            .in0(N__15544),
            .in1(N__14329),
            .in2(N__14362),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5120_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_1_14_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_1_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__14323),
            .in2(N__14290),
            .in3(N__15976),
            .lcout(\POWERLED.N_5121_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_1_14_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_1_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_1_14_5  (
            .in0(N__15943),
            .in1(N__17047),
            .in2(N__14317),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5122_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_1_14_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_1_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__14305),
            .in2(N__20188),
            .in3(N__15898),
            .lcout(\POWERLED.N_5123_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_1_14_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_1_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_1_14_7  (
            .in0(N__15694),
            .in1(N__14299),
            .in2(N__14386),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5124_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_1_15_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_1_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14293),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_15_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_15_2  (
            .in0(N__18268),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_15_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18478),
            .lcout(\POWERLED.un85_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_15_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_15_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_1_15_4  (
            .in0(N__17281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_15_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_15_5  (
            .in0(N__16376),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_1_16_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_1_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16255),
            .lcout(\POWERLED.un85_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_1_16_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_1_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18085),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_16_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16428),
            .lcout(\POWERLED.un85_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_1_16_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_1_16_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_1_16_5  (
            .in0(N__17279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22231),
            .lcout(\POWERLED.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_2_1_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB5IA5_2_LC_2_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIB5IA5_2_LC_2_1_0  (
            .in0(N__14782),
            .in1(N__14590),
            .in2(N__14422),
            .in3(N__14524),
            .lcout(\HDA_STRAP.un4_count ),
            .ltout(\HDA_STRAP.un4_count_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_2_1_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_2_1_1 .LUT_INIT=16'b1000101010101010;
    LogicCell40 \HDA_STRAP.count_0_LC_2_1_1  (
            .in0(N__14650),
            .in1(N__15014),
            .in2(N__14644),
            .in3(N__14941),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34195),
            .ce(N__34688),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI2L821_2_LC_2_1_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI2L821_2_LC_2_1_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNI2L821_2_LC_2_1_2  (
            .in0(N__14640),
            .in1(N__14628),
            .in2(N__14617),
            .in3(N__14601),
            .lcout(\HDA_STRAP.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_2_1_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_2_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_2_1_3 .LUT_INIT=16'b1000110011001100;
    LogicCell40 \HDA_STRAP.count_17_LC_2_1_3  (
            .in0(N__15023),
            .in1(N__14584),
            .in2(N__14951),
            .in3(N__14710),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34195),
            .ce(N__34688),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_2_1_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI4CB61_17_LC_2_1_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \HDA_STRAP.count_RNI4CB61_17_LC_2_1_4  (
            .in0(N__14502),
            .in1(N__14575),
            .in2(N__14563),
            .in3(N__14538),
            .lcout(),
            .ltout(\HDA_STRAP.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_2_1_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIH7IR1_10_LC_2_1_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \HDA_STRAP.count_RNIH7IR1_10_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(N__14730),
            .in2(N__14527),
            .in3(N__14484),
            .lcout(\HDA_STRAP.un4_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_2_1_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_2_1_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_2_1_6 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \HDA_STRAP.count_16_LC_2_1_6  (
            .in0(N__14708),
            .in1(N__14937),
            .in2(N__14518),
            .in3(N__15027),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34195),
            .ce(N__34688),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_2_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_2_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_2_1_7 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \HDA_STRAP.count_10_LC_2_1_7  (
            .in0(N__14936),
            .in1(N__14491),
            .in2(N__15028),
            .in3(N__14709),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34195),
            .ce(N__34688),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_2_2_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIBJB61_7_LC_2_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \HDA_STRAP.count_RNIBJB61_7_LC_2_2_0  (
            .in0(N__14472),
            .in1(N__14460),
            .in2(N__14449),
            .in3(N__14433),
            .lcout(\HDA_STRAP.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_2_2_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDLB61_6_LC_2_2_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \HDA_STRAP.count_RNIDLB61_6_LC_2_2_1  (
            .in0(N__14808),
            .in1(N__14748),
            .in2(N__14797),
            .in3(N__14766),
            .lcout(\HDA_STRAP.un4_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_2_2_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_2_2_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_2_2_2 .LUT_INIT=16'b1000110011001100;
    LogicCell40 \HDA_STRAP.count_6_LC_2_2_2  (
            .in0(N__15019),
            .in1(N__14773),
            .in2(N__14953),
            .in3(N__14715),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34388),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_2_2_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_2_2_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_2_2_3 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \HDA_STRAP.count_8_LC_2_2_3  (
            .in0(N__14713),
            .in1(N__14755),
            .in2(N__14950),
            .in3(N__15021),
            .lcout(\HDA_STRAP.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34388),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_2_2_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_2_2_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_2_2_4 .LUT_INIT=16'b1000110011001100;
    LogicCell40 \HDA_STRAP.count_11_LC_2_2_4  (
            .in0(N__15018),
            .in1(N__14737),
            .in2(N__14952),
            .in3(N__14714),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34388),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_2_2_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_2_2_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_2_2_5 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_2_2_5  (
            .in0(N__14712),
            .in1(N__15020),
            .in2(N__14949),
            .in3(N__18764),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34388),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_1_2_LC_2_2_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_1_2_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_1_2_LC_2_2_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_1_2_LC_2_2_6  (
            .in0(N__15017),
            .in1(N__14929),
            .in2(_gnd_net_),
            .in3(N__14711),
            .lcout(),
            .ltout(\HDA_STRAP.N_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_2_2_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_2_2_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_2_2_7 .LUT_INIT=16'b0010111000001100;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_2_2_7  (
            .in0(N__15022),
            .in1(N__14676),
            .in2(N__14719),
            .in3(N__14872),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34388),
            .ce(N__34710),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_2_3_0 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_0_LC_2_3_0 .LUT_INIT=16'b1010101000111111;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_0_LC_2_3_0  (
            .in0(N__14716),
            .in1(N__20436),
            .in2(N__31177),
            .in3(N__14923),
            .lcout(\HDA_STRAP.curr_state_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_2_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_2_3_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_2_3_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_2_3_2  (
            .in0(N__15016),
            .in1(N__14677),
            .in2(_gnd_net_),
            .in3(N__14928),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34322),
            .ce(N__34706),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_1_0_LC_2_3_3 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_1_0_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_1_0_LC_2_3_3 .LUT_INIT=16'b0111111101110000;
    LogicCell40 \HDA_STRAP.curr_state_RNO_1_0_LC_2_3_3  (
            .in0(N__20437),
            .in1(N__31176),
            .in2(N__14948),
            .in3(N__15040),
            .lcout(),
            .ltout(\HDA_STRAP.curr_state_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_2_3_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_2_3_4 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_2_3_4  (
            .in0(_gnd_net_),
            .in1(N__15015),
            .in2(N__14962),
            .in3(N__14959),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34322),
            .ce(N__34706),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_2_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNO_0_2_LC_2_3_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \HDA_STRAP.curr_state_RNO_0_2_LC_2_3_6  (
            .in0(_gnd_net_),
            .in1(N__14924),
            .in2(_gnd_net_),
            .in3(N__18753),
            .lcout(\HDA_STRAP.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_2_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_2_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_2_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25620),
            .lcout(\POWERLED.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34390),
            .ce(N__25596),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_2_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_2_4_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_2_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_5_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25755),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34390),
            .ce(N__25596),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_2_4_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_2_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_6_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25689),
            .lcout(\POWERLED.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34390),
            .ce(N__25596),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_2_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_2_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_8_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19015),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34390),
            .ce(N__25596),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_5_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_5_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_5_1  (
            .in0(N__14865),
            .in1(N__14853),
            .in2(N__14842),
            .in3(N__14823),
            .lcout(),
            .ltout(\DSW_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_5_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_2_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIB8TE4_0_LC_2_5_2  (
            .in0(N__15157),
            .in1(N__15214),
            .in2(N__14812),
            .in3(N__16501),
            .lcout(\DSW_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_2_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_2_5_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__21300),
            .in2(_gnd_net_),
            .in3(N__21805),
            .lcout(\POWERLED.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_2_5_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_2_5_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIH71P_2_LC_2_5_4  (
            .in0(N__15264),
            .in1(N__15252),
            .in2(N__15241),
            .in3(N__15225),
            .lcout(\DSW_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_5_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_5_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_2_6_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_2_6_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DSW_PWRGD.count_RNIBCB91_0_LC_2_6_0  (
            .in0(N__15207),
            .in1(N__15195),
            .in2(N__15184),
            .in3(N__15168),
            .lcout(\DSW_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.DSW_PWROK_LC_2_6_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.DSW_PWROK_LC_2_6_1 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_LC_2_6_1  (
            .in0(N__15134),
            .in1(N__15111),
            .in2(N__15088),
            .in3(_gnd_net_),
            .lcout(dsw_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(N__34713),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_2_6_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_2_6_2 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \DSW_PWRGD.curr_state_RNIADII_0_LC_2_6_2  (
            .in0(N__15116),
            .in1(N__15075),
            .in2(_gnd_net_),
            .in3(N__15132),
            .lcout(\DSW_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_0_LC_2_6_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_0_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_0_LC_2_6_3 .LUT_INIT=16'b0100101001000000;
    LogicCell40 \DSW_PWRGD.curr_state_0_LC_2_6_3  (
            .in0(N__15135),
            .in1(N__15112),
            .in2(N__15087),
            .in3(N__15054),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(N__34713),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_1_LC_2_6_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_1_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_1_LC_2_6_4 .LUT_INIT=16'b0001000101010000;
    LogicCell40 \DSW_PWRGD.curr_state_1_LC_2_6_4  (
            .in0(N__15085),
            .in1(N__15058),
            .in2(N__15118),
            .in3(N__15136),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34439),
            .ce(N__34713),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_6_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_6_5 .LUT_INIT=16'b1111000111111011;
    LogicCell40 \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_6_5  (
            .in0(N__15133),
            .in1(N__15117),
            .in2(N__15086),
            .in3(N__15053),
            .lcout(),
            .ltout(DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_27_LC_2_6_6 .C_ON=1'b0;
    defparam \POWERLED.G_27_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_27_LC_2_6_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \POWERLED.G_27_LC_2_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15334),
            .in3(N__34841),
            .lcout(G_27),
            .ltout(G_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_2_6_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_2_6_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \DSW_PWRGD.count_esr_RNO_0_15_LC_2_6_7  (
            .in0(N__34842),
            .in1(_gnd_net_),
            .in2(N__15295),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.N_29_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_9_LC_2_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_2_7_0 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_9_LC_2_7_0  (
            .in0(N__21125),
            .in1(N__20968),
            .in2(_gnd_net_),
            .in3(N__20809),
            .lcout(),
            .ltout(\POWERLED.d_i1_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_16_9_LC_2_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_16_9_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_16_9_LC_2_7_1 .LUT_INIT=16'b1000100000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_16_9_LC_2_7_1  (
            .in0(N__19314),
            .in1(N__16489),
            .in2(N__15283),
            .in3(N__15273),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_16Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_2_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_2_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_2_7_2  (
            .in0(N__21568),
            .in1(N__20811),
            .in2(N__15280),
            .in3(N__21949),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_9_LC_2_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_9_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_9_LC_2_7_3 .LUT_INIT=16'b0001000000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_9_LC_2_7_3  (
            .in0(N__20808),
            .in1(N__21124),
            .in2(N__20971),
            .in3(N__27160),
            .lcout(\POWERLED.un1_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_9_LC_2_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_2_7_4 .LUT_INIT=16'b0011010011010011;
    LogicCell40 \POWERLED.dutycycle_RNI_5_9_LC_2_7_4  (
            .in0(N__27161),
            .in1(N__20969),
            .in2(N__21137),
            .in3(N__20810),
            .lcout(),
            .ltout(\POWERLED.d_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_2_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_2_7_5 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_2_7_5  (
            .in0(N__23278),
            .in1(N__16653),
            .in2(N__15277),
            .in3(N__15274),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_2_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_2_7_6 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_2_7_6  (
            .in0(N__22140),
            .in1(N__21777),
            .in2(N__23797),
            .in3(N__26599),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_0_LC_2_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_2_7_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.dutycycle_RNI_1_0_LC_2_7_7  (
            .in0(N__21776),
            .in1(N__22139),
            .in2(_gnd_net_),
            .in3(N__22383),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_LC_2_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_LC_2_8_0 .LUT_INIT=16'b1100001110000111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_LC_2_8_0  (
            .in0(N__21802),
            .in1(N__22141),
            .in2(N__15346),
            .in3(N__26604),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_2_LC_2_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_2_8_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_2_LC_2_8_1  (
            .in0(N__23792),
            .in1(_gnd_net_),
            .in2(N__15349),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_2_LC_2_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_2_8_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \POWERLED.dutycycle_RNI_1_2_LC_2_8_2  (
            .in0(N__21296),
            .in1(N__23791),
            .in2(_gnd_net_),
            .in3(N__27117),
            .lcout(\POWERLED.un1_dutycycle_53_axb_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_9_LC_2_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_2_8_3 .LUT_INIT=16'b1110101010101000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_9_LC_2_8_3  (
            .in0(N__27118),
            .in1(N__20815),
            .in2(N__16654),
            .in3(N__21129),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_LC_2_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_2_8_4 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_2_8_4  (
            .in0(N__21130),
            .in1(N__20937),
            .in2(N__15337),
            .in3(N__21451),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_0_LC_2_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_2_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_0_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__21298),
            .in2(_gnd_net_),
            .in3(N__22382),
            .lcout(\POWERLED.mult1_un145_sum ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_10_LC_2_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_2_8_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_10_LC_2_8_6  (
            .in0(N__20938),
            .in1(N__21955),
            .in2(_gnd_net_),
            .in3(N__27119),
            .lcout(\POWERLED.g0_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_3_LC_2_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_2_8_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.dutycycle_RNI_7_3_LC_2_8_7  (
            .in0(N__21131),
            .in1(N__21803),
            .in2(_gnd_net_),
            .in3(N__21297),
            .lcout(\POWERLED.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_2_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_9_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15772),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34445),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIJKSP_10_LC_2_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIJKSP_10_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIJKSP_10_LC_2_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNIJKSP_10_LC_2_9_2  (
            .in0(N__15559),
            .in1(N__15502),
            .in2(_gnd_net_),
            .in3(N__30604),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_2_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_2_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_10_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15558),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34445),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNISEFN_2_LC_2_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNISEFN_2_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNISEFN_2_LC_2_9_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNISEFN_2_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__15496),
            .in2(N__15403),
            .in3(N__30603),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_2_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_2_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_2_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15402),
            .lcout(\POWERLED.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34445),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNISF4O_11_LC_2_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNISF4O_11_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNISF4O_11_LC_2_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNISF4O_11_LC_2_9_6  (
            .in0(N__15517),
            .in1(N__15490),
            .in2(_gnd_net_),
            .in3(N__30605),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_2_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_11_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15516),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34445),
            .ce(N__30783),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_2_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_2_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__15480),
            .in2(N__15462),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_2_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_2_10_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIB209_LC_2_10_1  (
            .in0(N__15838),
            .in1(N__15422),
            .in2(_gnd_net_),
            .in3(N__15391),
            .lcout(\POWERLED.count_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_2_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_2_10_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIC419_LC_2_10_2  (
            .in0(N__15841),
            .in1(N__15383),
            .in2(_gnd_net_),
            .in3(N__15352),
            .lcout(\POWERLED.count_1_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2 ),
            .carryout(\POWERLED.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_2_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_2_10_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNID629_LC_2_10_3  (
            .in0(N__15837),
            .in1(N__15668),
            .in2(_gnd_net_),
            .in3(N__15637),
            .lcout(\POWERLED.count_1_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3 ),
            .carryout(\POWERLED.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_2_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_2_10_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNIE839_LC_2_10_4  (
            .in0(N__15842),
            .in1(N__15629),
            .in2(_gnd_net_),
            .in3(N__15598),
            .lcout(\POWERLED.count_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_2_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_2_10_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNIFA49_LC_2_10_5  (
            .in0(N__15839),
            .in1(N__15736),
            .in2(_gnd_net_),
            .in3(N__15595),
            .lcout(\POWERLED.count_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_2_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_2_10_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIGC59_LC_2_10_6  (
            .in0(N__15843),
            .in1(N__16072),
            .in2(_gnd_net_),
            .in3(N__15592),
            .lcout(\POWERLED.count_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_2_10_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_2_10_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIHE69_LC_2_10_7  (
            .in0(N__15840),
            .in1(N__16026),
            .in2(_gnd_net_),
            .in3(N__15589),
            .lcout(\POWERLED.count_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_2_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_2_11_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNIIG79_LC_2_11_0  (
            .in0(N__15844),
            .in1(N__15753),
            .in2(_gnd_net_),
            .in3(N__15586),
            .lcout(\POWERLED.count_1_9 ),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_2_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_2_11_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNIJI89_LC_2_11_1  (
            .in0(N__15849),
            .in1(N__15578),
            .in2(_gnd_net_),
            .in3(N__15547),
            .lcout(\POWERLED.count_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_2_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_2_11_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_2_11_2  (
            .in0(N__15846),
            .in1(N__15536),
            .in2(_gnd_net_),
            .in3(N__15505),
            .lcout(\POWERLED.count_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_2_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_2_11_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNISEH7_LC_2_11_3  (
            .in0(N__15848),
            .in1(N__15974),
            .in2(_gnd_net_),
            .in3(N__15946),
            .lcout(\POWERLED.count_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11_cZ0 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_2_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_2_11_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNITGI7_LC_2_11_4  (
            .in0(N__15845),
            .in1(N__15941),
            .in2(_gnd_net_),
            .in3(N__15901),
            .lcout(\POWERLED.count_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_2_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_2_11_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_2_11_5  (
            .in0(N__15847),
            .in1(N__15897),
            .in2(_gnd_net_),
            .in3(N__15859),
            .lcout(\POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13_cZ0 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_2_11_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_2_11_6  (
            .in0(N__15687),
            .in1(N__15850),
            .in2(_gnd_net_),
            .in3(N__15787),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIA4NN_9_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIA4NN_9_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIA4NN_9_LC_2_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNIA4NN_9_LC_2_11_7  (
            .in0(N__30606),
            .in1(N__15784),
            .in2(_gnd_net_),
            .in3(N__15768),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI4RJN_6_LC_2_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI4RJN_6_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI4RJN_6_LC_2_12_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI4RJN_6_LC_2_12_0  (
            .in0(N__15700),
            .in1(N__30600),
            .in2(_gnd_net_),
            .in3(N__15711),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_2_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_2_12_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_6_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15715),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34459),
            .ce(N__30785),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI4S8O_15_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI4S8O_15_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI4S8O_15_LC_2_12_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI4S8O_15_LC_2_12_2  (
            .in0(N__16078),
            .in1(N__30599),
            .in2(_gnd_net_),
            .in3(N__16086),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_2_12_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_15_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16090),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34459),
            .ce(N__30785),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI6UKN_7_LC_2_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI6UKN_7_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI6UKN_7_LC_2_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI6UKN_7_LC_2_12_4  (
            .in0(N__16036),
            .in1(N__30601),
            .in2(_gnd_net_),
            .in3(N__16047),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_2_12_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_7_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16051),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34459),
            .ce(N__30785),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI81MN_8_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI81MN_8_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI81MN_8_LC_2_12_6 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \POWERLED.count_RNI81MN_8_LC_2_12_6  (
            .in0(N__15991),
            .in1(N__30602),
            .in2(N__16006),
            .in3(_gnd_net_),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_2_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_8_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16005),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34459),
            .ce(N__30785),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__19711),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__16873),
            .in2(N__16214),
            .in3(N__15985),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__16126),
            .in2(N__16216),
            .in3(N__15982),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__16117),
            .in2(N__16253),
            .in3(N__15979),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__16108),
            .in2(N__16254),
            .in3(N__16144),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_13_5  (
            .in0(N__16989),
            .in1(N__16099),
            .in2(N__16215),
            .in3(N__16141),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_13_6  (
            .in0(N__16267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16138),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(\POWERLED.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16135),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_2_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_2_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__19672),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_2_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_2_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__16765),
            .in2(N__16350),
            .in3(N__16120),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_2_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_2_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__16346),
            .in2(N__16192),
            .in3(N__16111),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_2_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_2_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__16180),
            .in2(N__16383),
            .in3(N__16102),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_2_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_2_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__16171),
            .in2(N__16384),
            .in3(N__16093),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_2_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_2_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_2_14_5  (
            .in0(N__16243),
            .in1(N__16162),
            .in2(N__16351),
            .in3(N__16261),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_2_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_2_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_2_14_6  (
            .in0(N__16153),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16258),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16242),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__19633),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__16397),
            .in2(N__20092),
            .in3(N__16183),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__16333),
            .in2(N__16402),
            .in3(N__16174),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__16424),
            .in2(N__16324),
            .in3(N__16165),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__16312),
            .in2(N__16429),
            .in3(N__16156),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_2_15_5  (
            .in0(N__16375),
            .in1(N__16401),
            .in2(N__16303),
            .in3(N__16147),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__16276),
            .in2(_gnd_net_),
            .in3(N__16387),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(\POWERLED.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_2_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_2_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16354),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__20116),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__16287),
            .in2(N__20236),
            .in3(N__16327),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2_c ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__17026),
            .in2(N__16291),
            .in3(N__16315),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3_c ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__17353),
            .in2(N__17280),
            .in3(N__16306),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4_c ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__17275),
            .in2(N__17341),
            .in3(N__16294),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5_c ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_16_5  (
            .in0(N__16423),
            .in1(N__16286),
            .in2(N__17326),
            .in3(N__16270),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6_c ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_16_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_16_6  (
            .in0(N__17296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16432),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(\POWERLED.mult1_un96_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16405),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_2_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_4_2_0  (
            .in0(N__17212),
            .in1(N__17192),
            .in2(N__17146),
            .in3(N__17168),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_4_2_1 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_4_2_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_3_LC_4_2_1  (
            .in0(N__17169),
            .in1(N__25096),
            .in2(_gnd_net_),
            .in3(N__17155),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34267),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_4_2_2 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_4_2_2 .LUT_INIT=16'b0000011000000110;
    LogicCell40 \COUNTER.counter_1_LC_4_2_2  (
            .in0(N__17223),
            .in1(N__17241),
            .in2(N__25119),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34267),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_4_2_3 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_4_2_3 .LUT_INIT=16'b0001001000010010;
    LogicCell40 \COUNTER.counter_6_LC_4_2_3  (
            .in0(N__17409),
            .in1(N__25099),
            .in2(N__17395),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34267),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_4_2_4 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_4_2_4 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \COUNTER.counter_2_LC_4_2_4  (
            .in0(N__17179),
            .in1(_gnd_net_),
            .in2(N__25120),
            .in3(N__17193),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34267),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_4_2_5 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_4_2_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_4_LC_4_2_5  (
            .in0(N__17145),
            .in1(N__25097),
            .in2(_gnd_net_),
            .in3(N__17125),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34267),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_4_2_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_4_2_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_4_2_6  (
            .in0(N__17382),
            .in1(N__17408),
            .in2(N__17440),
            .in3(N__17240),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_4_2_7 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_4_2_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_5_LC_4_2_7  (
            .in0(N__17439),
            .in1(N__25098),
            .in2(_gnd_net_),
            .in3(N__17419),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34267),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI94A94_LC_4_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI94A94_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI94A94_LC_4_3_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI94A94_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__20430),
            .in2(_gnd_net_),
            .in3(N__31166),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_4_3_5 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_4_3_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_4_3_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \COUNTER.counter_0_LC_4_3_5  (
            .in0(_gnd_net_),
            .in1(N__25106),
            .in2(_gnd_net_),
            .in3(N__17219),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34321),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIV3O1A_4_LC_4_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIV3O1A_4_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIV3O1A_4_LC_4_4_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.count_off_RNIV3O1A_4_LC_4_4_0  (
            .in0(N__26918),
            .in1(N__16459),
            .in2(N__25591),
            .in3(N__19074),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_4_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_4_4_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_3_LC_4_4_1  (
            .in0(N__19105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26920),
            .lcout(\POWERLED.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34271),
            .ce(N__25597),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_4_4_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_4_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_4_LC_4_4_2  (
            .in0(N__26919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19075),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34271),
            .ce(N__25597),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI7GS1A_8_LC_4_4_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI7GS1A_8_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI7GS1A_8_LC_4_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNI7GS1A_8_LC_4_4_3  (
            .in0(N__16453),
            .in1(N__19011),
            .in2(_gnd_net_),
            .in3(N__25579),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(\POWERLED.count_offZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_3_LC_4_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_3_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_3_LC_4_4_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_3_LC_4_4_4  (
            .in0(N__19119),
            .in1(N__19053),
            .in2(N__16444),
            .in3(N__19090),
            .lcout(\POWERLED.un34_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIT0N1A_3_LC_4_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIT0N1A_3_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIT0N1A_3_LC_4_4_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \POWERLED.count_off_RNIT0N1A_3_LC_4_4_5  (
            .in0(N__19104),
            .in1(N__25574),
            .in2(N__16441),
            .in3(N__26917),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_4_4_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_4_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_7_LC_4_4_6  (
            .in0(N__19039),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34271),
            .ce(N__25597),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI5DR1A_7_LC_4_4_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI5DR1A_7_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI5DR1A_7_LC_4_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNI5DR1A_7_LC_4_4_7  (
            .in0(N__16573),
            .in1(N__19038),
            .in2(_gnd_net_),
            .in3(N__25578),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_4_5_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_4_5_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_RNIKA1P_1_LC_4_5_1  (
            .in0(N__16567),
            .in1(N__16552),
            .in2(N__16537),
            .in3(N__16516),
            .lcout(\DSW_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_4_5_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_4_5_2 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_4_5_2  (
            .in0(N__21105),
            .in1(_gnd_net_),
            .in2(N__21278),
            .in3(N__21766),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_4_5_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_4_5_3 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_4_5_3  (
            .in0(N__20942),
            .in1(N__21796),
            .in2(N__16492),
            .in3(N__26603),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_4_5_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_4_5_4 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_4_5_4  (
            .in0(N__21241),
            .in1(N__21762),
            .in2(_gnd_net_),
            .in3(N__20940),
            .lcout(\POWERLED.un1_dutycycle_53_20_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_4_5_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_4_5_5 .LUT_INIT=16'b0000011100011111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_4_5_5  (
            .in0(N__20941),
            .in1(N__21242),
            .in2(N__21801),
            .in3(N__21104),
            .lcout(),
            .ltout(\POWERLED.o2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_9_LC_4_5_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_4_5_6 .LUT_INIT=16'b0111011100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_9_LC_4_5_6  (
            .in0(N__19297),
            .in1(N__16482),
            .in2(N__16471),
            .in3(N__20805),
            .lcout(\POWERLED.un1_dutycycle_53_axb_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_4_5_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_4_5_7 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_4_5_7  (
            .in0(N__20939),
            .in1(N__21240),
            .in2(N__21800),
            .in3(N__21103),
            .lcout(\POWERLED.un1_dutycycle_53_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_9_LC_4_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_4_6_0 .LUT_INIT=16'b1010100110100110;
    LogicCell40 \POWERLED.dutycycle_RNI_0_9_LC_4_6_0  (
            .in0(N__16594),
            .in1(N__20806),
            .in2(N__16468),
            .in3(N__27152),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_10_LC_4_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_4_6_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_10_LC_4_6_1  (
            .in0(N__21900),
            .in1(_gnd_net_),
            .in2(N__16600),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_4_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_4_6_2 .LUT_INIT=16'b1110110011001000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_4_6_2  (
            .in0(N__21062),
            .in1(N__21728),
            .in2(N__21279),
            .in3(N__20949),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_3 ),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_9_LC_4_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_4_6_3 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_9_LC_4_6_3  (
            .in0(N__20807),
            .in1(N__27151),
            .in2(N__16597),
            .in3(N__26602),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_10_LC_4_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_4_6_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_10_LC_4_6_4  (
            .in0(N__21063),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21896),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_1_LC_4_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_4_6_5 .LUT_INIT=16'b0000111101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_1_LC_4_6_5  (
            .in0(N__21729),
            .in1(_gnd_net_),
            .in2(N__22145),
            .in3(N__26601),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_4_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_4_6_6 .LUT_INIT=16'b1010111100001010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_4_6_6  (
            .in0(N__21249),
            .in1(N__19732),
            .in2(N__16588),
            .in3(N__27153),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_4_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_4_6_7 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_4_6_7  (
            .in0(N__20950),
            .in1(_gnd_net_),
            .in2(N__21926),
            .in3(N__21064),
            .lcout(\POWERLED.un1_dutycycle_53_8_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_11_LC_4_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_4_7_0 .LUT_INIT=16'b0000101000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_3_11_LC_4_7_0  (
            .in0(N__16585),
            .in1(N__21385),
            .in2(N__21450),
            .in3(N__23265),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_11_LC_4_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_11_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_11_LC_4_7_1 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_11_LC_4_7_1  (
            .in0(N__16639),
            .in1(N__16612),
            .in2(N__16579),
            .in3(N__16660),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_8_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_4_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_4_7_2 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_4_7_2  (
            .in0(N__21566),
            .in1(N__16618),
            .in2(N__16576),
            .in3(N__27142),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_4_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_4_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_4_7_3  (
            .in0(N__21102),
            .in1(N__21892),
            .in2(N__23273),
            .in3(N__20920),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_3Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_4_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_4_7_4 .LUT_INIT=16'b0000011100001110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_4_7_4  (
            .in0(N__21894),
            .in1(N__20776),
            .in2(N__16663),
            .in3(N__23261),
            .lcout(\POWERLED.un1_dutycycle_53_8_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_4_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_4_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_4_7_5  (
            .in0(N__16640),
            .in1(N__20924),
            .in2(N__23274),
            .in3(N__21895),
            .lcout(\POWERLED.un1_dutycycle_53_56_a0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_4_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_4_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_4_7_6  (
            .in0(N__21893),
            .in1(N__27141),
            .in2(N__20951),
            .in3(N__23260),
            .lcout(\POWERLED.un1_dutycycle_53_56_a1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_9_LC_4_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_4_7_7 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_9_LC_4_7_7  (
            .in0(N__20775),
            .in1(N__20919),
            .in2(N__21388),
            .in3(N__21891),
            .lcout(\POWERLED.un1_dutycycle_53_50_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_4_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_4_8_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_4_8_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \POWERLED.dutycycle_8_LC_4_8_0  (
            .in0(N__16696),
            .in1(N__20830),
            .in2(N__29811),
            .in3(N__16690),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34368),
            .ce(),
            .sr(N__23685));
    defparam \POWERLED.dutycycle_RNI2O4A1_13_LC_4_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_13_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_13_LC_4_8_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_13_LC_4_8_1  (
            .in0(N__26049),
            .in1(N__21555),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_45_and_i_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5MDM4_13_LC_4_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5MDM4_13_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5MDM4_13_LC_4_8_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI5MDM4_13_LC_4_8_2  (
            .in0(N__23372),
            .in1(N__25861),
            .in2(N__16606),
            .in3(N__23464),
            .lcout(),
            .ltout(\POWERLED.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRBF58_13_LC_4_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRBF58_13_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRBF58_13_LC_4_8_3 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \POWERLED.dutycycle_RNIRBF58_13_LC_4_8_3  (
            .in0(N__26767),
            .in1(N__29774),
            .in2(N__16603),
            .in3(N__23073),
            .lcout(\POWERLED.dutycycle_en_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3U8C3_8_LC_4_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3U8C3_8_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3U8C3_8_LC_4_8_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI3U8C3_8_LC_4_8_4  (
            .in0(N__23371),
            .in1(N__26048),
            .in2(N__25872),
            .in3(N__20913),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQN4F7_8_LC_4_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQN4F7_8_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQN4F7_8_LC_4_8_5 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \POWERLED.dutycycle_RNIQN4F7_8_LC_4_8_5  (
            .in0(N__23463),
            .in1(N__26765),
            .in2(N__16699),
            .in3(N__23072),
            .lcout(\POWERLED.dutycycle_eena_3 ),
            .ltout(\POWERLED.dutycycle_eena_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITTBN9_8_LC_4_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITTBN9_8_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITTBN9_8_LC_4_8_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNITTBN9_8_LC_4_8_6  (
            .in0(N__29773),
            .in1(N__16689),
            .in2(N__16678),
            .in3(N__20829),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(\POWERLED.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_10_LC_4_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_4_8_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.dutycycle_RNI_4_10_LC_4_8_7  (
            .in0(N__21925),
            .in1(_gnd_net_),
            .in2(N__16675),
            .in3(N__21061),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_9_LC_4_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_9_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_9_LC_4_9_1 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_9_LC_4_9_1  (
            .in0(N__20931),
            .in1(N__20812),
            .in2(N__21387),
            .in3(N__21106),
            .lcout(\POWERLED.un1_dutycycle_53_4_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_4_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_4_9_2 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__21380),
            .in2(N__21951),
            .in3(N__23247),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_4_9_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_4_9_3 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_4_9_3  (
            .in0(N__20932),
            .in1(N__19315),
            .in2(N__16672),
            .in3(N__16669),
            .lcout(\POWERLED.un1_dutycycle_53_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__17754),
            .in2(_gnd_net_),
            .in3(N__17907),
            .lcout(\POWERLED.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_14_LC_4_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_4_9_5 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_14_LC_4_9_5  (
            .in0(N__21381),
            .in1(_gnd_net_),
            .in2(N__23268),
            .in3(N__25376),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_13_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_4_9_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_13_LC_4_9_6  (
            .in0(N__20813),
            .in1(N__21567),
            .in2(N__16729),
            .in3(N__25405),
            .lcout(\POWERLED.un2_count_clk_17_0_a2_5 ),
            .ltout(\POWERLED.un2_count_clk_17_0_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_3_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_4_9_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_3_LC_4_9_7  (
            .in0(N__20933),
            .in1(N__21307),
            .in2(N__16726),
            .in3(N__21107),
            .lcout(\POWERLED.m18_e_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19771),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16774),
            .in3(N__16723),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__16705),
            .in2(N__17707),
            .in3(N__16720),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__34556),
            .in2(N__17686),
            .in3(N__16717),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__34561),
            .in2(N__17923),
            .in3(N__16714),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_4_10_5  (
            .in0(N__18214),
            .in1(N__18004),
            .in2(N__17986),
            .in3(N__16711),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_10_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(N__17908),
            .in2(N__17758),
            .in3(N__16708),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_10_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_4_10_7  (
            .in0(N__17702),
            .in1(N__17703),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.slp_s3n_signal_i_LC_4_11_1 .C_ON=1'b0;
    defparam \POWERLED.slp_s3n_signal_i_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.slp_s3n_signal_i_LC_4_11_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.slp_s3n_signal_i_LC_4_11_1  (
            .in0(N__27340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26412),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19882),
            .lcout(\POWERLED.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_4_11_4  (
            .in0(N__22147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_4_11_6  (
            .in0(N__19632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_SUSn_RNIN4K9_LC_4_11_7.C_ON=1'b0;
    defparam SLP_SUSn_RNIN4K9_LC_4_11_7.SEQ_MODE=4'b0000;
    defparam SLP_SUSn_RNIN4K9_LC_4_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 SLP_SUSn_RNIN4K9_LC_4_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24886),
            .lcout(v33a_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_4_12_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_4_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_4_12_0  (
            .in0(N__17103),
            .in1(N__16935),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_12_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19389),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_4_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_4_12_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_4_12_2  (
            .in0(N__17102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_4_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_4_12_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__17104),
            .in2(_gnd_net_),
            .in3(N__16887),
            .lcout(\POWERLED.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_10_LC_4_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_4_12_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_10_LC_4_12_4  (
            .in0(N__20943),
            .in1(N__24114),
            .in2(N__19943),
            .in3(N__21952),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_12_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19707),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19671),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__19390),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__16973),
            .in2(N__16861),
            .in3(N__16852),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__16849),
            .in2(N__16978),
            .in3(N__16840),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__16837),
            .in2(N__17002),
            .in3(N__16828),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__17001),
            .in2(N__16825),
            .in3(N__16813),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_4_13_5  (
            .in0(N__17101),
            .in1(N__16977),
            .in2(N__16810),
            .in3(N__16798),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_4_13_6  (
            .in0(N__17014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17005),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_4_13_7  (
            .in0(N__16997),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__20290),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__17077),
            .in2(N__16963),
            .in3(N__16951),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(N__16948),
            .in2(N__16939),
            .in3(N__16924),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(N__17106),
            .in2(N__16921),
            .in3(N__16912),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_14_4  (
            .in0(_gnd_net_),
            .in1(N__16909),
            .in2(N__17110),
            .in3(N__16903),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_14_5  (
            .in0(N__18465),
            .in1(N__16900),
            .in2(N__16891),
            .in3(N__16876),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_14_6  (
            .in0(N__17119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17113),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17105),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_4_15_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_4_15_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_4_15_1  (
            .in0(N__19558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18251),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_4_15_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_4_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(N__30213),
            .in2(_gnd_net_),
            .in3(N__17071),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18553),
            .lcout(\POWERLED.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_15_7  (
            .in0(N__18466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_4_16_0  (
            .in0(_gnd_net_),
            .in1(N__20257),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_16_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__17309),
            .in2(N__17035),
            .in3(N__17017),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_4_16_2  (
            .in0(_gnd_net_),
            .in1(N__17311),
            .in2(N__18379),
            .in3(N__17344),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_4_16_3  (
            .in0(_gnd_net_),
            .in1(N__18355),
            .in2(N__18267),
            .in3(N__17329),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_4_16_4  (
            .in0(_gnd_net_),
            .in1(N__18263),
            .in2(N__18334),
            .in3(N__17314),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_16_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_4_16_5  (
            .in0(N__17260),
            .in1(N__17310),
            .in2(N__18313),
            .in3(N__17287),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_16_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_4_16_6  (
            .in0(_gnd_net_),
            .in1(N__18289),
            .in2(_gnd_net_),
            .in3(N__17284),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_5_1_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_5_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_5_1_0  (
            .in0(_gnd_net_),
            .in1(N__17242),
            .in2(N__17227),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_1_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_1_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__17194),
            .in2(_gnd_net_),
            .in3(N__17173),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_1_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(N__17170),
            .in2(_gnd_net_),
            .in3(N__17149),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_1_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_1_3  (
            .in0(_gnd_net_),
            .in1(N__17144),
            .in2(_gnd_net_),
            .in3(N__17443),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_1_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_1_4  (
            .in0(_gnd_net_),
            .in1(N__17438),
            .in2(_gnd_net_),
            .in3(N__17413),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_1_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_1_5  (
            .in0(_gnd_net_),
            .in1(N__17410),
            .in2(_gnd_net_),
            .in3(N__17386),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_5_1_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_5_1_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_5_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(N__17383),
            .in2(_gnd_net_),
            .in3(N__17371),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__34020),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_5_1_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_5_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_5_1_7  (
            .in0(_gnd_net_),
            .in1(N__18697),
            .in2(_gnd_net_),
            .in3(N__17368),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__34020),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_5_2_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_5_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__18672),
            .in2(_gnd_net_),
            .in3(N__17365),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_5_2_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_5_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__18685),
            .in2(_gnd_net_),
            .in3(N__17362),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_5_2_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_5_2_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_5_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__18658),
            .in2(_gnd_net_),
            .in3(N__17359),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_5_2_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_5_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__18621),
            .in2(_gnd_net_),
            .in3(N__17356),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_5_2_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_5_2_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_5_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__18634),
            .in2(_gnd_net_),
            .in3(N__17470),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_5_2_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_5_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__18646),
            .in2(_gnd_net_),
            .in3(N__17467),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_5_2_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_5_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__18607),
            .in2(_gnd_net_),
            .in3(N__17464),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_5_2_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_5_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__18841),
            .in2(_gnd_net_),
            .in3(N__17461),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__34163),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_5_3_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_5_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__18802),
            .in2(_gnd_net_),
            .in3(N__17458),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_5_3_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_5_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__18829),
            .in2(_gnd_net_),
            .in3(N__17455),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_5_3_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_5_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__18816),
            .in2(_gnd_net_),
            .in3(N__17452),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_5_3_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_5_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__18922),
            .in2(_gnd_net_),
            .in3(N__17449),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_5_3_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_5_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(N__18936),
            .in2(_gnd_net_),
            .in3(N__17446),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_5_3_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_5_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__18949),
            .in2(_gnd_net_),
            .in3(N__17497),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_5_3_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_5_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(N__18961),
            .in2(_gnd_net_),
            .in3(N__17494),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_5_3_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_5_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(N__18901),
            .in2(_gnd_net_),
            .in3(N__17491),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__34185),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_5_4_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_5_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__18862),
            .in2(_gnd_net_),
            .in3(N__17488),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_5_4_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_5_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__18876),
            .in2(_gnd_net_),
            .in3(N__17485),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_5_4_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_5_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__18889),
            .in2(_gnd_net_),
            .in3(N__17482),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_5_4_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_5_4_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_28_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17566),
            .in3(N__17479),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_5_4_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_5_4_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_29_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17530),
            .in3(N__17476),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_5_4_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_5_4_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_30_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17545),
            .in3(N__17473),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_5_4_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_5_4_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.counter_31_LC_5_4_6  (
            .in0(N__17554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17569),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_5_4_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_5_4_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_5_4_7  (
            .in0(N__17562),
            .in1(N__17553),
            .in2(N__17544),
            .in3(N__17526),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_5_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_5_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_9_LC_5_5_0  (
            .in0(N__18988),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34196),
            .ce(N__25590),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI9JT1A_9_LC_5_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI9JT1A_9_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI9JT1A_9_LC_5_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNI9JT1A_9_LC_5_5_1  (
            .in0(N__17518),
            .in1(N__25550),
            .in2(_gnd_net_),
            .in3(N__18987),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(\POWERLED.count_offZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_10_LC_5_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_10_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_10_LC_5_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_10_LC_5_5_2  (
            .in0(N__19189),
            .in1(N__19215),
            .in2(N__17512),
            .in3(N__19165),
            .lcout(\POWERLED.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIIT20A_10_LC_5_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIIT20A_10_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIIT20A_10_LC_5_5_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIIT20A_10_LC_5_5_3  (
            .in0(N__17509),
            .in1(N__25551),
            .in2(_gnd_net_),
            .in3(N__19200),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_5_5_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_5_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_10_LC_5_5_4  (
            .in0(N__19201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34196),
            .ce(N__25590),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIR4GU9_11_LC_5_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIR4GU9_11_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIR4GU9_11_LC_5_5_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIR4GU9_11_LC_5_5_5  (
            .in0(N__17503),
            .in1(N__25552),
            .in2(_gnd_net_),
            .in3(N__19176),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_5_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_5_5_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_11_LC_5_5_6  (
            .in0(N__19177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34196),
            .ce(N__25590),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIT7HU9_12_LC_5_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIT7HU9_12_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIT7HU9_12_LC_5_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIT7HU9_12_LC_5_5_7  (
            .in0(N__19129),
            .in1(N__25553),
            .in2(_gnd_net_),
            .in3(N__19140),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3U8C3_3_LC_5_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3U8C3_3_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3U8C3_3_LC_5_6_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI3U8C3_3_LC_5_6_0  (
            .in0(N__26047),
            .in1(N__25865),
            .in2(N__23380),
            .in3(N__21267),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQN4F7_3_LC_5_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQN4F7_3_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQN4F7_3_LC_5_6_1 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \POWERLED.dutycycle_RNIQN4F7_3_LC_5_6_1  (
            .in0(N__23070),
            .in1(N__26770),
            .in2(N__17617),
            .in3(N__23459),
            .lcout(\POWERLED.dutycycle_eena_8 ),
            .ltout(\POWERLED.dutycycle_eena_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJE6N9_3_LC_5_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJE6N9_3_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJE6N9_3_LC_5_6_2 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_RNIJE6N9_3_LC_5_6_2  (
            .in0(N__21184),
            .in1(N__29821),
            .in2(N__17614),
            .in3(N__17604),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_5_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_5_6_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_5_6_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_3_LC_5_6_3  (
            .in0(N__17605),
            .in1(N__17611),
            .in2(N__29830),
            .in3(N__21183),
            .lcout(\POWERLED.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34349),
            .ce(),
            .sr(N__23698));
    defparam \POWERLED.dutycycle_RNI8U6P9_10_LC_5_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8U6P9_10_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8U6P9_10_LC_5_6_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_RNI8U6P9_10_LC_5_6_4  (
            .in0(N__17577),
            .in1(N__29820),
            .in2(N__17590),
            .in3(N__20682),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(\POWERLED.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3U8C3_10_LC_5_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3U8C3_10_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3U8C3_10_LC_5_6_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI3U8C3_10_LC_5_6_5  (
            .in0(N__25864),
            .in1(N__23376),
            .in2(N__17596),
            .in3(N__26046),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQN4F7_10_LC_5_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQN4F7_10_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQN4F7_10_LC_5_6_6 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \POWERLED.dutycycle_RNIQN4F7_10_LC_5_6_6  (
            .in0(N__26769),
            .in1(N__23458),
            .in2(N__17593),
            .in3(N__23069),
            .lcout(\POWERLED.dutycycle_eena_4 ),
            .ltout(\POWERLED.dutycycle_eena_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_5_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_5_6_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_5_6_7 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_10_LC_5_6_7  (
            .in0(N__20683),
            .in1(N__29825),
            .in2(N__17581),
            .in3(N__17578),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34349),
            .ce(),
            .sr(N__23698));
    defparam \POWERLED.dutycycle_RNIQN4F7_7_LC_5_7_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQN4F7_7_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQN4F7_7_LC_5_7_0 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \POWERLED.dutycycle_RNIQN4F7_7_LC_5_7_0  (
            .in0(N__26741),
            .in1(N__23460),
            .in2(N__23074),
            .in3(N__17668),
            .lcout(\POWERLED.dutycycle_eena_5 ),
            .ltout(\POWERLED.dutycycle_eena_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNII46M9_7_LC_5_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNII46M9_7_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNII46M9_7_LC_5_7_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_RNII46M9_7_LC_5_7_1  (
            .in0(N__29812),
            .in1(N__17628),
            .in2(N__17674),
            .in3(N__20985),
            .lcout(\POWERLED.dutycycleZ1Z_5 ),
            .ltout(\POWERLED.dutycycleZ1Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3U8C3_7_LC_5_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3U8C3_7_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3U8C3_7_LC_5_7_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI3U8C3_7_LC_5_7_2  (
            .in0(N__25862),
            .in1(N__23374),
            .in2(N__17671),
            .in3(N__26036),
            .lcout(\POWERLED.dutycycle_eena_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILH7N9_4_LC_5_7_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILH7N9_4_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILH7N9_4_LC_5_7_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_RNILH7N9_4_LC_5_7_3  (
            .in0(N__17646),
            .in1(N__17656),
            .in2(N__29828),
            .in3(N__21166),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3U8C3_4_LC_5_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3U8C3_4_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3U8C3_4_LC_5_7_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI3U8C3_4_LC_5_7_4  (
            .in0(N__25863),
            .in1(N__23375),
            .in2(N__17662),
            .in3(N__26037),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQN4F7_4_LC_5_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQN4F7_4_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQN4F7_4_LC_5_7_5 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \POWERLED.dutycycle_RNIQN4F7_4_LC_5_7_5  (
            .in0(N__23461),
            .in1(N__26742),
            .in2(N__17659),
            .in3(N__23068),
            .lcout(\POWERLED.dutycycle_eena_6 ),
            .ltout(\POWERLED.dutycycle_eena_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_5_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_5_7_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_5_7_6 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_4_LC_5_7_6  (
            .in0(N__17647),
            .in1(N__29816),
            .in2(N__17650),
            .in3(N__21162),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34323),
            .ce(),
            .sr(N__23696));
    defparam \POWERLED.dutycycle_7_LC_5_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_5_7_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_5_7_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \POWERLED.dutycycle_7_LC_5_7_7  (
            .in0(N__17635),
            .in1(N__20986),
            .in2(N__29829),
            .in3(N__17629),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34323),
            .ce(),
            .sr(N__23696));
    defparam \POWERLED.dutycycle_RNI5MDM4_15_LC_5_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5MDM4_15_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5MDM4_15_LC_5_8_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.dutycycle_RNI5MDM4_15_LC_5_8_0  (
            .in0(N__17740),
            .in1(N__23462),
            .in2(N__25873),
            .in3(N__23373),
            .lcout(),
            .ltout(\POWERLED.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRBF58_15_LC_5_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRBF58_15_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRBF58_15_LC_5_8_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \POWERLED.dutycycle_RNIRBF58_15_LC_5_8_1  (
            .in0(N__26766),
            .in1(N__23071),
            .in2(N__17620),
            .in3(N__29778),
            .lcout(\POWERLED.dutycycle_en_12 ),
            .ltout(\POWERLED.dutycycle_en_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_5_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_5_8_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_5_8_2 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_15_LC_5_8_2  (
            .in0(N__17727),
            .in1(N__29987),
            .in2(N__17743),
            .in3(N__21463),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34223),
            .ce(),
            .sr(N__23670));
    defparam \POWERLED.dutycycle_RNI2O4A1_15_LC_5_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_15_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_15_LC_5_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_15_LC_5_8_3  (
            .in0(N__26050),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25406),
            .lcout(\POWERLED.un1_clk_100khz_48_and_i_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIPUS6A_15_LC_5_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIPUS6A_15_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIPUS6A_15_LC_5_8_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.dutycycle_RNIPUS6A_15_LC_5_8_4  (
            .in0(N__17734),
            .in1(N__29986),
            .in2(N__17728),
            .in3(N__21462),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(\POWERLED.dutycycleZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_5_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_5_8_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17716),
            .in3(N__23267),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_5_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_5_8_6 .LUT_INIT=16'b1110000100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_5_8_6  (
            .in0(N__17767),
            .in1(N__19459),
            .in2(N__17713),
            .in3(N__21434),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_5_8_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17710),
            .in3(N__25407),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19878),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17968),
            .in3(N__17689),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17977),
            .in3(N__17677),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__34537),
            .in2(N__18013),
            .in3(N__17914),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4 .C_ON=1'b0;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17911),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_0_LC_5_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_5_9_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNI_6_0_LC_5_9_5  (
            .in0(N__22146),
            .in1(N__32968),
            .in2(N__22384),
            .in3(N__21109),
            .lcout(\POWERLED.g2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_LC_5_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_5_9_6 .LUT_INIT=16'b1010111101010000;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_5_9_6  (
            .in0(N__19453),
            .in1(N__25378),
            .in2(N__17896),
            .in3(N__21529),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_5_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_5_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_5_9_7  (
            .in0(N__21784),
            .in1(N__21280),
            .in2(_gnd_net_),
            .in3(N__21108),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_5_10_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_5_10_0 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \POWERLED.curr_state_0_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__17887),
            .in2(N__17851),
            .in3(N__17818),
            .lcout(\POWERLED.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34357),
            .ce(N__30782),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_9_LC_5_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_9_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_9_LC_5_10_1 .LUT_INIT=16'b0001000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_9_LC_5_10_1  (
            .in0(N__17776),
            .in1(N__19237),
            .in2(N__20814),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_9Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_2 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_5_10_2  (
            .in0(N__19857),
            .in1(_gnd_net_),
            .in2(N__19816),
            .in3(N__19836),
            .lcout(\POWERLED.mult1_un40_sum_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_3 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__19856),
            .in2(N__19837),
            .in3(N__19812),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_10_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_5_10_5  (
            .in0(N__18002),
            .in1(N__18003),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19858),
            .in3(N__19832),
            .lcout(\POWERLED.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_5_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_5_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19852),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_11_0  (
            .in0(_gnd_net_),
            .in1(N__19794),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__19753),
            .in2(N__18192),
            .in3(N__17959),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_11_2  (
            .in0(_gnd_net_),
            .in1(N__18188),
            .in2(N__17956),
            .in3(N__17947),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__17944),
            .in2(N__18220),
            .in3(N__17938),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__18218),
            .in2(N__17935),
            .in3(N__17926),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_11_5  (
            .in0(N__18070),
            .in1(N__18133),
            .in2(N__18193),
            .in3(N__18127),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18124),
            .in3(N__18115),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(\POWERLED.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18112),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19990),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(N__19783),
            .in2(N__18033),
            .in3(N__18109),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(N__18029),
            .in2(N__18106),
            .in3(N__18097),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__18094),
            .in2(N__18078),
            .in3(N__18088),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__18074),
            .in2(N__18052),
            .in3(N__18043),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_12_5  (
            .in0(N__20212),
            .in1(N__18040),
            .in2(N__18034),
            .in3(N__18016),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__18229),
            .in2(_gnd_net_),
            .in3(N__18223),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18219),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20170),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__18389),
            .in2(N__19972),
            .in3(N__18175),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__18172),
            .in2(N__18394),
            .in3(N__18166),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__18163),
            .in2(N__20221),
            .in3(N__18157),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__18154),
            .in2(N__20220),
            .in3(N__18148),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_13_5  (
            .in0(N__18543),
            .in1(N__18393),
            .in2(N__18145),
            .in3(N__18136),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_13_6  (
            .in0(N__18403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18397),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20213),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__19554),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__18518),
            .in2(N__20152),
            .in3(N__18367),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__18364),
            .in2(N__18523),
            .in3(N__18346),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__18545),
            .in2(N__18343),
            .in3(N__18322),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__18319),
            .in2(N__18552),
            .in3(N__18301),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_14_5  (
            .in0(N__18250),
            .in1(N__18522),
            .in2(N__18298),
            .in3(N__18280),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_14_6  (
            .in0(N__18277),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18271),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18544),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_5_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_5_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__20143),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_5_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__18434),
            .in2(N__20266),
            .in3(N__18508),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_5_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__18505),
            .in2(N__18439),
            .in3(N__18499),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_5_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__18467),
            .in2(N__18496),
            .in3(N__18487),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_5_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__18484),
            .in2(N__18474),
            .in3(N__18442),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_5_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_5_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_5_15_5  (
            .in0(N__20323),
            .in1(N__18438),
            .in2(N__18424),
            .in3(N__18415),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_5_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_5_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_5_15_6  (
            .in0(N__18412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18406),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(\POWERLED.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_15_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18712),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_6_1_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_6_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_6_1_0  (
            .in0(N__18696),
            .in1(N__18684),
            .in2(N__18673),
            .in3(N__18657),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_6_1_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_6_1_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_6_1_1  (
            .in0(N__18645),
            .in1(N__18633),
            .in2(N__18622),
            .in3(N__18606),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_6_2_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_6_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18595),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_6_2_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_6_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18583),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_6_2_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_6_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_6_2_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_6_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18562),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_6_2_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_6_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18790),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_6_2_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_6_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_6_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18910),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_6_2_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_6_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18850),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_6_2_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_6_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18976),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(COUNTER_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_3_0.C_ON=1'b0;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_3_0.SEQ_MODE=4'b0000;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18964),
            .lcout(COUNTER_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_6_3_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_6_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_6_3_2  (
            .in0(N__18960),
            .in1(N__18948),
            .in2(N__18937),
            .in3(N__18921),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_6_3_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_6_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_6_3_3  (
            .in0(N__18900),
            .in1(N__18888),
            .in2(N__18877),
            .in3(N__18861),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_6_3_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_6_3_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_6_3_6  (
            .in0(N__18840),
            .in1(N__18828),
            .in2(N__18817),
            .in3(N__18801),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_PWRGD_LC_6_3_7 .C_ON=1'b0;
    defparam \POWERLED.VCCST_PWRGD_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_PWRGD_LC_6_3_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.VCCST_PWRGD_LC_6_3_7  (
            .in0(N__18757),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30424),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_6_4_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_6_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__22945),
            .in2(N__22846),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI22EQ2_LC_6_4_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI22EQ2_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI22EQ2_LC_6_4_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNI22EQ2_LC_6_4_1  (
            .in0(N__26907),
            .in1(N__25456),
            .in2(_gnd_net_),
            .in3(N__19123),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_4_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__19120),
            .in2(_gnd_net_),
            .in3(N__19093),
            .lcout(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_4_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__19089),
            .in2(_gnd_net_),
            .in3(N__19063),
            .lcout(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI58HQ2_LC_6_4_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI58HQ2_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI58HQ2_LC_6_4_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNI58HQ2_LC_6_4_4  (
            .in0(N__26908),
            .in1(N__25735),
            .in2(_gnd_net_),
            .in3(N__19060),
            .lcout(\POWERLED.count_off_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI6AIQ2_LC_6_4_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI6AIQ2_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI6AIQ2_LC_6_4_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNI6AIQ2_LC_6_4_5  (
            .in0(N__26905),
            .in1(N__25669),
            .in2(_gnd_net_),
            .in3(N__19057),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI7CJQ2_LC_6_4_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI7CJQ2_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI7CJQ2_LC_6_4_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNI7CJQ2_LC_6_4_6  (
            .in0(N__26909),
            .in1(N__19054),
            .in2(_gnd_net_),
            .in3(N__19027),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI8EKQ2_LC_6_4_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI8EKQ2_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI8EKQ2_LC_6_4_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNI8EKQ2_LC_6_4_7  (
            .in0(N__26906),
            .in1(N__19024),
            .in2(_gnd_net_),
            .in3(N__18997),
            .lcout(\POWERLED.count_off_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNI9GLQ2_LC_6_5_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNI9GLQ2_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNI9GLQ2_LC_6_5_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNI9GLQ2_LC_6_5_0  (
            .in0(N__26910),
            .in1(N__18994),
            .in2(_gnd_net_),
            .in3(N__18979),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIAIMQ2_LC_6_5_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIAIMQ2_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIAIMQ2_LC_6_5_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNIAIMQ2_LC_6_5_1  (
            .in0(N__26913),
            .in1(_gnd_net_),
            .in2(N__19216),
            .in3(N__19192),
            .lcout(\POWERLED.count_off_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIIO3P2_LC_6_5_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIIO3P2_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIIO3P2_LC_6_5_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNIIO3P2_LC_6_5_2  (
            .in0(N__26911),
            .in1(N__19188),
            .in2(_gnd_net_),
            .in3(N__19168),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIJQ4P2_LC_6_5_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIJQ4P2_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIJQ4P2_LC_6_5_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNIJQ4P2_LC_6_5_3  (
            .in0(N__26914),
            .in1(N__19164),
            .in2(_gnd_net_),
            .in3(N__19153),
            .lcout(\POWERLED.count_off_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIKS5P2_LC_6_5_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIKS5P2_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIKS5P2_LC_6_5_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNIKS5P2_LC_6_5_4  (
            .in0(N__26912),
            .in1(N__20553),
            .in2(_gnd_net_),
            .in3(N__19150),
            .lcout(\POWERLED.count_off_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNILU6P2_LC_6_5_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNILU6P2_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNILU6P2_LC_6_5_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNILU6P2_LC_6_5_5  (
            .in0(N__26915),
            .in1(N__20538),
            .in2(_gnd_net_),
            .in3(N__19147),
            .lcout(\POWERLED.count_off_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIM08P2_LC_6_5_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIM08P2_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIM08P2_LC_6_5_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIM08P2_LC_6_5_6  (
            .in0(N__20560),
            .in1(N__26916),
            .in2(_gnd_net_),
            .in3(N__19144),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNIM08PZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_6_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_6_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_12_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19141),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34013),
            .ce(N__25592),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_LC_6_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_LC_6_6_0 .LUT_INIT=16'b1110111011001000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_LC_6_6_0  (
            .in0(N__21889),
            .in1(N__20772),
            .in2(N__21122),
            .in3(N__20964),
            .lcout(\POWERLED.un1_dutycycle_53_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_6_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_6_6_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_6_6_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \POWERLED.dutycycle_14_LC_6_6_1  (
            .in0(N__29994),
            .in1(N__23115),
            .in2(N__19270),
            .in3(N__21481),
            .lcout(\POWERLED.dutycycleZ1Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34085),
            .ce(),
            .sr(N__23697));
    defparam \POWERLED.dutycycle_RNI_13_9_LC_6_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_9_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_9_LC_6_6_2 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \POWERLED.dutycycle_RNI_13_9_LC_6_6_2  (
            .in0(N__27054),
            .in1(N__20771),
            .in2(N__21121),
            .in3(N__21775),
            .lcout(\POWERLED.dutycycle_RNI_13Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI03FP9_14_LC_6_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI03FP9_14_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI03FP9_14_LC_6_6_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI03FP9_14_LC_6_6_3  (
            .in0(N__19266),
            .in1(N__29984),
            .in2(N__23116),
            .in3(N__21480),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_6_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_6_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_6_6_4  (
            .in0(N__21890),
            .in1(_gnd_net_),
            .in2(N__19258),
            .in3(N__21433),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_9_LC_6_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_9_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_9_LC_6_6_5 .LUT_INIT=16'b1111000010110100;
    LogicCell40 \POWERLED.dutycycle_RNI_14_9_LC_6_6_5  (
            .in0(N__19255),
            .in1(N__19249),
            .in2(N__19243),
            .in3(N__19236),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_6_6_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_6_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19240),
            .in3(N__25341),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_4_LC_6_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_6_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_1_4_LC_6_6_7  (
            .in0(N__20963),
            .in1(N__21888),
            .in2(N__21804),
            .in3(N__27053),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI4J2O7_1_LC_6_7_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4J2O7_1_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4J2O7_1_LC_6_7_0 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \POWERLED.func_state_RNI4J2O7_1_LC_6_7_0  (
            .in0(N__23143),
            .in1(N__19363),
            .in2(N__26768),
            .in3(N__29780),
            .lcout(\POWERLED.dutycycle_en_7 ),
            .ltout(\POWERLED.dutycycle_en_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_6_7_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_6_7_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_6_7_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.dutycycle_11_LC_6_7_1  (
            .in0(N__29992),
            .in1(N__19333),
            .in2(N__19219),
            .in3(N__21583),
            .lcout(\POWERLED.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33998),
            .ce(),
            .sr(N__23668));
    defparam \POWERLED.dutycycle_9_LC_6_7_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_9_LC_6_7_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_9_LC_6_7_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.dutycycle_9_LC_6_7_2  (
            .in0(N__19354),
            .in1(N__29993),
            .in2(N__19348),
            .in3(N__20695),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33998),
            .ce(),
            .sr(N__23668));
    defparam \POWERLED.func_state_RNI2O4A1_0_1_LC_6_7_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_0_1_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_0_1_LC_6_7_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_0_1_LC_6_7_3  (
            .in0(N__30049),
            .in1(N__23173),
            .in2(_gnd_net_),
            .in3(N__21386),
            .lcout(\POWERLED.un1_clk_100khz_39_and_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_9_LC_6_7_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_9_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_9_LC_6_7_4 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_9_LC_6_7_4  (
            .in0(N__23172),
            .in1(N__30048),
            .in2(_gnd_net_),
            .in3(N__20773),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_30_and_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4J2O7_9_LC_6_7_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4J2O7_9_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4J2O7_9_LC_6_7_5 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \POWERLED.dutycycle_RNI4J2O7_9_LC_6_7_5  (
            .in0(N__29779),
            .in1(N__26755),
            .in2(N__19357),
            .in3(N__23142),
            .lcout(\POWERLED.dutycycle_RNI4J2O7Z0Z_9 ),
            .ltout(\POWERLED.dutycycle_RNI4J2O7Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI880A9_9_LC_6_7_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI880A9_9_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI880A9_9_LC_6_7_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI880A9_9_LC_6_7_6  (
            .in0(N__19344),
            .in1(N__29990),
            .in2(N__19336),
            .in3(N__20694),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQPBP9_11_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQPBP9_11_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQPBP9_11_LC_6_7_7 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.dutycycle_RNIQPBP9_11_LC_6_7_7  (
            .in0(N__29991),
            .in1(N__19332),
            .in2(N__19324),
            .in3(N__21582),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILOQ6A_13_LC_6_8_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILOQ6A_13_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILOQ6A_13_LC_6_8_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.dutycycle_RNILOQ6A_13_LC_6_8_0  (
            .in0(N__19485),
            .in1(N__29988),
            .in2(N__19504),
            .in3(N__21492),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_9_LC_6_8_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_9_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_9_LC_6_8_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \POWERLED.dutycycle_RNI_8_9_LC_6_8_1  (
            .in0(N__21066),
            .in1(N__21359),
            .in2(_gnd_net_),
            .in3(N__20763),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_3_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_13_LC_6_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_6_8_2 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_13_LC_6_8_2  (
            .in0(N__19313),
            .in1(N__23266),
            .in2(N__19276),
            .in3(N__21528),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_13_LC_6_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_13_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_13_LC_6_8_3 .LUT_INIT=16'b0100000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_13_LC_6_8_3  (
            .in0(N__19452),
            .in1(N__19476),
            .in2(N__19273),
            .in3(N__21361),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_6_8_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_6_8_4 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_6_8_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.dutycycle_13_LC_6_8_4  (
            .in0(N__19500),
            .in1(N__29989),
            .in2(N__19489),
            .in3(N__21493),
            .lcout(\POWERLED.dutycycleZ1Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34086),
            .ce(),
            .sr(N__23646));
    defparam \POWERLED.dutycycle_RNI_12_9_LC_6_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_9_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_9_LC_6_8_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNI_12_9_LC_6_8_5  (
            .in0(N__21067),
            .in1(N__21360),
            .in2(N__21806),
            .in3(N__20764),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_12Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_9_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_9_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_9_LC_6_8_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \POWERLED.dutycycle_RNI_15_9_LC_6_8_6  (
            .in0(N__19477),
            .in1(_gnd_net_),
            .in2(N__19462),
            .in3(N__19451),
            .lcout(\POWERLED.dutycycle_RNI_15Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_9_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_9_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_9_LC_6_8_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_11_9_LC_6_8_7  (
            .in0(N__21065),
            .in1(N__20762),
            .in2(N__27145),
            .in3(N__21358),
            .lcout(\POWERLED.dutycycle_RNI_11Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_6_9_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_6_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__22357),
            .in2(N__21301),
            .in3(N__22129),
            .lcout(\POWERLED.m18_e_0 ),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_6_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_6_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__19438),
            .in2(N__22376),
            .in3(N__19423),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_6_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_6_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__23786),
            .in2(N__19420),
            .in3(N__19405),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_6_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_6_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__19402),
            .in2(N__23796),
            .in3(N__19366),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_6_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_6_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__19744),
            .in2(N__19728),
            .in3(N__19690),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_6_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_6_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__26595),
            .in2(N__19687),
            .in3(N__19648),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_6_9_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_6_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__19645),
            .in2(N__26605),
            .in3(N__19609),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_6_9_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_6_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__21939),
            .in2(N__19606),
            .in3(N__19591),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_6_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_6_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__19588),
            .in2(N__21449),
            .in3(N__19576),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_6_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__23269),
            .in2(N__19573),
            .in3(N__19537),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_6_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__19534),
            .in2(N__21562),
            .in3(N__19522),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_6_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__25366),
            .in2(N__19519),
            .in3(N__19507),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_6_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__25422),
            .in2(N__19921),
            .in3(N__19909),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_6_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_6_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__21551),
            .in2(N__19906),
            .in3(N__19891),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_6_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_6_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__19888),
            .in2(N__25377),
            .in3(N__19861),
            .lcout(\POWERLED.mult1_un47_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_6_10_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_6_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(N__25285),
            .in2(N__25431),
            .in3(N__19840),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_6_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_6_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__25426),
            .in2(N__19804),
            .in3(N__19822),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_6_11_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_6_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19819),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_6_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_6_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__25365),
            .in2(_gnd_net_),
            .in3(N__25305),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19795),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19767),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILP0F_0_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILP0F_0_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILP0F_0_LC_6_11_5 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \POWERLED.dutycycle_RNILP0F_0_LC_6_11_5  (
            .in0(N__31132),
            .in1(N__23908),
            .in2(N__20035),
            .in3(N__20017),
            .lcout(\POWERLED.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_9_5_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_9_5_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_9_5_LC_6_11_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_RNO_9_5_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__20970),
            .in2(_gnd_net_),
            .in3(N__21953),
            .lcout(\POWERLED.g3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_3_LC_6_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_3_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_3_LC_6_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_3_LC_6_12_1  (
            .in0(N__21139),
            .in1(N__21314),
            .in2(N__19948),
            .in3(N__21809),
            .lcout(),
            .ltout(\POWERLED.g0_4_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_12_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_0_LC_6_12_2  (
            .in0(N__22378),
            .in1(N__20008),
            .in2(N__19993),
            .in3(N__22143),
            .lcout(\POWERLED.N_398_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19989),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_10_5_LC_6_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_10_5_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_10_5_LC_6_12_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNO_10_5_LC_6_12_4  (
            .in0(N__21808),
            .in1(N__22142),
            .in2(N__21316),
            .in3(N__21138),
            .lcout(),
            .ltout(\POWERLED.g3_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_8_5_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_8_5_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_8_5_LC_6_12_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.dutycycle_RNO_8_5_LC_6_12_5  (
            .in0(N__19960),
            .in1(N__22377),
            .in2(N__19954),
            .in3(N__27154),
            .lcout(),
            .ltout(\POWERLED.g3_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_7_5_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_7_5_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_7_5_LC_6_12_6 .LUT_INIT=16'b1111101110111011;
    LogicCell40 \POWERLED.dutycycle_RNO_7_5_LC_6_12_6  (
            .in0(N__27430),
            .in1(N__32944),
            .in2(N__19951),
            .in3(N__19944),
            .lcout(\POWERLED.un2_count_clk_17_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20073),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20211),
            .lcout(\POWERLED.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_6_13_1  (
            .in0(N__20166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20139),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_6_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22460),
            .lcout(\POWERLED.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_6_13_7  (
            .in0(N__20115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__20077),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__20300),
            .in2(N__20056),
            .in3(N__20047),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__20044),
            .in2(N__20305),
            .in3(N__20038),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__20374),
            .in2(N__20329),
            .in3(N__20368),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__20328),
            .in2(N__20365),
            .in3(N__20356),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_6_14_5  (
            .in0(N__22213),
            .in1(N__20304),
            .in2(N__20353),
            .in3(N__20344),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_6_14_6  (
            .in0(N__20341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20335),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(\POWERLED.mult1_un145_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20332),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_15_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20324),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_15_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_15_7  (
            .in0(N__20283),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_16_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20250),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_15_LC_7_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_7_1_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_7_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_15_LC_7_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22717),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33853),
            .ce(N__27844),
            .sr(N__28226));
    defparam \PCH_PWRGD.count_RNIS94O4_13_LC_7_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIS94O4_13_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIS94O4_13_LC_7_1_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIS94O4_13_LC_7_1_1  (
            .in0(N__20391),
            .in1(N__22763),
            .in2(_gnd_net_),
            .in3(N__27807),
            .lcout(\PCH_PWRGD.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_13_LC_7_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_7_1_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_7_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_13_LC_7_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22765),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33853),
            .ce(N__27844),
            .sr(N__28226));
    defparam \PCH_PWRGD.count_RNI0G6O4_15_LC_7_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI0G6O4_15_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI0G6O4_15_LC_7_1_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNI0G6O4_15_LC_7_1_3  (
            .in0(N__22716),
            .in1(N__20398),
            .in2(_gnd_net_),
            .in3(N__27808),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(\PCH_PWRGD.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIS94O4_0_13_LC_7_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIS94O4_0_13_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIS94O4_0_13_LC_7_1_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \PCH_PWRGD.count_RNIS94O4_0_13_LC_7_1_4  (
            .in0(N__27809),
            .in1(N__20392),
            .in2(N__20383),
            .in3(N__22764),
            .lcout(\PCH_PWRGD.count_1_i_a2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIAKA42_LC_7_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIAKA42_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIAKA42_LC_7_1_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNIAKA42_LC_7_1_5  (
            .in0(N__27702),
            .in1(N__22659),
            .in2(N__22675),
            .in3(N__28225),
            .lcout(\PCH_PWRGD.count_rst_10 ),
            .ltout(\PCH_PWRGD.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISVPK4_4_LC_7_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISVPK4_4_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISVPK4_4_LC_7_1_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNISVPK4_4_LC_7_1_6  (
            .in0(N__27810),
            .in1(_gnd_net_),
            .in2(N__20380),
            .in3(N__24159),
            .lcout(\PCH_PWRGD.un2_count_1_axb_4 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_7_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_7_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_7_1_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_4_LC_7_1_7  (
            .in0(N__27703),
            .in1(N__28227),
            .in2(N__20377),
            .in3(N__22660),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33853),
            .ce(N__27844),
            .sr(N__28226));
    defparam \PCH_PWRGD.count_14_LC_7_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_7_2_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_7_2_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \PCH_PWRGD.count_14_LC_7_2_0  (
            .in0(N__22741),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28224),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33996),
            .ce(N__27834),
            .sr(N__28243));
    defparam \PCH_PWRGD.count_RNIOPNK4_2_LC_7_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOPNK4_2_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOPNK4_2_LC_7_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIOPNK4_2_LC_7_2_1  (
            .in0(N__20454),
            .in1(N__27833),
            .in2(_gnd_net_),
            .in3(N__22523),
            .lcout(\PCH_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_2_LC_7_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_7_2_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_7_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_2_LC_7_2_2  (
            .in0(N__22525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33996),
            .ce(N__27834),
            .sr(N__28243));
    defparam \PCH_PWRGD.count_RNIUC5O4_14_LC_7_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIUC5O4_14_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIUC5O4_14_LC_7_2_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \PCH_PWRGD.count_RNIUC5O4_14_LC_7_2_3  (
            .in0(N__28223),
            .in1(N__22740),
            .in2(N__20464),
            .in3(N__27832),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(\PCH_PWRGD.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOPNK4_0_2_LC_7_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOPNK4_0_2_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOPNK4_0_2_LC_7_2_4 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \PCH_PWRGD.count_RNIOPNK4_0_2_LC_7_2_4  (
            .in0(N__22524),
            .in1(N__20455),
            .in2(N__20446),
            .in3(N__27811),
            .lcout(\PCH_PWRGD.count_1_i_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_12_LC_7_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_7_2_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_7_2_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_12_LC_7_2_6  (
            .in0(N__22783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33996),
            .ce(N__27834),
            .sr(N__28243));
    defparam \PCH_PWRGD.count_RNIQ63O4_12_LC_7_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQ63O4_12_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQ63O4_12_LC_7_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIQ63O4_12_LC_7_2_7  (
            .in0(N__20443),
            .in1(N__22782),
            .in2(_gnd_net_),
            .in3(N__27831),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_0_LC_7_3_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_0_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_0_LC_7_3_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_0_LC_7_3_1  (
            .in0(_gnd_net_),
            .in1(N__22692),
            .in2(_gnd_net_),
            .in3(N__22707),
            .lcout(\RSMRST_PWRGD.m4_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIKA9Q3_LC_7_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIKA9Q3_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIKA9Q3_LC_7_3_3 .LUT_INIT=16'b1110111100100000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIKA9Q3_LC_7_3_3  (
            .in0(N__24710),
            .in1(N__20416),
            .in2(N__30811),
            .in3(N__20406),
            .lcout(PCH_PWRGD_delayed_vccin_ok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_7_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_7_3_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_7_3_4  (
            .in0(_gnd_net_),
            .in1(N__28278),
            .in2(N__31267),
            .in3(N__28300),
            .lcout(\PCH_PWRGD.N_250_0 ),
            .ltout(\PCH_PWRGD.N_250_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_7_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_7_3_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_7_3_5 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_7_3_5  (
            .in0(N__30807),
            .in1(N__20407),
            .in2(N__20410),
            .in3(N__24711),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33875),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_0_LC_7_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_0_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI2UUH1_0_LC_7_3_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI2UUH1_0_LC_7_3_7  (
            .in0(N__28299),
            .in1(N__31263),
            .in2(_gnd_net_),
            .in3(N__28384),
            .lcout(\PCH_PWRGD.curr_state_RNI2UUH1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI39MT5_0_LC_7_4_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI39MT5_0_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI39MT5_0_LC_7_4_0 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \POWERLED.dutycycle_RNI39MT5_0_LC_7_4_0  (
            .in0(N__20472),
            .in1(N__29807),
            .in2(N__20515),
            .in3(N__20524),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(\POWERLED.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNII3LM3_0_LC_7_4_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNII3LM3_0_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNII3LM3_0_LC_7_4_1 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \POWERLED.dutycycle_RNII3LM3_0_LC_7_4_1  (
            .in0(N__26715),
            .in1(N__31158),
            .in2(N__20527),
            .in3(N__21327),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(\POWERLED.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_7_4_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_7_4_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_7_4_2 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_0_LC_7_4_2  (
            .in0(N__20473),
            .in1(N__20514),
            .in2(N__20518),
            .in3(N__29809),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33997),
            .ce(),
            .sr(N__23669));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_4_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_4_3 .LUT_INIT=16'b1100111101011111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_4_3  (
            .in0(N__20626),
            .in1(N__26164),
            .in2(N__25027),
            .in3(N__29332),
            .lcout(\POWERLED.dutycycle_1_0_1 ),
            .ltout(\POWERLED.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_7_4_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_7_4_4 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_7_4_4 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \POWERLED.dutycycle_1_LC_7_4_4  (
            .in0(N__20497),
            .in1(N__20485),
            .in2(N__20500),
            .in3(N__29810),
            .lcout(\POWERLED.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33997),
            .ce(),
            .sr(N__23669));
    defparam \POWERLED.dutycycle_RNII3LM3_1_LC_7_4_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNII3LM3_1_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNII3LM3_1_LC_7_4_5 .LUT_INIT=16'b1010101011111011;
    LogicCell40 \POWERLED.dutycycle_RNII3LM3_1_LC_7_4_5  (
            .in0(N__26716),
            .in1(N__31159),
            .in2(N__22106),
            .in3(N__21328),
            .lcout(\POWERLED.dutycycle_eena_0 ),
            .ltout(\POWERLED.dutycycle_eena_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI7KKU5_1_LC_7_4_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI7KKU5_1_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI7KKU5_1_LC_7_4_6 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_RNI7KKU5_1_LC_7_4_6  (
            .in0(N__20491),
            .in1(N__20484),
            .in2(N__20476),
            .in3(N__29808),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_7_4_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_0_LC_7_4_7 .LUT_INIT=16'b1100111110101111;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_0_LC_7_4_7  (
            .in0(N__22322),
            .in1(N__26163),
            .in2(N__25026),
            .in3(N__29331),
            .lcout(\POWERLED.dutycycle_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNISKPU6_0_LC_7_5_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNISKPU6_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNISKPU6_0_LC_7_5_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \POWERLED.func_state_RNISKPU6_0_LC_7_5_0  (
            .in0(N__24282),
            .in1(N__29985),
            .in2(N__26092),
            .in3(N__29772),
            .lcout(\POWERLED.func_state_RNISKPU6Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNISKPU6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIVAIU9_13_LC_7_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIVAIU9_13_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIVAIU9_13_LC_7_5_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \POWERLED.count_off_RNIVAIU9_13_LC_7_5_1  (
            .in0(N__20608),
            .in1(_gnd_net_),
            .in2(N__20611),
            .in3(N__20599),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_7_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_7_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_13_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20607),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34293),
            .ce(N__25557),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_7_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_7_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_15_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20577),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34293),
            .ce(N__25557),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_7_5_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_7_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_14_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20593),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34293),
            .ce(N__25557),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI1EJU9_14_LC_7_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI1EJU9_14_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI1EJU9_14_LC_7_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNI1EJU9_14_LC_7_5_5  (
            .in0(N__20592),
            .in1(N__20584),
            .in2(_gnd_net_),
            .in3(N__25517),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI3HKU9_15_LC_7_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI3HKU9_15_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI3HKU9_15_LC_7_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.count_off_RNI3HKU9_15_LC_7_5_6  (
            .in0(N__25558),
            .in1(N__20578),
            .in2(_gnd_net_),
            .in3(N__20566),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(\POWERLED.count_offZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_7_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_7_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_7_5_7  (
            .in0(N__20554),
            .in1(N__22839),
            .in2(N__20542),
            .in3(N__20539),
            .lcout(\POWERLED.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_3_LC_7_6_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_3_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_3_LC_7_6_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_3_LC_7_6_0  (
            .in0(N__21299),
            .in1(N__21807),
            .in2(N__20647),
            .in3(N__27423),
            .lcout(\POWERLED.dutycycle_RNI_10Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_7_6_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_7_6_1 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_7_6_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.dutycycle_6_LC_7_6_1  (
            .in0(N__23982),
            .in1(N__20665),
            .in2(N__29806),
            .in3(N__22882),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34084),
            .ce(),
            .sr(N__23695));
    defparam \POWERLED.dutycycle_RNIEP8SA_6_LC_7_6_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEP8SA_6_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEP8SA_6_LC_7_6_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_RNIEP8SA_6_LC_7_6_2  (
            .in0(N__20664),
            .in1(N__29759),
            .in2(N__23983),
            .in3(N__22881),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(\POWERLED.dutycycleZ1Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_0_LC_7_6_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_7_6_3 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_0_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__22094),
            .in2(N__20653),
            .in3(N__22343),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNI_5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_LC_7_6_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_LC_7_6_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20650),
            .in3(N__26579),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_0_LC_7_6_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_7_6_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_0_LC_7_6_5  (
            .in0(N__32969),
            .in1(N__22093),
            .in2(_gnd_net_),
            .in3(N__22342),
            .lcout(\POWERLED.un1_dutycycle_96_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_1_LC_7_6_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_1_LC_7_6_6 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \POWERLED.func_state_RNI_6_1_LC_7_6_6  (
            .in0(N__32971),
            .in1(N__27424),
            .in2(N__20638),
            .in3(N__23881),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_3_LC_7_6_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_3_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_3_LC_7_6_7 .LUT_INIT=16'b1100111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_13_3_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__26239),
            .in2(N__20629),
            .in3(N__26476),
            .lcout(\POWERLED.un1_dutycycle_172_m3s4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_7_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_7_7_0 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \POWERLED.dutycycle_RNI_3_0_LC_7_7_0  (
            .in0(N__22086),
            .in1(_gnd_net_),
            .in2(N__22356),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__23005),
            .in2(N__22112),
            .in3(N__20617),
            .lcout(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__23009),
            .in2(N__23790),
            .in3(N__20614),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI765B1_LC_7_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI765B1_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI765B1_LC_7_7_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI765B1_LC_7_7_3  (
            .in0(N__29944),
            .in1(N__23006),
            .in2(N__21315),
            .in3(N__21169),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI765BZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI886B1_LC_7_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI886B1_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI886B1_LC_7_7_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI886B1_LC_7_7_4  (
            .in0(N__29983),
            .in1(N__23010),
            .in2(N__21813),
            .in3(N__21148),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI886BZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__23007),
            .in2(N__26600),
            .in3(N__21145),
            .lcout(\POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_7_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__23011),
            .in2(N__27078),
            .in3(N__21142),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4A1_LC_7_7_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4A1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4A1_LC_7_7_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4A1_LC_7_7_7  (
            .in0(N__29943),
            .in1(N__23008),
            .in2(N__21123),
            .in3(N__20974),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI2O4AZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNICGAB1_LC_7_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNICGAB1_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNICGAB1_LC_7_8_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNICGAB1_LC_7_8_0  (
            .in0(N__29916),
            .in1(N__23002),
            .in2(N__20962),
            .in3(N__20818),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNICGABZ0Z1 ),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_7_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_7_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__23012),
            .in2(N__20774),
            .in3(N__20686),
            .lcout(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCB1_LC_7_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCB1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCB1_LC_7_8_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCB1_LC_7_8_2  (
            .in0(N__29917),
            .in1(N__23003),
            .in2(N__21954),
            .in3(N__20668),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNIEKCBZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__23013),
            .in2(N__21438),
            .in3(N__21574),
            .lcout(\POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__23004),
            .in2(N__23229),
            .in3(N__21571),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__23014),
            .in2(N__21547),
            .in3(N__21484),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_8_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__23001),
            .in2(N__25370),
            .in3(N__21469),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_8_7 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_7_8_7  (
            .in0(N__25427),
            .in1(_gnd_net_),
            .in2(N__27411),
            .in3(N__21466),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_7_9_0 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_7_9_0  (
            .in0(N__24233),
            .in1(N__21621),
            .in2(N__26156),
            .in3(N__24246),
            .lcout(\POWERLED.N_396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_7_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_7_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21439),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_2_2_LC_7_9_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_2_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_2_LC_7_9_2 .LUT_INIT=16'b0101110111011101;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_2_2_LC_7_9_2  (
            .in0(N__25019),
            .in1(N__32956),
            .in2(N__24235),
            .in3(N__21620),
            .lcout(\POWERLED.dutycycle_RNI2O4A1_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIA02P1_1_LC_7_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIA02P1_1_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIA02P1_1_LC_7_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \POWERLED.func_state_RNIA02P1_1_LC_7_9_3  (
            .in0(N__23346),
            .in1(N__26212),
            .in2(_gnd_net_),
            .in3(N__21651),
            .lcout(\POWERLED.N_115_f0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_6_LC_7_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_7_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_6_LC_7_9_4  (
            .in0(N__26594),
            .in1(N__29426),
            .in2(N__24082),
            .in3(N__27069),
            .lcout(\POWERLED.N_366 ),
            .ltout(\POWERLED.N_366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_6_LC_7_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_6_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_6_LC_7_9_5 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_6_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__29914),
            .in2(N__21640),
            .in3(N__24234),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI2O4A1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI4G9K2_1_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4G9K2_1_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4G9K2_1_LC_7_9_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \POWERLED.func_state_RNI4G9K2_1_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__27412),
            .in2(N__21637),
            .in3(N__21634),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI68EU3_1_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI68EU3_1_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI68EU3_1_LC_7_9_7 .LUT_INIT=16'b1111000001110111;
    LogicCell40 \POWERLED.func_state_RNI68EU3_1_LC_7_9_7  (
            .in0(N__29425),
            .in1(N__29913),
            .in2(N__21628),
            .in3(N__26470),
            .lcout(\POWERLED.func_state_RNI68EU3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_0_o2_0_6_LC_7_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_0_o2_0_6_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_0_o2_0_6_LC_7_10_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_0_o2_0_6_LC_7_10_0  (
            .in0(N__29061),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21965),
            .lcout(\POWERLED.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_7_10_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_7_10_1  (
            .in0(N__24228),
            .in1(N__21625),
            .in2(_gnd_net_),
            .in3(N__26151),
            .lcout(\POWERLED.func_state_RNI_0Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_0_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_0_LC_7_10_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \POWERLED.func_state_RNIOGRS_0_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__28962),
            .in2(N__21604),
            .in3(N__31116),
            .lcout(\POWERLED.func_state_RNIOGRSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_fast_LC_7_10_3 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_fast_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_fast_LC_7_10_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \COUNTER.tmp_0_fast_LC_7_10_3  (
            .in0(N__21967),
            .in1(_gnd_net_),
            .in2(N__25123),
            .in3(_gnd_net_),
            .lcout(SUSWARN_N_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34240),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIT69J5_1_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIT69J5_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIT69J5_1_LC_7_10_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \POWERLED.func_state_RNIT69J5_1_LC_7_10_4  (
            .in0(N__25860),
            .in1(N__31115),
            .in2(_gnd_net_),
            .in3(N__21601),
            .lcout(\POWERLED.func_state_RNIT69J5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI98TE_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI98TE_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI98TE_LC_7_10_5 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI98TE_LC_7_10_5  (
            .in0(N__21595),
            .in1(N__29474),
            .in2(N__27348),
            .in3(N__29318),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI919H1_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI919H1_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI919H1_LC_7_10_6 .LUT_INIT=16'b1000111111001111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI919H1_LC_7_10_6  (
            .in0(N__29062),
            .in1(N__27335),
            .in2(N__21970),
            .in3(N__21966),
            .lcout(\POWERLED.un1_dutycycle_94_cry_4_c_RNI919HZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_4_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_7_10_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_4_LC_7_10_7  (
            .in0(N__21950),
            .in1(N__21820),
            .in2(N__21814),
            .in3(N__27140),
            .lcout(\POWERLED.m18_e_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_eena_14_0_0_LC_7_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_eena_14_0_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_eena_14_0_0_LC_7_11_0 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \POWERLED.dutycycle_eena_14_0_0_LC_7_11_0  (
            .in0(N__28901),
            .in1(N__26404),
            .in2(N__27339),
            .in3(N__29712),
            .lcout(\POWERLED.dutycycle_eena_14_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_7_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_2_LC_7_11_2 .LUT_INIT=16'b0011010100111111;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_2_LC_7_11_2  (
            .in0(N__29459),
            .in1(N__23757),
            .in2(N__26249),
            .in3(N__29995),
            .lcout(\POWERLED.un1_dutycycle_172_m1_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_rep1_LC_7_11_3 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_rep1_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_rep1_LC_7_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_0_rep1_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__23534),
            .in2(_gnd_net_),
            .in3(N__25117),
            .lcout(SUSWARN_N_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34162),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_m2_0_a2_iso_LC_7_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_m2_0_a2_iso_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_m2_0_a2_iso_LC_7_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_m2_0_a2_iso_LC_7_11_4  (
            .in0(N__27315),
            .in1(N__23473),
            .in2(N__26411),
            .in3(N__30574),
            .lcout(\POWERLED.func_m2_0_a2_isoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIVR902_LC_7_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIVR902_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIVR902_LC_7_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIVR902_LC_7_11_5  (
            .in0(N__34565),
            .in1(N__21661),
            .in2(_gnd_net_),
            .in3(N__30190),
            .lcout(\POWERLED.dutycycle_1_0_5 ),
            .ltout(\POWERLED.dutycycle_1_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIBFCJ3_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIBFCJ3_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIBFCJ3_LC_7_11_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIBFCJ3_LC_7_11_6  (
            .in0(N__23535),
            .in1(N__25118),
            .in2(N__21655),
            .in3(N__26210),
            .lcout(\POWERLED.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJ2BQ2_2_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJ2BQ2_2_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJ2BQ2_2_LC_7_11_7 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \POWERLED.dutycycle_RNIJ2BQ2_2_LC_7_11_7  (
            .in0(N__26682),
            .in1(N__26209),
            .in2(N__21994),
            .in3(N__21652),
            .lcout(\POWERLED.dutycycle_eena_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_155_LC_7_12_0 .C_ON=1'b0;
    defparam \POWERLED.G_155_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_155_LC_7_12_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.G_155_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23536),
            .in3(N__25110),
            .lcout(G_155),
            .ltout(G_155_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJDU46_2_LC_7_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJDU46_2_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJDU46_2_LC_7_12_1 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_RNIJDU46_2_LC_7_12_1  (
            .in0(N__22021),
            .in1(N__22002),
            .in2(N__22024),
            .in3(N__22014),
            .lcout(\POWERLED.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIFRMD2_LC_7_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIFRMD2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIFRMD2_LC_7_12_2 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIFRMD2_LC_7_12_2  (
            .in0(N__21976),
            .in1(N__29469),
            .in2(N__26947),
            .in3(N__29316),
            .lcout(\POWERLED.N_73 ),
            .ltout(\POWERLED.N_73_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_7_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_7_12_3 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_7_12_3 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \POWERLED.dutycycle_2_LC_7_12_3  (
            .in0(N__29711),
            .in1(N__22015),
            .in2(N__22006),
            .in3(N__22003),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34224),
            .ce(),
            .sr(N__23615));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_12_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_12_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_12_4  (
            .in0(N__23760),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILP0F_2_LC_7_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILP0F_2_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILP0F_2_LC_7_12_5 .LUT_INIT=16'b0100010011001000;
    LogicCell40 \POWERLED.dutycycle_RNILP0F_2_LC_7_12_5  (
            .in0(N__29317),
            .in1(N__31120),
            .in2(N__29481),
            .in3(N__23759),
            .lcout(\POWERLED.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_12_6 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIF01V_LC_7_12_6  (
            .in0(N__30238),
            .in1(N__21985),
            .in2(N__31154),
            .in3(N__29315),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOBHB2_0_LC_7_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOBHB2_0_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOBHB2_0_LC_7_12_7 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \POWERLED.func_state_RNIOBHB2_0_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__29458),
            .in2(N__26001),
            .in3(N__26942),
            .lcout(\POWERLED.func_state_1_m2_am_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_7_13_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_7_13_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_7_13_0  (
            .in0(N__23875),
            .in1(N__23761),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_331 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__22267),
            .in2(N__22179),
            .in3(N__22261),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__22175),
            .in2(N__22258),
            .in3(N__22249),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__22246),
            .in2(N__22223),
            .in3(N__22240),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__22237),
            .in2(N__22224),
            .in3(N__22192),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_13_5  (
            .in0(N__22459),
            .in1(N__22189),
            .in2(N__22180),
            .in3(N__22162),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_13_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__22159),
            .in2(_gnd_net_),
            .in3(N__22153),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(\POWERLED.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_7_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_7_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22150),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_7_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_7_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__22144),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__22433),
            .in2(N__22510),
            .in3(N__22495),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__22492),
            .in2(N__22438),
            .in3(N__22486),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__22461),
            .in2(N__22483),
            .in3(N__22474),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__22471),
            .in2(N__22465),
            .in3(N__22441),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_14_5  (
            .in0(N__22600),
            .in1(N__22437),
            .in2(N__22423),
            .in3(N__22414),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_14_6  (
            .in0(N__22411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22405),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(\POWERLED.mult1_un159_sum_s_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_14_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22402),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_7_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__22366),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_7_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_7_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(N__22580),
            .in2(N__22282),
            .in3(N__22601),
            .lcout(G_2078),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_7_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_7_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__22627),
            .in2(N__22585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_7_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_7_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__22602),
            .in2(N__22621),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_7_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_7_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__22612),
            .in2(N__22606),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_7_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_7_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(N__22584),
            .in2(N__22570),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_7_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_7_15_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_7_15_6  (
            .in0(N__22561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22555),
            .lcout(\POWERLED.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_9_LC_7_16_6 .C_ON=1'b0;
    defparam \POWERLED.G_9_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_9_LC_7_16_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.G_9_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__30612),
            .in2(_gnd_net_),
            .in3(N__25122),
            .lcout(G_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_8_1_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_LC_8_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__27605),
            .in2(N__27628),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI8G842_LC_8_1_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI8G842_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI8G842_LC_8_1_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNI8G842_LC_8_1_1  (
            .in0(N__28218),
            .in1(N__22531),
            .in2(_gnd_net_),
            .in3(N__22513),
            .lcout(\PCH_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_8_1_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_8_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__24140),
            .in2(_gnd_net_),
            .in3(N__22678),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_8_1_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_8_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__22671),
            .in2(_gnd_net_),
            .in3(N__22651),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_8_1_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_8_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__27973),
            .in2(_gnd_net_),
            .in3(N__22648),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_8_1_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_8_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__24484),
            .in2(_gnd_net_),
            .in3(N__22645),
            .lcout(\PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_8_1_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_8_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28009),
            .in3(N__22642),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_8_1_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_8_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_8_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27464),
            .in3(N__22639),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_8_2_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_8_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__27525),
            .in2(_gnd_net_),
            .in3(N__22636),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIG0H42_LC_8_2_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIG0H42_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIG0H42_LC_8_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNIG0H42_LC_8_2_1  (
            .in0(N__28204),
            .in1(N__24352),
            .in2(_gnd_net_),
            .in3(N__22633),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_8_2_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_8_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27898),
            .in3(N__22630),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIP94V1_LC_8_2_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIP94V1_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIP94V1_LC_8_2_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNIP94V1_LC_8_2_3  (
            .in0(N__28205),
            .in1(N__24438),
            .in2(_gnd_net_),
            .in3(N__22774),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIQB5V1_LC_8_2_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIQB5V1_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIQB5V1_LC_8_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNIQB5V1_LC_8_2_4  (
            .in0(N__28222),
            .in1(N__22771),
            .in2(_gnd_net_),
            .in3(N__22750),
            .lcout(\PCH_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_8_2_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_8_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__22747),
            .in2(_gnd_net_),
            .in3(N__22729),
            .lcout(\PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNISF7V1_LC_8_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNISF7V1_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNISF7V1_LC_8_2_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNISF7V1_LC_8_2_6  (
            .in0(N__22726),
            .in1(N__28206),
            .in2(_gnd_net_),
            .in3(N__22720),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIHNMD2_1_LC_8_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIHNMD2_1_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIHNMD2_1_LC_8_2_7 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIHNMD2_1_LC_8_2_7  (
            .in0(N__28203),
            .in1(N__28357),
            .in2(_gnd_net_),
            .in3(N__29827),
            .lcout(\PCH_PWRGD.curr_state_RNIHNMD2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_8_3_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_8_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_8_3_0  (
            .in0(N__34858),
            .in1(N__24742),
            .in2(N__24805),
            .in3(N__24804),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_1_LC_8_3_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_8_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_8_3_1  (
            .in0(N__34851),
            .in1(N__22708),
            .in2(_gnd_net_),
            .in3(N__22696),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_2_LC_8_3_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_8_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_8_3_2  (
            .in0(N__34859),
            .in1(N__22693),
            .in2(_gnd_net_),
            .in3(N__22681),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_3_LC_8_3_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_8_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_8_3_3  (
            .in0(N__34852),
            .in1(N__24520),
            .in2(_gnd_net_),
            .in3(N__22810),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_4_LC_8_3_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_8_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_8_3_4  (
            .in0(N__34860),
            .in1(N__24631),
            .in2(_gnd_net_),
            .in3(N__22807),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_5_LC_8_3_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_8_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_8_3_5  (
            .in0(N__34853),
            .in1(N__24559),
            .in2(_gnd_net_),
            .in3(N__22804),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_6_LC_8_3_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_8_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_8_3_6  (
            .in0(N__34861),
            .in1(N__24547),
            .in2(_gnd_net_),
            .in3(N__22801),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_7_LC_8_3_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_8_3_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_8_3_7  (
            .in0(N__34854),
            .in1(N__24534),
            .in2(_gnd_net_),
            .in3(N__22798),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__34144),
            .ce(),
            .sr(N__25165));
    defparam \RSMRST_PWRGD.count_8_LC_8_4_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_8_4_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_8_4_0  (
            .in0(N__34850),
            .in1(N__24643),
            .in2(_gnd_net_),
            .in3(N__22795),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.count_9_LC_8_4_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_8_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_8_4_1  (
            .in0(N__34846),
            .in1(N__24655),
            .in2(_gnd_net_),
            .in3(N__22792),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.count_10_LC_8_4_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_8_4_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_8_4_2  (
            .in0(N__34847),
            .in1(N__24781),
            .in2(_gnd_net_),
            .in3(N__22789),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.count_11_LC_8_4_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_8_4_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_8_4_3  (
            .in0(N__34844),
            .in1(N__24616),
            .in2(_gnd_net_),
            .in3(N__22786),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.count_12_LC_8_4_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_8_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_8_4_4  (
            .in0(N__34848),
            .in1(N__24577),
            .in2(_gnd_net_),
            .in3(N__22867),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.count_13_LC_8_4_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_8_4_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_8_4_5  (
            .in0(N__34845),
            .in1(N__24769),
            .in2(_gnd_net_),
            .in3(N__22864),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.count_14_LC_8_4_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_8_4_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_8_4_6  (
            .in0(N__34849),
            .in1(N__24604),
            .in2(_gnd_net_),
            .in3(N__22861),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__34080),
            .ce(),
            .sr(N__25173));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(N__34557),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_8_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__24591),
            .in2(_gnd_net_),
            .in3(N__22858),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34324),
            .ce(N__25135),
            .sr(N__25180));
    defparam \POWERLED.count_off_RNIBQDB2_0_LC_8_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIBQDB2_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIBQDB2_0_LC_8_6_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_off_RNIBQDB2_0_LC_8_6_0  (
            .in0(N__26862),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22837),
            .lcout(),
            .ltout(\POWERLED.count_off_RNIBQDB2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI2KLI9_0_LC_8_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI2KLI9_0_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI2KLI9_0_LC_8_6_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNI2KLI9_0_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__22816),
            .in2(N__22855),
            .in3(N__25496),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(\POWERLED.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_8_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_8_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22852),
            .in3(N__22941),
            .lcout(\POWERLED.count_off_RNIZ0Z_1 ),
            .ltout(\POWERLED.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_8_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_8_6_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.count_off_1_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22849),
            .in3(N__26864),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34233),
            .ce(N__25583),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_8_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_8_6_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_off_0_LC_8_6_4  (
            .in0(N__26863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22838),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34233),
            .ce(N__25583),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI3LLI9_1_LC_8_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI3LLI9_1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI3LLI9_1_LC_8_6_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.count_off_RNI3LLI9_1_LC_8_6_5  (
            .in0(N__22960),
            .in1(N__25495),
            .in2(N__22954),
            .in3(N__26861),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(\POWERLED.count_offZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_1_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_1_LC_8_6_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_1_LC_8_6_6  (
            .in0(N__25734),
            .in1(N__25668),
            .in2(N__22927),
            .in3(N__25455),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_10_LC_8_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_10_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_10_LC_8_6_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_10_LC_8_6_7  (
            .in0(N__22924),
            .in1(N__22918),
            .in2(N__22906),
            .in3(N__22903),
            .lcout(\POWERLED.count_off_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIRGL41_LC_8_7_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIRGL41_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIRGL41_LC_8_7_0 .LUT_INIT=16'b1010100011111101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIRGL41_LC_8_7_0  (
            .in0(N__31026),
            .in1(N__29382),
            .in2(N__23089),
            .in3(N__22891),
            .lcout(),
            .ltout(\POWERLED.N_220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI4L823_LC_8_7_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI4L823_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI4L823_LC_8_7_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI4L823_LC_8_7_1  (
            .in0(N__30149),
            .in1(N__26693),
            .in2(N__22885),
            .in3(N__29305),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNI4LZ0Z823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_0_0_LC_8_7_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_0_0_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_0_0_LC_8_7_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \POWERLED.func_state_RNIOGRS_0_0_LC_8_7_2  (
            .in0(N__31027),
            .in1(N__29383),
            .in2(N__29573),
            .in3(N__28984),
            .lcout(),
            .ltout(\POWERLED.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHGMD3_1_LC_8_7_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHGMD3_1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHGMD3_1_LC_8_7_3 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \POWERLED.func_state_RNIHGMD3_1_LC_8_7_3  (
            .in0(N__23026),
            .in1(N__26694),
            .in2(N__22870),
            .in3(N__29306),
            .lcout(\POWERLED.func_state_1_ss0_i_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_0_LC_8_7_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_0_LC_8_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_2_0_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26155),
            .lcout(\POWERLED.N_2216_i ),
            .ltout(\POWERLED.N_2216_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJ9IE1_1_LC_8_7_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJ9IE1_1_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJ9IE1_1_LC_8_7_5 .LUT_INIT=16'b1101110111001101;
    LogicCell40 \POWERLED.func_state_RNIJ9IE1_1_LC_8_7_5  (
            .in0(N__29333),
            .in1(N__26692),
            .in2(N__23095),
            .in3(N__23848),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m2s2_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIN2PE3_1_LC_8_7_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIN2PE3_1_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIN2PE3_1_LC_8_7_6 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \POWERLED.func_state_RNIN2PE3_1_LC_8_7_6  (
            .in0(N__29307),
            .in1(N__25186),
            .in2(N__23092),
            .in3(N__23025),
            .lcout(\POWERLED.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIMJCH1_10_LC_8_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIMJCH1_10_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIMJCH1_10_LC_8_7_7 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \POWERLED.count_off_RNIMJCH1_10_LC_8_7_7  (
            .in0(N__28983),
            .in1(N__23088),
            .in2(N__29574),
            .in3(N__31028),
            .lcout(\POWERLED.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_1_0_LC_8_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_1_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_1_0_LC_8_8_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_1_0_LC_8_8_0  (
            .in0(N__29915),
            .in1(N__32952),
            .in2(_gnd_net_),
            .in3(N__30037),
            .lcout(\POWERLED.N_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.slp_s3n_signal_2_LC_8_8_1 .C_ON=1'b0;
    defparam \POWERLED.slp_s3n_signal_2_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.slp_s3n_signal_2_LC_8_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.slp_s3n_signal_2_LC_8_8_1  (
            .in0(N__27346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26969),
            .lcout(slp_s3n_signal),
            .ltout(slp_s3n_signal_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_8_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_8_2 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_8_8_2  (
            .in0(N__28982),
            .in1(_gnd_net_),
            .in2(N__23029),
            .in3(N__30465),
            .lcout(\POWERLED.N_183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_m1_0_a2_LC_8_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_m1_0_a2_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_m1_0_a2_LC_8_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.un1_m1_0_a2_LC_8_8_3  (
            .in0(N__27347),
            .in1(N__29040),
            .in2(_gnd_net_),
            .in3(N__26070),
            .lcout(\POWERLED.un1_N_3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_8_8_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_8_8_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29392),
            .in3(N__29301),
            .lcout(\POWERLED.func_state_RNIZ0Z_1 ),
            .ltout(\POWERLED.func_state_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_8_1_LC_8_8_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_8_1_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_8_1_LC_8_8_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_8_1_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23017),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_162_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIET094_1_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIET094_1_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIET094_1_LC_8_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_RNIET094_1_LC_8_8_6  (
            .in0(N__25817),
            .in1(N__26211),
            .in2(N__23457),
            .in3(N__23345),
            .lcout(\POWERLED.N_399_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIV0AS_1_LC_8_8_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIV0AS_1_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIV0AS_1_LC_8_8_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.func_state_RNIV0AS_1_LC_8_8_7  (
            .in0(N__27345),
            .in1(N__26069),
            .in2(N__29330),
            .in3(N__29371),
            .lcout(\POWERLED.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4J2O7_12_LC_8_9_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4J2O7_12_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4J2O7_12_LC_8_9_0 .LUT_INIT=16'b1000100010001010;
    LogicCell40 \POWERLED.dutycycle_RNI4J2O7_12_LC_8_9_0  (
            .in0(N__29744),
            .in1(N__26678),
            .in2(N__23136),
            .in3(N__23179),
            .lcout(\POWERLED.dutycycle_en_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_8_9_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.dutycycle_12_LC_8_9_1  (
            .in0(N__23287),
            .in1(N__23311),
            .in2(N__23302),
            .in3(N__29939),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34449),
            .ce(),
            .sr(N__23664));
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_1_LC_8_9_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_1_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__24991),
            .in2(_gnd_net_),
            .in3(N__29202),
            .lcout(\POWERLED.func_state_RNI2O4A1Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI2O4A1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_1_1_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_1_1_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_1_1_LC_8_9_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_1_1_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23314),
            .in3(_gnd_net_),
            .lcout(\POWERLED.func_state_RNI2O4A1_1Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI2O4A1_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNISSCP9_12_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNISSCP9_12_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNISSCP9_12_LC_8_9_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.dutycycle_RNISSCP9_12_LC_8_9_4  (
            .in0(N__23310),
            .in1(N__23298),
            .in2(N__23290),
            .in3(N__23286),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(\POWERLED.dutycycleZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_12_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_12_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_12_LC_8_9_5 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_12_LC_8_9_5  (
            .in0(N__30038),
            .in1(_gnd_net_),
            .in2(N__23182),
            .in3(N__23162),
            .lcout(\POWERLED.un1_clk_100khz_42_and_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_14_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_14_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_14_LC_8_9_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_14_LC_8_9_6  (
            .in0(N__30050),
            .in1(N__25375),
            .in2(_gnd_net_),
            .in3(N__23166),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_47_and_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4J2O7_14_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4J2O7_14_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4J2O7_14_LC_8_9_7 .LUT_INIT=16'b1000100010001100;
    LogicCell40 \POWERLED.dutycycle_RNI4J2O7_14_LC_8_9_7  (
            .in0(N__26677),
            .in1(N__29743),
            .in2(N__23146),
            .in3(N__23129),
            .lcout(\POWERLED.dutycycle_en_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_3_LC_8_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_3_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_3_LC_8_10_0 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \POWERLED.dutycycle_RNI_11_3_LC_8_10_0  (
            .in0(N__27420),
            .in1(N__23494),
            .in2(N__32970),
            .in3(N__23479),
            .lcout(\POWERLED.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_8_10_1 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.func_state_0_LC_8_10_1  (
            .in0(N__23392),
            .in1(N__30165),
            .in2(N__25903),
            .in3(N__23398),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34425),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_m2_0_a2_0_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_m2_0_a2_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_m2_0_a2_0_LC_8_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.func_m2_0_a2_0_LC_8_10_2  (
            .in0(N__29060),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28979),
            .lcout(\POWERLED.func_m2_0_a2Z0Z_0 ),
            .ltout(\POWERLED.func_m2_0_a2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_m2_0_a2_LC_8_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_m2_0_a2_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_m2_0_a2_LC_8_10_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_m2_0_a2_LC_8_10_3  (
            .in0(N__26386),
            .in1(N__27319),
            .in2(N__23467),
            .in3(N__23532),
            .lcout(\POWERLED.func_N_5_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2O4A1_0_10_LC_8_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2O4A1_0_10_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2O4A1_0_10_LC_8_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_RNI2O4A1_0_10_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__29896),
            .in2(_gnd_net_),
            .in3(N__32951),
            .lcout(\POWERLED.count_clk_RNI2O4A1_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI91IA4_0_1_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI91IA4_0_1_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI91IA4_0_1_LC_8_10_5 .LUT_INIT=16'b0101000001010001;
    LogicCell40 \POWERLED.func_state_RNI91IA4_0_1_LC_8_10_5  (
            .in0(N__25996),
            .in1(N__27419),
            .in2(N__25963),
            .in3(N__29588),
            .lcout(),
            .ltout(\POWERLED.func_state_RNI91IA4_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI4CHA7_0_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4CHA7_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4CHA7_0_LC_8_10_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.func_state_RNI4CHA7_0_LC_8_10_6  (
            .in0(N__25939),
            .in1(_gnd_net_),
            .in2(N__23401),
            .in3(N__23503),
            .lcout(\POWERLED.func_state_1_m2_0 ),
            .ltout(\POWERLED.func_state_1_m2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIA20K9_0_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIA20K9_0_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIA20K9_0_LC_8_10_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.func_state_RNIA20K9_0_LC_8_10_7  (
            .in0(N__23391),
            .in1(N__30164),
            .in2(N__23383),
            .in3(N__25896),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE1QU7_5_LC_8_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE1QU7_5_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE1QU7_5_LC_8_11_0 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \POWERLED.dutycycle_RNIE1QU7_5_LC_8_11_0  (
            .in0(N__23931),
            .in1(N__23829),
            .in2(N__26308),
            .in3(N__26199),
            .lcout(),
            .ltout(\POWERLED.g0_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILMBVD_5_LC_8_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILMBVD_5_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILMBVD_5_LC_8_11_1 .LUT_INIT=16'b1000000000001010;
    LogicCell40 \POWERLED.dutycycle_RNILMBVD_5_LC_8_11_1  (
            .in0(N__23887),
            .in1(N__29678),
            .in2(N__23713),
            .in3(N__26304),
            .lcout(),
            .ltout(\POWERLED.dutycycle_fb_15_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1DAA11_5_LC_8_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1DAA11_5_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1DAA11_5_LC_8_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI1DAA11_5_LC_8_11_2  (
            .in0(N__23542),
            .in1(N__23707),
            .in2(N__23710),
            .in3(N__23566),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBQG35_5_LC_8_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBQG35_5_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBQG35_5_LC_8_11_3 .LUT_INIT=16'b0011101100001010;
    LogicCell40 \POWERLED.dutycycle_RNIBQG35_5_LC_8_11_3  (
            .in0(N__23806),
            .in1(N__23577),
            .in2(N__24019),
            .in3(N__23828),
            .lcout(\POWERLED.dutycycle_fb_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_5_LC_8_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_0_5_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_5_LC_8_11_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \POWERLED.dutycycle_RNO_0_5_LC_8_11_4  (
            .in0(N__23576),
            .in1(N__26689),
            .in2(_gnd_net_),
            .in3(N__23992),
            .lcout(),
            .ltout(\POWERLED.dutycycle_en_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_8_11_5 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_8_11_5 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \POWERLED.dutycycle_5_LC_8_11_5  (
            .in0(N__26690),
            .in1(N__23826),
            .in2(N__23701),
            .in3(N__23930),
            .lcout(\POWERLED.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34458),
            .ce(),
            .sr(N__23616));
    defparam \POWERLED.dutycycle_RNIN2958_5_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN2958_5_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN2958_5_LC_8_11_6 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \POWERLED.dutycycle_RNIN2958_5_LC_8_11_6  (
            .in0(N__23578),
            .in1(N__24018),
            .in2(N__23917),
            .in3(N__26691),
            .lcout(\POWERLED.dutycycle_fb_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIAP426_5_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIAP426_5_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIAP426_5_LC_8_11_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \POWERLED.dutycycle_RNIAP426_5_LC_8_11_7  (
            .in0(N__23557),
            .in1(N__23551),
            .in2(N__24040),
            .in3(N__23827),
            .lcout(\POWERLED.dutycycle_fb_15_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_2_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_2_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_2_LC_8_12_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_0_2_LC_8_12_0  (
            .in0(N__23533),
            .in1(N__28941),
            .in2(N__29068),
            .in3(N__31163),
            .lcout(\POWERLED.N_340 ),
            .ltout(\POWERLED.N_340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRAVV2_0_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRAVV2_0_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRAVV2_0_LC_8_12_1 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \POWERLED.func_state_RNIRAVV2_0_LC_8_12_1  (
            .in0(N__26002),
            .in1(N__29589),
            .in2(N__23506),
            .in3(N__26113),
            .lcout(\POWERLED.func_state_RNIRAVV2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKLAF2_0_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKLAF2_0_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKLAF2_0_LC_8_12_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNIKLAF2_0_LC_8_12_2  (
            .in0(N__24312),
            .in1(N__24052),
            .in2(N__31167),
            .in3(N__23932),
            .lcout(\POWERLED.dutycycle_fb_15_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_6_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_8_12_3 .LUT_INIT=16'b0000000010111111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_6_LC_8_12_3  (
            .in0(N__26545),
            .in1(N__23880),
            .in2(N__27144),
            .in3(N__24313),
            .lcout(\POWERLED.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILP0F_0_0_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILP0F_0_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILP0F_0_0_LC_8_12_4 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \POWERLED.dutycycle_RNILP0F_0_0_LC_8_12_4  (
            .in0(N__24331),
            .in1(N__23896),
            .in2(N__32967),
            .in3(N__31164),
            .lcout(\POWERLED.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_LC_8_12_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_LC_8_12_5  (
            .in0(N__24083),
            .in1(N__23879),
            .in2(_gnd_net_),
            .in3(N__27110),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_6_LC_8_12_7  (
            .in0(N__24084),
            .in1(N__24217),
            .in2(N__27143),
            .in3(N__26516),
            .lcout(\POWERLED.func_state_1_m2s2_i_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8OIL_5_LC_8_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8OIL_5_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8OIL_5_LC_8_13_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.dutycycle_RNI8OIL_5_LC_8_13_0  (
            .in0(N__24306),
            .in1(N__24051),
            .in2(N__23836),
            .in3(N__31147),
            .lcout(\POWERLED.dutycycle_fb_14_a4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNINH5P1_2_LC_8_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNINH5P1_2_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNINH5P1_2_LC_8_13_1 .LUT_INIT=16'b1100010111001111;
    LogicCell40 \POWERLED.dutycycle_RNINH5P1_2_LC_8_13_1  (
            .in0(N__23719),
            .in1(N__24292),
            .in2(N__31165),
            .in3(N__23758),
            .lcout(\POWERLED.dutycycle_RNINH5P1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_2_0_LC_8_13_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_2_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_2_0_LC_8_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_2_0_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(N__30003),
            .in2(_gnd_net_),
            .in3(N__29460),
            .lcout(\POWERLED.count_off_1_sqmuxa ),
            .ltout(\POWERLED.count_off_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4G9K2_5_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4G9K2_5_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4G9K2_5_LC_8_13_3 .LUT_INIT=16'b1111000000100010;
    LogicCell40 \POWERLED.dutycycle_RNI4G9K2_5_LC_8_13_3  (
            .in0(N__26577),
            .in1(N__25018),
            .in2(N__24127),
            .in3(N__24124),
            .lcout(\POWERLED.dutycycle_RNI4G9K2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_6_LC_8_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_8_13_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_6_LC_8_13_4  (
            .in0(N__24342),
            .in1(N__32963),
            .in2(_gnd_net_),
            .in3(N__26576),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_6 ),
            .ltout(\POWERLED.dutycycle_RNI_4Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_0_LC_8_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_8_13_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_0_LC_8_13_5  (
            .in0(N__32964),
            .in1(N__24118),
            .in2(N__24088),
            .in3(N__24085),
            .lcout(\POWERLED.dutycycle_RNI_8Z0Z_0 ),
            .ltout(\POWERLED.dutycycle_RNI_8Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_2_5_LC_8_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_2_5_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_2_5_LC_8_13_6 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \POWERLED.dutycycle_RNO_2_5_LC_8_13_6  (
            .in0(N__24036),
            .in1(N__24009),
            .in2(N__23998),
            .in3(N__31145),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNO_2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_1_5_LC_8_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_1_5_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_1_5_LC_8_13_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \POWERLED.dutycycle_RNO_1_5_LC_8_13_7  (
            .in0(N__31146),
            .in1(N__24305),
            .in2(N__23995),
            .in3(N__23938),
            .lcout(\POWERLED.N_240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_4_5_LC_8_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_4_5_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_4_5_LC_8_14_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \POWERLED.dutycycle_RNO_4_5_LC_8_14_0  (
            .in0(N__29479),
            .in1(N__29981),
            .in2(_gnd_net_),
            .in3(N__26474),
            .lcout(\POWERLED.g3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILG3T6_6_LC_8_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILG3T6_6_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILG3T6_6_LC_8_14_1 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \POWERLED.dutycycle_RNILG3T6_6_LC_8_14_1  (
            .in0(N__27001),
            .in1(N__26700),
            .in2(N__24265),
            .in3(N__24190),
            .lcout(\POWERLED.dutycycle_eena_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_5_5_LC_8_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_5_5_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_5_5_LC_8_14_2 .LUT_INIT=16'b0110111000001111;
    LogicCell40 \POWERLED.dutycycle_RNO_5_5_LC_8_14_2  (
            .in0(N__26250),
            .in1(N__26287),
            .in2(N__24184),
            .in3(N__23959),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_3_5_LC_8_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_3_5_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_3_5_LC_8_14_3 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \POWERLED.dutycycle_RNO_3_5_LC_8_14_3  (
            .in0(N__26475),
            .in1(N__23947),
            .in2(N__23941),
            .in3(N__26575),
            .lcout(\POWERLED.dutycycle_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_6_LC_8_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_8_14_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_6_LC_8_14_4  (
            .in0(N__24346),
            .in1(N__24330),
            .in2(_gnd_net_),
            .in3(N__32965),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2O4A1_10_LC_8_14_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2O4A1_10_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2O4A1_10_LC_8_14_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.count_clk_RNI2O4A1_10_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__29982),
            .in2(_gnd_net_),
            .in3(N__32966),
            .lcout(\POWERLED.count_clk_RNI2O4A1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_1_LC_8_14_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_8_14_7 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_8_14_7  (
            .in0(N__29313),
            .in1(N__29478),
            .in2(_gnd_net_),
            .in3(N__26574),
            .lcout(\POWERLED.N_239 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI88TE_0_LC_8_15_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI88TE_0_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI88TE_0_LC_8_15_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \POWERLED.func_state_RNI88TE_0_LC_8_15_4  (
            .in0(N__24286),
            .in1(N__27277),
            .in2(_gnd_net_),
            .in3(N__26397),
            .lcout(\POWERLED.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_8_15_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIMQ0F_1_LC_8_15_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNIMQ0F_1_LC_8_15_6  (
            .in0(N__24253),
            .in1(N__30189),
            .in2(N__24229),
            .in3(N__29302),
            .lcout(\POWERLED.N_272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_6_5_LC_8_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_6_5_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_6_5_LC_8_16_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.dutycycle_RNO_6_5_LC_8_16_7  (
            .in0(N__27264),
            .in1(N__28885),
            .in2(_gnd_net_),
            .in3(N__26387),
            .lcout(\POWERLED.dutycycle_N_3_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISVPK4_0_4_LC_9_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISVPK4_0_4_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISVPK4_0_4_LC_9_1_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \PCH_PWRGD.count_RNISVPK4_0_4_LC_9_1_0  (
            .in0(N__24172),
            .in1(N__24163),
            .in2(N__27858),
            .in3(N__24141),
            .lcout(\PCH_PWRGD.count_1_i_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNI9I942_LC_9_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNI9I942_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNI9I942_LC_9_1_1 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNI9I942_LC_9_1_1  (
            .in0(N__27692),
            .in1(N__28208),
            .in2(N__24145),
            .in3(N__24387),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQSOK4_3_LC_9_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQSOK4_3_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQSOK4_3_LC_9_1_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIQSOK4_3_LC_9_1_2  (
            .in0(N__27780),
            .in1(_gnd_net_),
            .in2(N__24148),
            .in3(N__24379),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(\PCH_PWRGD.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_3_LC_9_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_9_1_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_9_1_3 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_3_LC_9_1_3  (
            .in0(N__27693),
            .in1(N__28210),
            .in2(N__24391),
            .in3(N__24388),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34055),
            .ce(N__27845),
            .sr(N__28228));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIESE42_LC_9_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIESE42_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIESE42_LC_9_1_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNIESE42_LC_9_1_4  (
            .in0(N__28207),
            .in1(N__27691),
            .in2(N__27465),
            .in3(N__24366),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI4CUK4_8_LC_9_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI4CUK4_8_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI4CUK4_8_LC_9_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNI4CUK4_8_LC_9_1_5  (
            .in0(_gnd_net_),
            .in1(N__24358),
            .in2(N__24373),
            .in3(N__27779),
            .lcout(\PCH_PWRGD.countZ0Z_8 ),
            .ltout(\PCH_PWRGD.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_8_LC_9_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_9_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_9_1_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_8_LC_9_1_6  (
            .in0(N__28209),
            .in1(N__27694),
            .in2(N__24370),
            .in3(N__24367),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34055),
            .ce(N__27845),
            .sr(N__28228));
    defparam \PCH_PWRGD.count_9_LC_9_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_9_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_9_1_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_9_LC_9_1_7  (
            .in0(N__27695),
            .in1(N__28211),
            .in2(N__27526),
            .in3(N__27501),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34055),
            .ce(N__27845),
            .sr(N__28228));
    defparam \PCH_PWRGD.count_10_LC_9_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_9_2_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_9_2_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \PCH_PWRGD.count_10_LC_9_2_0  (
            .in0(_gnd_net_),
            .in1(N__24465),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34197),
            .ce(N__27838),
            .sr(N__28217));
    defparam \PCH_PWRGD.count_6_LC_9_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_9_2_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_9_2_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \PCH_PWRGD.count_6_LC_9_2_1  (
            .in0(N__24493),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28216),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34197),
            .ce(N__27838),
            .sr(N__28217));
    defparam \PCH_PWRGD.count_RNIFRFT4_10_LC_9_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFRFT4_10_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFRFT4_10_LC_9_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIFRFT4_10_LC_9_2_2  (
            .in0(N__24477),
            .in1(N__24464),
            .in2(_gnd_net_),
            .in3(N__27802),
            .lcout(\PCH_PWRGD.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_9_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_9_2_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_9_2_3 .LUT_INIT=16'b0000001000001010;
    LogicCell40 \PCH_PWRGD.count_0_LC_9_2_3  (
            .in0(N__24678),
            .in1(N__24669),
            .in2(N__28240),
            .in3(N__27553),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34197),
            .ce(N__27838),
            .sr(N__28217));
    defparam \PCH_PWRGD.count_RNI06SK4_6_LC_9_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI06SK4_6_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI06SK4_6_LC_9_2_4 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \PCH_PWRGD.count_RNI06SK4_6_LC_9_2_4  (
            .in0(N__24502),
            .in1(N__24492),
            .in2(N__28239),
            .in3(N__27803),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(\PCH_PWRGD.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIFRFT4_0_10_LC_9_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFRFT4_0_10_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFRFT4_0_10_LC_9_2_5 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \PCH_PWRGD.count_RNIFRFT4_0_10_LC_9_2_5  (
            .in0(N__27804),
            .in1(N__24478),
            .in2(N__24469),
            .in3(N__24466),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI3VBAE_2_LC_9_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI3VBAE_2_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI3VBAE_2_LC_9_2_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI3VBAE_2_LC_9_2_6  (
            .in0(N__24451),
            .in1(N__24442),
            .in2(N__24427),
            .in3(N__24424),
            .lcout(\PCH_PWRGD.count_1_i_a2_11_0 ),
            .ltout(\PCH_PWRGD.count_1_i_a2_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIM6A821_1_LC_9_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIM6A821_1_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIM6A821_1_LC_9_2_7 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \PCH_PWRGD.count_RNIM6A821_1_LC_9_2_7  (
            .in0(N__24679),
            .in1(N__28212),
            .in2(N__24412),
            .in3(N__27552),
            .lcout(\PCH_PWRGD.count_RNIM6A821Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIO73V1_LC_9_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIO73V1_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIO73V1_LC_9_3_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNIO73V1_LC_9_3_0  (
            .in0(N__28166),
            .in1(N__27921),
            .in2(N__27905),
            .in3(N__27685),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIO32O4_11_LC_9_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIO32O4_11_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIO32O4_11_LC_9_3_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIO32O4_11_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(N__27871),
            .in2(N__24409),
            .in3(N__27805),
            .lcout(\PCH_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_3_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_3_2 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_3_2  (
            .in0(N__30951),
            .in1(_gnd_net_),
            .in2(N__25234),
            .in3(N__25266),
            .lcout(),
            .ltout(N_253_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_11_LC_9_3_3 .C_ON=1'b0;
    defparam \POWERLED.G_11_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_11_LC_9_3_3 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \POWERLED.G_11_LC_9_3_3  (
            .in0(N__24818),
            .in1(N__34839),
            .in2(N__24406),
            .in3(N__25232),
            .lcout(G_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI4EPO41_0_LC_9_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI4EPO41_0_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI4EPO41_0_LC_9_3_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNI4EPO41_0_LC_9_3_4  (
            .in0(N__27806),
            .in1(N__24403),
            .in2(_gnd_net_),
            .in3(N__24397),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(\PCH_PWRGD.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI_0_LC_9_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI_0_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI_0_LC_9_3_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.count_RNI_0_LC_9_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24682),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2173_i ),
            .ltout(\PCH_PWRGD.N_2173_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI63UG01_1_LC_9_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI63UG01_1_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI63UG01_1_LC_9_3_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI63UG01_1_LC_9_3_6  (
            .in0(_gnd_net_),
            .in1(N__24670),
            .in2(N__24658),
            .in3(N__27551),
            .lcout(\PCH_PWRGD.N_364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_9_3_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_9_3_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_9_3_7 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_9_3_7  (
            .in0(N__25267),
            .in1(N__30950),
            .in2(N__24825),
            .in3(N__25233),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34069),
            .ce(N__34687),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_9_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_9_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28376),
            .lcout(\PCH_PWRGD.N_2171_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_11_LC_9_4_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_11_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_11_LC_9_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_11_LC_9_4_1  (
            .in0(N__24654),
            .in1(N__24642),
            .in2(N__25273),
            .in3(N__24630),
            .lcout(),
            .ltout(\RSMRST_PWRGD.m4_0_a2_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_LC_9_4_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_LC_9_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_LC_9_4_2  (
            .in0(N__24565),
            .in1(N__24508),
            .in2(N__24619),
            .in3(N__24730),
            .lcout(N_382),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_10_LC_9_4_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_10_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_10_LC_9_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_10_LC_9_4_3  (
            .in0(N__24615),
            .in1(N__24603),
            .in2(N__24592),
            .in3(N__24576),
            .lcout(\RSMRST_PWRGD.m4_0_a2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_9_LC_9_4_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_9_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_9_LC_9_4_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_9_LC_9_4_4  (
            .in0(N__24558),
            .in1(N__24546),
            .in2(N__24535),
            .in3(N__24519),
            .lcout(\RSMRST_PWRGD.m4_0_a2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_12_LC_9_4_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_12_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_12_LC_9_4_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a2_12_LC_9_4_5  (
            .in0(N__24780),
            .in1(N__24768),
            .in2(N__24757),
            .in3(N__24741),
            .lcout(\RSMRST_PWRGD.m4_0_a2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_5_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_5_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_5_0  (
            .in0(N__32172),
            .in1(N__31988),
            .in2(N__28557),
            .in3(N__31798),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_5_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_5_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__24955),
            .in2(N__24724),
            .in3(N__31620),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_9_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_9_5_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_9_5_3  (
            .in0(N__28333),
            .in1(N__28270),
            .in2(_gnd_net_),
            .in3(N__24720),
            .lcout(\PCH_PWRGD.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34294),
            .ce(N__30778),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_9_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_9_5_4 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_9_5_4  (
            .in0(N__24721),
            .in1(N__28271),
            .in2(_gnd_net_),
            .in3(N__28332),
            .lcout(),
            .ltout(\PCH_PWRGD.m4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI0EA52_0_LC_9_5_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI0EA52_0_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI0EA52_0_LC_9_5_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNI0EA52_0_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__24694),
            .in2(N__24688),
            .in3(N__30531),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_6_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_6_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_6_0  (
            .in0(N__32166),
            .in1(N__31790),
            .in2(N__30850),
            .in3(N__31980),
            .lcout(\VPP_VDDQ.count_2_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_9_6_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_9_6_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_9_6_1  (
            .in0(N__31791),
            .in1(N__32167),
            .in2(N__28599),
            .in3(N__31981),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_9_6_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIPM861_8_LC_9_6_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIPM861_8_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__24970),
            .in2(N__24685),
            .in3(N__31626),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_8_LC_9_6_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_8_LC_9_6_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_9_6_3  (
            .in0(N__31794),
            .in1(N__32171),
            .in2(N__28600),
            .in3(N__31984),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34210),
            .ce(N__31631),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_9_6_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_9_LC_9_6_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_9_6_4  (
            .in0(N__32169),
            .in1(N__31795),
            .in2(N__31990),
            .in3(N__28578),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34210),
            .ce(N__31631),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_6_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_6_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_6_5  (
            .in0(N__31792),
            .in1(N__32168),
            .in2(N__28579),
            .in3(N__31982),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_9_6_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIRP961_9_LC_9_6_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIRP961_9_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__24964),
            .in2(N__24958),
            .in3(N__31627),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_10_LC_9_6_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_10_LC_9_6_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_9_6_7  (
            .in0(N__31793),
            .in1(N__32170),
            .in2(N__28558),
            .in3(N__31983),
            .lcout(\VPP_VDDQ.count_2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34210),
            .ce(N__31631),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_9_7_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_9_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_9_7_1  (
            .in0(N__24935),
            .in1(N__24901),
            .in2(N__24882),
            .in3(N__24855),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(rsmrst_pwrgd_signal_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a3_0_LC_9_7_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a3_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a3_0_LC_9_7_2 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_a3_0_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__25208),
            .in2(N__24832),
            .in3(N__25269),
            .lcout(),
            .ltout(\RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_9_7_3 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_9_7_3  (
            .in0(N__25209),
            .in1(_gnd_net_),
            .in2(N__24829),
            .in3(N__24826),
            .lcout(RSMRST_PWRGD_curr_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34161),
            .ce(N__34696),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_7_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_7_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_7_4  (
            .in0(N__30941),
            .in1(N__25207),
            .in2(_gnd_net_),
            .in3(N__25268),
            .lcout(\RSMRST_PWRGD.N_254_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_7_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_7_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_7_5  (
            .in0(N__25271),
            .in1(_gnd_net_),
            .in2(N__25221),
            .in3(N__30940),
            .lcout(RSMRSTn_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34161),
            .ce(N__34696),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_7_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_7_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_7_6  (
            .in0(N__30939),
            .in1(N__25210),
            .in2(_gnd_net_),
            .in3(N__25272),
            .lcout(RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34161),
            .ce(N__34696),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_7_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_LC_9_7_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_LC_9_7_7  (
            .in0(N__25270),
            .in1(_gnd_net_),
            .in2(N__25220),
            .in3(N__30938),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34161),
            .ce(N__34696),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIU2UT_1_LC_9_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIU2UT_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIU2UT_1_LC_9_8_0 .LUT_INIT=16'b0011100000000000;
    LogicCell40 \POWERLED.func_state_RNIU2UT_1_LC_9_8_0  (
            .in0(N__26352),
            .in1(N__28960),
            .in2(N__31108),
            .in3(N__26617),
            .lcout(\POWERLED.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_en_LC_9_8_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_en_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_en_LC_9_8_1 .LUT_INIT=16'b1011111100000000;
    LogicCell40 \POWERLED.func_state_en_LC_9_8_1  (
            .in0(N__28961),
            .in1(N__26351),
            .in2(N__27349),
            .in3(N__29758),
            .lcout(\POWERLED.func_state_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_8_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_8_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__34840),
            .in2(_gnd_net_),
            .in3(N__25172),
            .lcout(\RSMRST_PWRGD.N_29_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_0_LC_9_8_3 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_0_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_0_LC_9_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.VCCST_EN_0_LC_9_8_3  (
            .in0(N__28958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26970),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_0_LC_9_8_5 .C_ON=1'b0;
    defparam \COUNTER.tmp_0_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_0_LC_9_8_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_0_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__30490),
            .in2(_gnd_net_),
            .in3(N__25121),
            .lcout(suswarn_n),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34328),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_m1_e_LC_9_8_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_m1_e_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_m1_e_LC_9_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.dutycycle_m1_e_LC_9_8_6  (
            .in0(N__27341),
            .in1(N__28959),
            .in2(_gnd_net_),
            .in3(N__26068),
            .lcout(\POWERLED.dutycycle_N_3_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIRCVD_7_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__25789),
            .in2(N__32305),
            .in3(N__33318),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_9_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_9_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_7_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32304),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34332),
            .ce(N__33332),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIVI1E_9_LC_9_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIVI1E_9_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIVI1E_9_LC_9_9_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIVI1E_9_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__25783),
            .in2(N__32284),
            .in3(N__33319),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_9_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_9_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_9_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32283),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34332),
            .ce(N__33332),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI17P1A_5_LC_9_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI17P1A_5_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI17P1A_5_LC_9_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNI17P1A_5_LC_9_9_4  (
            .in0(N__25777),
            .in1(N__25759),
            .in2(_gnd_net_),
            .in3(N__25569),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI3AQ1A_6_LC_9_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI3AQ1A_6_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI3AQ1A_6_LC_9_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNI3AQ1A_6_LC_9_9_5  (
            .in0(N__25570),
            .in1(N__25708),
            .in2(_gnd_net_),
            .in3(N__25690),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIRTL1A_2_LC_9_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIRTL1A_2_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIRTL1A_2_LC_9_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIRTL1A_2_LC_9_9_6  (
            .in0(N__25642),
            .in1(N__25624),
            .in2(_gnd_net_),
            .in3(N__25568),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_15_LC_9_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_9_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_1_15_LC_9_9_7  (
            .in0(N__25435),
            .in1(N__25371),
            .in2(_gnd_net_),
            .in3(N__25306),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_1_2_LC_9_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_1_2_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_1_2_LC_9_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_1_2_LC_9_10_0  (
            .in0(N__28980),
            .in1(N__29051),
            .in2(_gnd_net_),
            .in3(N__31139),
            .lcout(\POWERLED.N_340_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_9_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_9_10_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \POWERLED.func_state_1_LC_9_10_1  (
            .in0(N__25895),
            .in1(N__25915),
            .in2(N__30188),
            .in3(N__25921),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34361),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2O4A1_0_0_LC_9_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2O4A1_0_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2O4A1_0_0_LC_9_10_3 .LUT_INIT=16'b0000000011011111;
    LogicCell40 \POWERLED.func_state_RNI2O4A1_0_0_LC_9_10_3  (
            .in0(N__26074),
            .in1(N__28981),
            .in2(N__27334),
            .in3(N__30051),
            .lcout(\POWERLED.N_4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI91IA4_1_LC_9_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI91IA4_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI91IA4_1_LC_9_10_4 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \POWERLED.func_state_RNI91IA4_1_LC_9_10_4  (
            .in0(N__25997),
            .in1(N__27421),
            .in2(N__25962),
            .in3(N__29587),
            .lcout(),
            .ltout(\POWERLED.func_state_RNI91IA4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIKML48_1_LC_9_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIKML48_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIKML48_1_LC_9_10_5 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \POWERLED.func_state_RNIKML48_1_LC_9_10_5  (
            .in0(N__26626),
            .in1(N__25938),
            .in2(N__25924),
            .in3(_gnd_net_),
            .lcout(\POWERLED.func_state_1_m2_1 ),
            .ltout(\POWERLED.func_state_1_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRD4EA_1_LC_9_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRD4EA_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRD4EA_1_LC_9_10_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \POWERLED.func_state_RNIRD4EA_1_LC_9_10_6  (
            .in0(N__25914),
            .in1(N__30159),
            .in2(N__25906),
            .in3(N__25894),
            .lcout(\POWERLED.func_state ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_9_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_9_10_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_0_LC_9_10_7  (
            .in0(N__30160),
            .in1(N__25848),
            .in2(_gnd_net_),
            .in3(N__29424),
            .lcout(\POWERLED.un1_func_state25_6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_7_1_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_7_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_7_1_LC_9_11_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \POWERLED.func_state_RNI_7_1_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__27422),
            .in2(_gnd_net_),
            .in3(N__32915),
            .lcout(func_state_RNI_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_0_2_LC_9_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_0_2_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_0_2_LC_9_11_1 .LUT_INIT=16'b1011101100110011;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_0_2_LC_9_11_1  (
            .in0(N__26285),
            .in1(N__26295),
            .in2(_gnd_net_),
            .in3(N__26259),
            .lcout(),
            .ltout(N_4_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S3n_RNI75Q52_LC_9_11_2.C_ON=1'b0;
    defparam SLP_S3n_RNI75Q52_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam SLP_S3n_RNI75Q52_LC_9_11_2.LUT_INIT=16'b0100000000000000;
    LogicCell40 SLP_S3n_RNI75Q52_LC_9_11_2 (
            .in0(N__27303),
            .in1(N__28909),
            .in2(N__25792),
            .in3(N__26469),
            .lcout(),
            .ltout(G_34_0_a4_0_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_2_RNIH76R4_LC_9_11_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_2_RNIH76R4_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_2_RNIH76R4_LC_9_11_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_2_RNIH76R4_LC_9_11_3  (
            .in0(N__26353),
            .in1(N__26218),
            .in2(N__26311),
            .in3(N__26422),
            .lcout(POWERLED_un1_dutycycle_172_m3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_1_2_LC_9_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_1_2_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_1_2_LC_9_11_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_1_2_LC_9_11_4  (
            .in0(N__26296),
            .in1(N__26286),
            .in2(N__26263),
            .in3(N__26468),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_9_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_9_11_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.un1_clk_100khz_52_and_i_a2_0_LC_9_11_5  (
            .in0(N__26354),
            .in1(N__28908),
            .in2(_gnd_net_),
            .in3(N__27302),
            .lcout(\POWERLED.N_319_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_9_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_9_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__26147),
            .in2(_gnd_net_),
            .in3(N__29223),
            .lcout(\POWERLED.func_state_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3VDK_0_LC_9_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3VDK_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3VDK_0_LC_9_11_7 .LUT_INIT=16'b0111010000000000;
    LogicCell40 \POWERLED.func_state_RNI3VDK_0_LC_9_11_7  (
            .in0(N__30491),
            .in1(N__31133),
            .in2(N__26157),
            .in3(N__29626),
            .lcout(\POWERLED.N_297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIBVNS_1_LC_9_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIBVNS_1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIBVNS_1_LC_9_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_clk_RNIBVNS_1_LC_9_12_0  (
            .in0(N__28755),
            .in1(N__32494),
            .in2(N__28827),
            .in3(N__29504),
            .lcout(\POWERLED.N_284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_2_LC_9_12_1 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_2_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_2_LC_9_12_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_2_LC_9_12_1  (
            .in0(N__32496),
            .in1(N__28756),
            .in2(N__28820),
            .in3(N__29246),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_o_N_296_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_12_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_9_12_2  (
            .in0(N__26107),
            .in1(N__26785),
            .in2(N__26098),
            .in3(N__29625),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_9_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_9_12_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_9_12_3  (
            .in0(N__26815),
            .in1(N__27428),
            .in2(N__26095),
            .in3(N__29582),
            .lcout(\POWERLED.un1_func_state25_6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI0RLE1_8_LC_9_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI0RLE1_8_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI0RLE1_8_LC_9_12_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \POWERLED.count_clk_RNI0RLE1_8_LC_9_12_4  (
            .in0(N__26946),
            .in1(_gnd_net_),
            .in2(N__29593),
            .in3(N__32497),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBQDB2_0_LC_9_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBQDB2_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBQDB2_0_LC_9_12_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \POWERLED.func_state_RNIBQDB2_0_LC_9_12_5  (
            .in0(N__26803),
            .in1(N__29115),
            .in2(N__26929),
            .in3(N__26926),
            .lcout(\POWERLED.func_state_RNIBQDB2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_9_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_9_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_9_12_6  (
            .in0(N__29116),
            .in1(N__26814),
            .in2(N__26802),
            .in3(N__32495),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_294_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBL3Q3_1_LC_9_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBL3Q3_1_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBL3Q3_1_LC_9_12_7 .LUT_INIT=16'b0000101000111011;
    LogicCell40 \POWERLED.func_state_RNIBL3Q3_1_LC_9_12_7  (
            .in0(N__29505),
            .in1(N__26779),
            .in2(N__26759),
            .in3(N__29583),
            .lcout(\POWERLED.func_state_RNIBL3Q3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_0_1_LC_9_13_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_0_1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_0_1_LC_9_13_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \POWERLED.func_state_RNIOGRS_0_1_LC_9_13_0  (
            .in0(N__29303),
            .in1(N__31148),
            .in2(_gnd_net_),
            .in3(N__28957),
            .lcout(\POWERLED.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_9_1_LC_9_13_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_9_1_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_9_1_LC_9_13_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI_9_1_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__29451),
            .in2(_gnd_net_),
            .in3(N__29509),
            .lcout(\POWERLED.func_state_1_m2s2_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2O4A1_5_LC_9_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2O4A1_5_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2O4A1_5_LC_9_13_6 .LUT_INIT=16'b1010101000101010;
    LogicCell40 \POWERLED.dutycycle_RNI2O4A1_5_LC_9_13_6  (
            .in0(N__26578),
            .in1(N__30004),
            .in2(N__29473),
            .in3(N__26456),
            .lcout(N_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIBVNS_0_LC_9_13_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIBVNS_0_LC_9_13_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.func_state_RNIBVNS_0_LC_9_13_7  (
            .in0(N__28956),
            .in1(N__26355),
            .in2(N__27333),
            .in3(N__29447),
            .lcout(\POWERLED.func_state_RNIBVNSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_0_1_LC_9_14_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_0_1_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_0_1_LC_9_14_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \POWERLED.func_state_RNI34G9_0_1_LC_9_14_0  (
            .in0(N__27429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29066),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_a2_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8H551_6_LC_9_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8H551_6_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8H551_6_LC_9_14_1 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \POWERLED.dutycycle_RNI8H551_6_LC_9_14_1  (
            .in0(N__28911),
            .in1(N__27265),
            .in2(N__27187),
            .in3(N__27163),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_a2_6_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIRKB61_6_LC_9_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIRKB61_6_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIRKB61_6_LC_9_14_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIRKB61_6_LC_9_14_2  (
            .in0(N__26981),
            .in1(_gnd_net_),
            .in2(N__27184),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_309_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPUGO_0_1_LC_9_14_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPUGO_0_1_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPUGO_0_1_LC_9_14_3 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \POWERLED.func_state_RNIPUGO_0_1_LC_9_14_3  (
            .in0(N__28912),
            .in1(N__26992),
            .in2(_gnd_net_),
            .in3(N__26982),
            .lcout(),
            .ltout(\POWERLED.func_state_RNIPUGO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI7N202_1_LC_9_14_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI7N202_1_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI7N202_1_LC_9_14_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.func_state_RNI7N202_1_LC_9_14_4  (
            .in0(N__31149),
            .in1(_gnd_net_),
            .in2(N__27181),
            .in3(N__26953),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_o2_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI44JG4_6_LC_9_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI44JG4_6_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI44JG4_6_LC_9_14_5 .LUT_INIT=16'b1011111110111011;
    LogicCell40 \POWERLED.dutycycle_RNI44JG4_6_LC_9_14_5  (
            .in0(N__27178),
            .in1(N__27172),
            .in2(N__27166),
            .in3(N__27162),
            .lcout(\POWERLED.N_145_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_1_LC_9_14_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_1_LC_9_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI34G9_1_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__29304),
            .in2(_gnd_net_),
            .in3(N__29067),
            .lcout(\POWERLED.un1_clk_100khz_51_and_i_a2_5_0 ),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPUGO_1_LC_9_14_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPUGO_1_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPUGO_1_LC_9_14_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.func_state_RNIPUGO_1_LC_9_14_7  (
            .in0(N__28913),
            .in1(N__29314),
            .in2(N__26986),
            .in3(N__26983),
            .lcout(\POWERLED.func_state_RNIPUGOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_9_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_9_15_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_9_15_2  (
            .in0(N__30310),
            .in1(N__30260),
            .in2(_gnd_net_),
            .in3(N__30076),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34417),
            .ce(N__34712),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_1_LC_11_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_11_1_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_11_1_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.count_1_LC_11_1_0  (
            .in0(N__28169),
            .in1(N__27624),
            .in2(_gnd_net_),
            .in3(N__27607),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33983),
            .ce(N__27859),
            .sr(N__28170));
    defparam \PCH_PWRGD.count_RNIVBR74_1_LC_11_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIVBR74_1_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIVBR74_1_LC_11_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \PCH_PWRGD.count_RNIVBR74_1_LC_11_1_1  (
            .in0(N__27576),
            .in1(N__27850),
            .in2(_gnd_net_),
            .in3(N__27583),
            .lcout(\PCH_PWRGD.un2_count_1_axb_1 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIG3CN1_1_LC_11_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIG3CN1_1_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIG3CN1_1_LC_11_1_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \PCH_PWRGD.count_RNIG3CN1_1_LC_11_1_2  (
            .in0(N__28168),
            .in1(_gnd_net_),
            .in2(N__27610),
            .in3(N__27606),
            .lcout(\PCH_PWRGD.count_rst_13 ),
            .ltout(\PCH_PWRGD.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIVBR74_0_1_LC_11_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIVBR74_0_1_LC_11_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIVBR74_0_1_LC_11_1_3 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \PCH_PWRGD.count_RNIVBR74_0_1_LC_11_1_3  (
            .in0(N__27577),
            .in1(N__27909),
            .in2(N__27568),
            .in3(N__27852),
            .lcout(),
            .ltout(\PCH_PWRGD.count_1_i_a2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI34I6I_1_LC_11_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI34I6I_1_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI34I6I_1_LC_11_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI34I6I_1_LC_11_1_4  (
            .in0(N__27436),
            .in1(N__27565),
            .in2(N__27556),
            .in3(N__28030),
            .lcout(\PCH_PWRGD.count_1_i_a2_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI6FVK4_9_LC_11_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI6FVK4_9_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI6FVK4_9_LC_11_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNI6FVK4_9_LC_11_1_5  (
            .in0(N__27477),
            .in1(N__27484),
            .in2(_gnd_net_),
            .in3(N__27849),
            .lcout(\PCH_PWRGD.un2_count_1_axb_9 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIFUF42_LC_11_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIFUF42_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIFUF42_LC_11_1_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNIFUF42_LC_11_1_6  (
            .in0(N__28167),
            .in1(N__27505),
            .in2(N__27487),
            .in3(N__27696),
            .lcout(\PCH_PWRGD.count_rst_5 ),
            .ltout(\PCH_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI6FVK4_0_9_LC_11_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI6FVK4_0_9_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI6FVK4_0_9_LC_11_1_7 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \PCH_PWRGD.count_RNI6FVK4_0_9_LC_11_1_7  (
            .in0(N__27478),
            .in1(N__27466),
            .in2(N__27439),
            .in3(N__27851),
            .lcout(\PCH_PWRGD.count_1_i_a2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI29TK4_7_LC_11_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI29TK4_7_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI29TK4_7_LC_11_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNI29TK4_7_LC_11_2_0  (
            .in0(N__28039),
            .in1(N__27985),
            .in2(_gnd_net_),
            .in3(N__27820),
            .lcout(\PCH_PWRGD.un2_count_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIDQD42_LC_11_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIDQD42_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIDQD42_LC_11_2_1 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNIDQD42_LC_11_2_1  (
            .in0(N__27701),
            .in1(N__28024),
            .in2(N__28235),
            .in3(N__28002),
            .lcout(\PCH_PWRGD.count_rst_7 ),
            .ltout(\PCH_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI29TK4_0_7_LC_11_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI29TK4_0_7_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI29TK4_0_7_LC_11_2_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \PCH_PWRGD.count_RNI29TK4_0_7_LC_11_2_2  (
            .in0(N__27857),
            .in1(N__27984),
            .in2(N__28033),
            .in3(N__27965),
            .lcout(\PCH_PWRGD.count_1_i_a2_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_7_LC_11_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_11_2_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_11_2_3 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.count_7_LC_11_2_3  (
            .in0(N__27699),
            .in1(N__28023),
            .in2(N__28234),
            .in3(N__28001),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34275),
            .ce(N__27856),
            .sr(N__28241));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIBMB42_LC_11_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIBMB42_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIBMB42_LC_11_2_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNIBMB42_LC_11_2_4  (
            .in0(N__28083),
            .in1(N__27966),
            .in2(N__27952),
            .in3(N__27700),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIU2RK4_5_LC_11_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIU2RK4_5_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIU2RK4_5_LC_11_2_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PCH_PWRGD.count_RNIU2RK4_5_LC_11_2_5  (
            .in0(N__27931),
            .in1(_gnd_net_),
            .in2(N__27976),
            .in3(N__27821),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(\PCH_PWRGD.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_5_LC_11_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_11_2_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_11_2_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_5_LC_11_2_6  (
            .in0(N__27948),
            .in1(N__28193),
            .in2(N__27934),
            .in3(N__27698),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34275),
            .ce(N__27856),
            .sr(N__28241));
    defparam \PCH_PWRGD.count_11_LC_11_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_11_2_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_11_2_7 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.count_11_LC_11_2_7  (
            .in0(N__27697),
            .in1(N__27925),
            .in2(N__27910),
            .in3(N__28242),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34275),
            .ce(N__27856),
            .sr(N__28241));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_a2_LC_11_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_a2_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_a2_LC_11_3_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_i_a2_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__28309),
            .in2(_gnd_net_),
            .in3(N__27670),
            .lcout(G_1939),
            .ltout(G_1939_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_11_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_11_3_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28387),
            .in3(N__28353),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34292),
            .ce(N__30779),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_o3_0_LC_11_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_o3_0_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_i_o3_0_LC_11_3_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_i_o3_0_LC_11_3_3  (
            .in0(N__31254),
            .in1(N__28290),
            .in2(_gnd_net_),
            .in3(N__28383),
            .lcout(N_218),
            .ltout(N_218_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_11_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_11_3_4 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_11_3_4  (
            .in0(N__28339),
            .in1(N__28326),
            .in2(N__28312),
            .in3(N__30575),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(\PCH_PWRGD.curr_state_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_0_1_LC_11_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_0_1_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIVGBJ_0_1_LC_11_3_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.curr_state_RNIVGBJ_0_1_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28303),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2190_i ),
            .ltout(\PCH_PWRGD.N_2190_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIG3CN1_1_LC_11_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIG3CN1_1_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIG3CN1_1_LC_11_3_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIG3CN1_1_LC_11_3_6  (
            .in0(N__28279),
            .in1(N__31253),
            .in2(N__28246),
            .in3(N__30576),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_0_LC_11_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_11_4_0 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_11_4_0  (
            .in0(N__31777),
            .in1(N__32069),
            .in2(N__30411),
            .in3(N__31908),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34374),
            .ce(N__30780),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_1_LC_11_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_11_4_1 .LUT_INIT=16'b0000010001010100;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_11_4_1  (
            .in0(N__31907),
            .in1(N__30406),
            .in2(N__32111),
            .in3(N__31778),
            .lcout(\VPP_VDDQ.curr_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34374),
            .ce(N__30780),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_4_2 .LUT_INIT=16'b1100111101110111;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_4_2  (
            .in0(N__31775),
            .in1(N__32068),
            .in2(N__30412),
            .in3(N__31909),
            .lcout(),
            .ltout(\VPP_VDDQ.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_4_3 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__28048),
            .in2(N__28042),
            .in3(N__30547),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_11_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_11_4_4 .LUT_INIT=16'b1111101011110011;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_11_4_4  (
            .in0(N__31774),
            .in1(N__30410),
            .in2(N__28417),
            .in3(N__32073),
            .lcout(),
            .ltout(\VPP_VDDQ.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_11_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_11_4_5 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__28414),
            .in2(N__28408),
            .in3(N__30546),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_4_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_4_6  (
            .in0(N__31776),
            .in1(N__28444),
            .in2(N__28405),
            .in3(N__31906),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_11_4_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIF7361_3_LC_11_4_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIF7361_3_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(N__28486),
            .in2(N__28402),
            .in3(N__31549),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_11_5_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_2_LC_11_5_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_11_5_0  (
            .in0(N__31744),
            .in1(N__28473),
            .in2(N__31953),
            .in3(N__32086),
            .lcout(\VPP_VDDQ.count_2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34378),
            .ce(N__31621),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_11_5_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_11_5_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_11_5_1  (
            .in0(N__32083),
            .in1(N__31901),
            .in2(N__28474),
            .in3(N__31742),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_11_5_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNID4261_2_LC_11_5_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNID4261_2_LC_11_5_2  (
            .in0(N__31547),
            .in1(_gnd_net_),
            .in2(N__28399),
            .in3(N__28396),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_2_LC_11_5_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_2_LC_11_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI_2_LC_11_5_3  (
            .in0(N__28621),
            .in1(N__31297),
            .in2(N__28390),
            .in3(N__28458),
            .lcout(\VPP_VDDQ.un9_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_11_5_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_15_LC_11_5_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_11_5_4  (
            .in0(N__31743),
            .in1(N__32085),
            .in2(N__28510),
            .in3(N__31927),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34378),
            .ce(N__31621),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_5_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_5_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_11_5_5  (
            .in0(N__32087),
            .in1(N__28509),
            .in2(N__31972),
            .in3(N__31745),
            .lcout(),
            .ltout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_11_5_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIL79C1_15_LC_11_5_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIL79C1_15_LC_11_5_6  (
            .in0(N__31548),
            .in1(_gnd_net_),
            .in2(N__28495),
            .in3(N__28492),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_11_5_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_3_LC_11_5_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_11_5_7  (
            .in0(N__32084),
            .in1(N__31902),
            .in2(N__31797),
            .in3(N__28443),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34378),
            .ce(N__31621),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_6_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__32248),
            .in2(N__32236),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_6_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__28480),
            .in2(_gnd_net_),
            .in3(N__28462),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_6_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__28459),
            .in2(_gnd_net_),
            .in3(N__28429),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_6_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__30891),
            .in2(_gnd_net_),
            .in3(N__28426),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_6_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__31296),
            .in2(_gnd_net_),
            .in3(N__28423),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_11_6_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_11_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__30898),
            .in2(_gnd_net_),
            .in3(N__28420),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_6_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__28666),
            .in2(_gnd_net_),
            .in3(N__28624),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_6_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__28617),
            .in2(_gnd_net_),
            .in3(N__28582),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_7_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__28716),
            .in2(_gnd_net_),
            .in3(N__28561),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_7_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__28689),
            .in2(_gnd_net_),
            .in3(N__28528),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_7_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__31480),
            .in2(_gnd_net_),
            .in3(N__28525),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_7_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__31428),
            .in2(_gnd_net_),
            .in3(N__28522),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_7_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__31453),
            .in2(_gnd_net_),
            .in3(N__28519),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_7_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__31410),
            .in2(_gnd_net_),
            .in3(N__28516),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_11_7_6  (
            .in0(N__31446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28513),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_7_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_7_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_11_7_7  (
            .in0(N__32164),
            .in1(N__31952),
            .in2(N__31365),
            .in3(N__31766),
            .lcout(\VPP_VDDQ.count_2_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_11_8_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_11_8_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_11_8_0  (
            .in0(N__31949),
            .in1(N__28656),
            .in2(N__32181),
            .in3(N__31784),
            .lcout(\VPP_VDDQ.count_2_1_7 ),
            .ltout(\VPP_VDDQ.count_2_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_11_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_0_7_LC_11_8_1 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_0_7_LC_11_8_1  (
            .in0(N__31606),
            .in1(N__28645),
            .in2(N__28720),
            .in3(N__28717),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_11_8_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_1_7_LC_11_8_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_1_7_LC_11_8_2  (
            .in0(N__31393),
            .in1(N__31479),
            .in2(N__28693),
            .in3(N__28690),
            .lcout(\VPP_VDDQ.un9_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_11_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINJ761_7_LC_11_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNINJ761_7_LC_11_8_3  (
            .in0(N__31605),
            .in1(N__28644),
            .in2(_gnd_net_),
            .in3(N__28672),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_11_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_7_LC_11_8_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_11_8_4  (
            .in0(N__31950),
            .in1(N__28657),
            .in2(N__32182),
            .in3(N__31786),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34434),
            .ce(N__31632),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_0_LC_11_8_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_0_LC_11_8_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \VPP_VDDQ.count_2_RNI_0_LC_11_8_5  (
            .in0(N__31783),
            .in1(N__32173),
            .in2(N__32235),
            .in3(N__31948),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_11_8_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIT1QU_0_LC_11_8_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIT1QU_0_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__31604),
            .in2(N__28636),
            .in3(N__28630),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_0_LC_11_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_0_LC_11_8_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_11_8_7  (
            .in0(N__31785),
            .in1(N__32177),
            .in2(N__28633),
            .in3(N__31951),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34434),
            .ce(N__31632),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJ0RD_3_LC_11_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJ0RD_3_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJ0RD_3_LC_11_9_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.count_clk_RNIJ0RD_3_LC_11_9_0  (
            .in0(N__28741),
            .in1(N__33289),
            .in2(N__33488),
            .in3(N__32349),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_11_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_11_9_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_3_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__33475),
            .in2(_gnd_net_),
            .in3(N__32350),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33999),
            .ce(N__33324),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_11_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_11_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_clk_13_LC_11_9_2  (
            .in0(N__32455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33483),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33999),
            .ce(N__33324),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINA66_14_LC_11_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINA66_14_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINA66_14_LC_11_9_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \POWERLED.count_clk_RNINA66_14_LC_11_9_3  (
            .in0(N__33291),
            .in1(N__28726),
            .in2(N__33490),
            .in3(N__32433),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(\POWERLED.count_clkZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_13_LC_11_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_13_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_13_LC_11_9_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.count_clk_RNI_13_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28735),
            .in3(N__32469),
            .lcout(\POWERLED.count_clk_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIL756_13_LC_11_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIL756_13_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIL756_13_LC_11_9_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \POWERLED.count_clk_RNIL756_13_LC_11_9_5  (
            .in0(N__33290),
            .in1(N__28732),
            .in2(N__33489),
            .in3(N__32454),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_11_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_clk_14_LC_11_9_6  (
            .in0(N__32434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33484),
            .lcout(\POWERLED.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33999),
            .ce(N__33324),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_11_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_11_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_4_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__33476),
            .in2(_gnd_net_),
            .in3(N__32335),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__33999),
            .ce(N__33324),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_11_10_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_11_10_0  (
            .in0(N__32613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33411),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNI_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIQF8B_0_LC_11_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIQF8B_0_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIQF8B_0_LC_11_10_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIQF8B_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__28762),
            .in2(N__28786),
            .in3(N__33285),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(\POWERLED.count_clkZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_11_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_11_10_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__33019),
            .in2(N__28783),
            .in3(N__33412),
            .lcout(),
            .ltout(\POWERLED.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIRG8B_1_LC_11_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIRG8B_1_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIRG8B_1_LC_11_10_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_clk_RNIRG8B_1_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__32587),
            .in2(N__28780),
            .in3(N__33286),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIP9UD_6_LC_11_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIP9UD_6_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIP9UD_6_LC_11_10_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \POWERLED.count_clk_RNIP9UD_6_LC_11_10_4  (
            .in0(N__33288),
            .in1(N__33416),
            .in2(N__28771),
            .in3(N__32316),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIL3SD_4_LC_11_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIL3SD_4_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIL3SD_4_LC_11_10_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \POWERLED.count_clk_RNIL3SD_4_LC_11_10_5  (
            .in0(N__28777),
            .in1(N__33287),
            .in2(N__33458),
            .in3(N__32334),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_11_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_6_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__32317),
            .in2(_gnd_net_),
            .in3(N__33418),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34438),
            .ce(N__33317),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_11_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_11_10_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_clk_0_LC_11_10_7  (
            .in0(N__33417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32612),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34438),
            .ce(N__33317),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_1_LC_11_11_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_1_LC_11_11_0  (
            .in0(N__32823),
            .in1(N__32735),
            .in2(N__33024),
            .in3(N__32414),
            .lcout(\POWERLED.count_clk_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_11_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_11_11_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_11_11_1  (
            .in0(N__32413),
            .in1(N__33014),
            .in2(N__32737),
            .in3(N__32822),
            .lcout(\POWERLED.count_clk_RNIZ0Z_1 ),
            .ltout(\POWERLED.count_clk_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_11_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_11_11_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_11_11_2  (
            .in0(N__29322),
            .in1(_gnd_net_),
            .in2(N__29119),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_1_1_LC_11_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_1_1_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_1_1_LC_11_11_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.func_state_RNIOGRS_1_1_LC_11_11_3  (
            .in0(N__31114),
            .in1(N__29109),
            .in2(N__29095),
            .in3(N__28910),
            .lcout(\POWERLED.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_4_LC_11_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_4_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_4_LC_11_11_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \POWERLED.count_clk_RNI_4_LC_11_11_4  (
            .in0(N__32540),
            .in1(N__33539),
            .in2(N__32418),
            .in3(N__32514),
            .lcout(\POWERLED.un2_count_clk_15_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI18EF2_1_LC_11_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI18EF2_1_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI18EF2_1_LC_11_11_5 .LUT_INIT=16'b1111111110101011;
    LogicCell40 \POWERLED.func_state_RNI18EF2_1_LC_11_11_5  (
            .in0(N__29092),
            .in1(N__30228),
            .in2(N__31153),
            .in3(N__29621),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIH9594_1_LC_11_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIH9594_1_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIH9594_1_LC_11_11_6 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \POWERLED.func_state_RNIH9594_1_LC_11_11_6  (
            .in0(N__29155),
            .in1(N__29077),
            .in2(N__29071),
            .in3(N__32484),
            .lcout(\POWERLED.func_state_RNIH9594_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOTGO_1_LC_11_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOTGO_1_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOTGO_1_LC_11_12_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.func_state_RNIOTGO_1_LC_11_12_0  (
            .in0(N__29591),
            .in1(N__29050),
            .in2(N__29334),
            .in3(N__31110),
            .lcout(\POWERLED.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_0_LC_11_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_0_LC_11_12_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.func_state_RNI34G9_0_LC_11_12_1  (
            .in0(N__29049),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29488),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_4_i_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIRKB61_1_LC_11_12_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIRKB61_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIRKB61_1_LC_11_12_2 .LUT_INIT=16'b0100110011111111;
    LogicCell40 \POWERLED.func_state_RNIRKB61_1_LC_11_12_2  (
            .in0(N__29518),
            .in1(N__28955),
            .in2(N__28831),
            .in3(N__31109),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIUHKR2_1_LC_11_12_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIUHKR2_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIUHKR2_1_LC_11_12_3 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \POWERLED.func_state_RNIUHKR2_1_LC_11_12_3  (
            .in0(N__28828),
            .in1(N__28795),
            .in2(N__28789),
            .in3(N__29620),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1U3S4_1_LC_11_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1U3S4_1_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1U3S4_1_LC_11_12_4 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \POWERLED.func_state_RNI1U3S4_1_LC_11_12_4  (
            .in0(N__30055),
            .in1(N__30002),
            .in2(N__29833),
            .in3(N__29713),
            .lcout(\POWERLED.count_clk_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_1_LC_11_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_1_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_1_LC_11_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.func_state_RNI_2_1_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29329),
            .in3(N__29590),
            .lcout(\POWERLED.func_state_RNI_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_11_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_11_12_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_11_12_6  (
            .in0(N__29592),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29294),
            .lcout(\POWERLED.N_176 ),
            .ltout(\POWERLED.N_176_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_1_LC_11_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_1_LC_11_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.func_state_RNI_5_1_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29512),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_2218_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOGRS_1_LC_11_13_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOGRS_1_LC_11_13_0 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \POWERLED.func_state_RNIOGRS_1_LC_11_13_0  (
            .in0(N__29480),
            .in1(N__29344),
            .in2(N__29335),
            .in3(N__32882),
            .lcout(\POWERLED.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_11_13_2  (
            .in0(N__29128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30218),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_13_3 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_11_13_3  (
            .in0(N__30371),
            .in1(N__30097),
            .in2(N__30229),
            .in3(N__30288),
            .lcout(),
            .ltout(\VPP_VDDQ.N_64_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_13_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_13_4 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_11_13_4  (
            .in0(N__29127),
            .in1(N__30303),
            .in2(N__29134),
            .in3(N__34855),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_pwrgd_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_13_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_13_5 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_13_5  (
            .in0(N__34856),
            .in1(_gnd_net_),
            .in2(N__29131),
            .in3(N__30319),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34143),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_13_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_13_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNILLP51_1_LC_11_13_6  (
            .in0(N__30273),
            .in1(N__30370),
            .in2(_gnd_net_),
            .in3(N__30214),
            .lcout(\VPP_VDDQ.curr_state_7_0 ),
            .ltout(\VPP_VDDQ.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI2OB42_0_LC_11_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI2OB42_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI2OB42_0_LC_11_13_7 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNI2OB42_0_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__30096),
            .in2(N__30313),
            .in3(N__30274),
            .lcout(\VPP_VDDQ.N_66_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_1 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_11_14_1  (
            .in0(N__30359),
            .in1(N__30095),
            .in2(N__30237),
            .in3(N__30276),
            .lcout(N_246),
            .ltout(N_246_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.G_43_LC_11_14_2 .C_ON=1'b0;
    defparam \POWERLED.G_43_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.G_43_LC_11_14_2 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \POWERLED.G_43_LC_11_14_2  (
            .in0(N__30289),
            .in1(N__30072),
            .in2(N__30292),
            .in3(N__34843),
            .lcout(G_43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNID2IU_0_LC_11_14_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNID2IU_0_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNID2IU_0_LC_11_14_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNID2IU_0_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__30094),
            .in2(_gnd_net_),
            .in3(N__30275),
            .lcout(N_381),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_11_14_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_11_14_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_11_14_7  (
            .in0(N__30358),
            .in1(N__30277),
            .in2(_gnd_net_),
            .in3(N__30233),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34431),
            .ce(N__34714),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_11_15_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_11_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_11_15_0  (
            .in0(N__33081),
            .in1(N__33096),
            .in2(N__33115),
            .in3(N__33657),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_11_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_11_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_11_15_1  (
            .in0(N__30649),
            .in1(N__30643),
            .in2(N__30079),
            .in3(N__30061),
            .lcout(VPP_VDDQ_un6_count),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_11_15_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_11_15_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_11_15_2  (
            .in0(N__33672),
            .in1(N__33144),
            .in2(N__33613),
            .in3(N__33129),
            .lcout(\VPP_VDDQ.un6_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_11_15_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_11_15_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_11_15_3  (
            .in0(N__33627),
            .in1(N__33642),
            .in2(N__33160),
            .in3(N__33594),
            .lcout(\VPP_VDDQ.un6_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_11_15_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_11_15_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_11_15_4  (
            .in0(N__34587),
            .in1(N__34473),
            .in2(N__33565),
            .in3(N__33579),
            .lcout(\VPP_VDDQ.un6_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_11_16_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_11_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__34857),
            .in2(_gnd_net_),
            .in3(N__33703),
            .lcout(\VPP_VDDQ.N_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_12_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_12_3_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32107),
            .lcout(\VPP_VDDQ.N_2192_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_4_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_4_0  (
            .in0(N__30399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30726),
            .lcout(\VPP_VDDQ.N_361_0 ),
            .ltout(\VPP_VDDQ.N_361_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_4_1 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_4_1  (
            .in0(N__30548),
            .in1(_gnd_net_),
            .in2(N__30433),
            .in3(N__31925),
            .lcout(\VPP_VDDQ.N_62 ),
            .ltout(\VPP_VDDQ.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_4_2 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_4_2  (
            .in0(N__30400),
            .in1(N__31971),
            .in2(N__30430),
            .in3(N__30808),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_en ),
            .ltout(\VPP_VDDQ.delayed_vddq_ok_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_3  (
            .in0(N__30328),
            .in1(N__30718),
            .in2(N__30427),
            .in3(N__30402),
            .lcout(VPP_VDDQ_delayed_vddq_ok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4  (
            .in0(N__30401),
            .in1(N__30327),
            .in2(N__30337),
            .in3(N__30717),
            .lcout(\VPP_VDDQ.delayed_vddq_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34222),
            .ce(),
            .sr(N__30703));
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_5 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_5  (
            .in0(N__30817),
            .in1(N__30803),
            .in2(N__30730),
            .in3(N__31926),
            .lcout(\VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30716),
            .lcout(\VPP_VDDQ.N_62_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_5_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_5_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_12_5_0  (
            .in0(N__32090),
            .in1(N__31912),
            .in2(N__31796),
            .in3(N__31342),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_12_5_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJ48C1_14_LC_12_5_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJ48C1_14_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__31324),
            .in2(N__30694),
            .in3(N__31552),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_12_5_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_12_5_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_12_5_2  (
            .in0(N__32088),
            .in1(N__31910),
            .in2(N__30687),
            .in3(N__31746),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_12_5_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIHA461_4_LC_12_5_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIHA461_4_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__30667),
            .in2(N__30691),
            .in3(N__31550),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_4_LC_12_5_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_4_LC_12_5_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_12_5_4  (
            .in0(N__32091),
            .in1(N__31913),
            .in2(N__30688),
            .in3(N__31748),
            .lcout(\VPP_VDDQ.count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34412),
            .ce(N__31633),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_5_LC_12_5_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_5_LC_12_5_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_12_5_5  (
            .in0(N__31914),
            .in1(N__30660),
            .in2(N__32150),
            .in3(N__31770),
            .lcout(\VPP_VDDQ.count_2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34412),
            .ce(N__31633),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_12_5_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_12_5_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_12_5_6  (
            .in0(N__32089),
            .in1(N__31911),
            .in2(N__30661),
            .in3(N__31747),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_12_5_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJD561_5_LC_12_5_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIJD561_5_LC_12_5_7  (
            .in0(N__31306),
            .in1(_gnd_net_),
            .in2(N__31300),
            .in3(N__31551),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_12_6_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_12_6_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_12_6_0  (
            .in0(N__31285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31140),
            .lcout(\PCH_PWRGD.N_174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_LC_12_6_2 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_LC_12_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_LC_12_6_2  (
            .in0(N__31236),
            .in1(N__31210),
            .in2(N__31198),
            .in3(N__31189),
            .lcout(),
            .ltout(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_12_6_3 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_12_6_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_12_6_3  (
            .in0(N__31141),
            .in1(_gnd_net_),
            .in2(N__30961),
            .in3(N__30958),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_12_6_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI38QU_6_LC_12_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI38QU_6_LC_12_6_4  (
            .in0(N__30879),
            .in1(N__30825),
            .in2(_gnd_net_),
            .in3(N__31589),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_12_6_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI38QU_0_6_LC_12_6_5 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \VPP_VDDQ.count_2_RNI38QU_0_6_LC_12_6_5  (
            .in0(N__31590),
            .in1(N__30892),
            .in2(N__30829),
            .in3(N__30880),
            .lcout(),
            .ltout(\VPP_VDDQ.un9_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_12_6_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIOUR33_1_LC_12_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIOUR33_1_LC_12_6_6  (
            .in0(N__31315),
            .in1(N__30868),
            .in2(N__30862),
            .in3(N__30859),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(\VPP_VDDQ.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_6_LC_12_6_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_6_LC_12_6_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_12_6_7  (
            .in0(N__30846),
            .in1(N__32165),
            .in2(N__30832),
            .in3(N__31943),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34350),
            .ce(N__31594),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_12_7_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIFU5C1_12_LC_12_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIFU5C1_12_LC_12_7_0  (
            .in0(N__31372),
            .in1(N__31618),
            .in2(_gnd_net_),
            .in3(N__31465),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_7_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_7_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_12_7_1  (
            .in0(N__32146),
            .in1(N__31941),
            .in2(N__31386),
            .in3(N__31762),
            .lcout(\VPP_VDDQ.count_2_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_12_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIH17C1_13_LC_12_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIH17C1_13_LC_12_7_2  (
            .in0(N__31348),
            .in1(N__31459),
            .in2(_gnd_net_),
            .in3(N__31619),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_15_LC_12_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_15_LC_12_7_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_15_LC_12_7_3  (
            .in0(N__31447),
            .in1(N__31429),
            .in2(N__31417),
            .in3(N__31414),
            .lcout(\VPP_VDDQ.un9_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_12_LC_12_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_12_LC_12_7_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_12_7_5  (
            .in0(N__32147),
            .in1(N__31942),
            .in2(N__31387),
            .in3(N__31764),
            .lcout(\VPP_VDDQ.count_2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34433),
            .ce(N__31622),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_13_LC_12_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_13_LC_12_7_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_12_7_6  (
            .in0(N__31763),
            .in1(N__32149),
            .in2(N__31366),
            .in3(N__31947),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34433),
            .ce(N__31622),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_14_LC_12_7_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_14_LC_12_7_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_12_7_7  (
            .in0(N__32148),
            .in1(N__31338),
            .in2(N__31979),
            .in3(N__31765),
            .lcout(\VPP_VDDQ.count_2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34433),
            .ce(N__31622),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_8_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_8_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_8_0  (
            .in0(N__32151),
            .in1(N__31973),
            .in2(N__32206),
            .in3(N__31779),
            .lcout(\VPP_VDDQ.count_2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_8_1 .LUT_INIT=16'b0001000100000011;
    LogicCell40 \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_8_1  (
            .in0(N__32257),
            .in1(N__32227),
            .in2(N__32194),
            .in3(N__31568),
            .lcout(\VPP_VDDQ.un9_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_8_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_8_2  (
            .in0(N__31567),
            .in1(N__32190),
            .in2(_gnd_net_),
            .in3(N__32256),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_1 ),
            .ltout(\VPP_VDDQ.un1_count_2_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32239),
            .in3(N__32228),
            .lcout(\VPP_VDDQ.count_2_RNIZ0Z_1 ),
            .ltout(\VPP_VDDQ.count_2_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_12_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_1_LC_12_8_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_12_8_4  (
            .in0(N__32152),
            .in1(N__31974),
            .in2(N__32197),
            .in3(N__31781),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34348),
            .ce(N__31569),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_11_LC_12_8_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_11_LC_12_8_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_12_8_5  (
            .in0(N__31780),
            .in1(N__32153),
            .in2(N__32002),
            .in3(N__31975),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34348),
            .ce(N__31569),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_8_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_8_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_8_6  (
            .in0(N__32154),
            .in1(N__32001),
            .in2(N__31989),
            .in3(N__31782),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_8_7 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__31642),
            .in2(N__31636),
            .in3(N__31566),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_12_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__32610),
            .in2(N__33020),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_9_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32635),
            .in3(N__31468),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_9_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33060),
            .in3(N__32338),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_9_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33543),
            .in3(N__32323),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_9_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_12_9_4  (
            .in0(N__33485),
            .in1(_gnd_net_),
            .in2(N__32419),
            .in3(N__32320),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_9_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32544),
            .in3(N__32308),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_9_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_9_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_12_9_6  (
            .in0(N__33486),
            .in1(_gnd_net_),
            .in2(N__32728),
            .in3(N__32290),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_9_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_9_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_12_9_7  (
            .in0(N__33487),
            .in1(N__32842),
            .in2(_gnd_net_),
            .in3(N__32287),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_10_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_12_10_0  (
            .in0(N__33453),
            .in1(_gnd_net_),
            .in2(N__32824),
            .in3(N__32266),
            .lcout(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33043),
            .in3(N__32263),
            .lcout(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_10_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32683),
            .in3(N__32260),
            .lcout(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_10_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_12_10_3  (
            .in0(N__33455),
            .in1(_gnd_net_),
            .in2(N__32752),
            .in3(N__32473),
            .lcout(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_10_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32470),
            .in3(N__32446),
            .lcout(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_12_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_12_10_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32443),
            .in3(N__32425),
            .lcout(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_10_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_12_10_6  (
            .in0(N__32356),
            .in1(N__33456),
            .in2(_gnd_net_),
            .in3(N__32422),
            .lcout(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_12_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_12_LC_12_10_7  (
            .in0(N__32766),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34430),
            .ce(N__33331),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIN6TD_5_LC_12_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIN6TD_5_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIN6TD_5_LC_12_11_0 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \POWERLED.count_clk_RNIN6TD_5_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__32377),
            .in2(N__33292),
            .in3(N__32388),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_12_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_12_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_5_LC_12_11_1  (
            .in0(N__32389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__33333),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_12_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_12_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_15_LC_12_11_2  (
            .in0(N__32365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__33333),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIPD76_15_LC_12_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIPD76_15_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIPD76_15_LC_12_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIPD76_15_LC_12_11_3  (
            .in0(N__33267),
            .in1(N__32371),
            .in2(_gnd_net_),
            .in3(N__32364),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(\POWERLED.count_clkZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_15_LC_12_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_15_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_15_LC_12_11_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.count_clk_RNI_15_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32617),
            .in3(N__32611),
            .lcout(\POWERLED.count_clk_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_12_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_12_11_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.count_clk_1_LC_12_11_5  (
            .in0(N__33471),
            .in1(N__32614),
            .in2(_gnd_net_),
            .in3(N__33018),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__33333),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNITF0E_8_LC_12_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNITF0E_8_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNITF0E_8_LC_12_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNITF0E_8_LC_12_11_6  (
            .in0(N__33257),
            .in1(N__32569),
            .in2(_gnd_net_),
            .in3(N__32580),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_12_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_12_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_8_LC_12_11_7  (
            .in0(N__32581),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34416),
            .ce(N__33333),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_12_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_12_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_clk_10_LC_12_12_0  (
            .in0(N__32557),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33457),
            .lcout(\POWERLED.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34421),
            .ce(N__33316),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8SH6_10_LC_12_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8SH6_10_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8SH6_10_LC_12_12_1 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \POWERLED.count_clk_RNI8SH6_10_LC_12_12_1  (
            .in0(N__32563),
            .in1(N__33454),
            .in2(N__33320),
            .in3(N__32556),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(\POWERLED.count_clkZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_10_LC_12_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_10_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_10_LC_12_12_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.count_clk_RNI_0_10_LC_12_12_2  (
            .in0(N__33067),
            .in1(N__32545),
            .in2(N__32521),
            .in3(N__32679),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_8_LC_12_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_8_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_8_LC_12_12_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_8_LC_12_12_3  (
            .in0(N__32841),
            .in1(N__32518),
            .in2(N__32500),
            .in3(N__33496),
            .lcout(\POWERLED.N_352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_10_LC_12_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_10_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_10_LC_12_12_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \POWERLED.count_clk_RNI_10_LC_12_12_4  (
            .in0(N__33066),
            .in1(N__33039),
            .in2(N__33025),
            .in3(N__33507),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_15_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_10_LC_12_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_10_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_10_LC_12_12_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_1_10_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__32782),
            .in2(N__32980),
            .in3(N__32977),
            .lcout(\POWERLED.un2_count_clk_15_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_8_LC_12_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_8_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_8_LC_12_12_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_8_LC_12_12_7  (
            .in0(N__32840),
            .in1(_gnd_net_),
            .in2(N__32692),
            .in3(N__32821),
            .lcout(\POWERLED.un2_count_clk_15_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJ446_12_LC_12_13_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJ446_12_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJ446_12_LC_12_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_clk_RNIJ446_12_LC_12_13_0  (
            .in0(N__33237),
            .in1(N__32776),
            .in2(_gnd_net_),
            .in3(N__32767),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(\POWERLED.count_clkZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_12_LC_12_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_12_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_12_LC_12_13_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.count_clk_RNI_12_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32740),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_RNIZ0Z_12 ),
            .ltout(\POWERLED.count_clk_RNIZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_11_LC_12_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_11_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_11_LC_12_13_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.count_clk_RNI_11_LC_12_13_2  (
            .in0(N__32631),
            .in1(N__32736),
            .in2(N__32695),
            .in3(N__32678),
            .lcout(\POWERLED.un2_count_clk_15_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIH136_11_LC_12_13_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIH136_11_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIH136_11_LC_12_13_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \POWERLED.count_clk_RNIH136_11_LC_12_13_3  (
            .in0(N__33469),
            .in1(N__33236),
            .in2(N__33343),
            .in3(N__33354),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_12_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_12_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_2_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__32658),
            .in2(_gnd_net_),
            .in3(N__33470),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34450),
            .ce(N__33334),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIHTPD_2_LC_12_13_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIHTPD_2_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIHTPD_2_LC_12_13_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \POWERLED.count_clk_RNIHTPD_2_LC_12_13_5  (
            .in0(N__32659),
            .in1(N__33459),
            .in2(N__32644),
            .in3(N__33235),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(\POWERLED.count_clkZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_2_LC_12_13_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_2_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_2_LC_12_13_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.count_clk_RNI_2_LC_12_13_6  (
            .in0(N__33547),
            .in1(N__33520),
            .in2(N__33514),
            .in3(N__33511),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_12_13_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_12_13_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_11_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__33460),
            .in2(_gnd_net_),
            .in3(N__33355),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34450),
            .ce(N__33334),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_12_14_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_12_14_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_12_14_0  (
            .in0(N__34880),
            .in1(N__33159),
            .in2(N__33175),
            .in3(N__33174),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_1_LC_12_14_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_12_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_12_14_1  (
            .in0(N__34870),
            .in1(N__33145),
            .in2(_gnd_net_),
            .in3(N__33133),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_2_LC_12_14_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_12_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_12_14_2  (
            .in0(N__34881),
            .in1(N__33130),
            .in2(_gnd_net_),
            .in3(N__33118),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_3_LC_12_14_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_12_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_12_14_3  (
            .in0(N__34871),
            .in1(N__33114),
            .in2(_gnd_net_),
            .in3(N__33100),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_4_LC_12_14_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_12_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_12_14_4  (
            .in0(N__34882),
            .in1(N__33097),
            .in2(_gnd_net_),
            .in3(N__33085),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_5_LC_12_14_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_12_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_12_14_5  (
            .in0(N__34872),
            .in1(N__33082),
            .in2(_gnd_net_),
            .in3(N__33070),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_6_LC_12_14_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_12_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_12_14_6  (
            .in0(N__34883),
            .in1(N__33673),
            .in2(_gnd_net_),
            .in3(N__33661),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_7_LC_12_14_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_12_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_12_14_7  (
            .in0(N__34873),
            .in1(N__33658),
            .in2(_gnd_net_),
            .in3(N__33646),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__34462),
            .ce(),
            .sr(N__33704));
    defparam \VPP_VDDQ.count_8_LC_12_15_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_12_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_12_15_0  (
            .in0(N__34887),
            .in1(N__33643),
            .in2(_gnd_net_),
            .in3(N__33631),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.count_9_LC_12_15_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_12_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_12_15_1  (
            .in0(N__34876),
            .in1(N__33628),
            .in2(_gnd_net_),
            .in3(N__33616),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.count_10_LC_12_15_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_12_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_12_15_2  (
            .in0(N__34884),
            .in1(N__33612),
            .in2(_gnd_net_),
            .in3(N__33598),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.count_11_LC_12_15_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_12_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_12_15_3  (
            .in0(N__34874),
            .in1(N__33595),
            .in2(_gnd_net_),
            .in3(N__33583),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.count_12_LC_12_15_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_12_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_12_15_4  (
            .in0(N__34885),
            .in1(N__33580),
            .in2(_gnd_net_),
            .in3(N__33568),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.count_13_LC_12_15_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_12_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_12_15_5  (
            .in0(N__34875),
            .in1(N__33564),
            .in2(_gnd_net_),
            .in3(N__33550),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.count_14_LC_12_15_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_12_15_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_12_15_6  (
            .in0(N__34886),
            .in1(N__34588),
            .in2(_gnd_net_),
            .in3(N__34576),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__34451),
            .ce(),
            .sr(N__33709));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_12_15_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_12_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__34573),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_12_16_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_12_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__34474),
            .in2(_gnd_net_),
            .in3(N__34477),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34461),
            .ce(N__33715),
            .sr(N__33705));
endmodule // TOP
