-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 9 2022 11:23:43

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : out std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__36183\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36181\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36173\ : std_logic;
signal \N__36172\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36163\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36136\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36127\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36100\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36091\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36002\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35965\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35956\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35947\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35939\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35921\ : std_logic;
signal \N__35920\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35911\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35894\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35884\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35876\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35858\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35840\ : std_logic;
signal \N__35839\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35822\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35804\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35785\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35750\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35740\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35723\ : std_logic;
signal \N__35722\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35697\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35687\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35670\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35659\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35634\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35626\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35605\ : std_logic;
signal \N__35602\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35591\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35576\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35557\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35551\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35542\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35512\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35504\ : std_logic;
signal \N__35495\ : std_logic;
signal \N__35492\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35480\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35475\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35472\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35462\ : std_logic;
signal \N__35459\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35446\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35385\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35358\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35346\ : std_logic;
signal \N__35345\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35286\ : std_logic;
signal \N__35279\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35256\ : std_logic;
signal \N__35249\ : std_logic;
signal \N__35240\ : std_logic;
signal \N__35237\ : std_logic;
signal \N__35232\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35183\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35153\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35126\ : std_logic;
signal \N__35123\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35111\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35097\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35049\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34969\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34960\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34941\ : std_logic;
signal \N__34938\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34925\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34886\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34880\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34830\ : std_logic;
signal \N__34821\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34811\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34808\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34754\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34715\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34708\ : std_logic;
signal \N__34705\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34700\ : std_logic;
signal \N__34699\ : std_logic;
signal \N__34696\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34690\ : std_logic;
signal \N__34687\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34685\ : std_logic;
signal \N__34682\ : std_logic;
signal \N__34681\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34678\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34676\ : std_logic;
signal \N__34673\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34664\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34660\ : std_logic;
signal \N__34657\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34652\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34622\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34616\ : std_logic;
signal \N__34613\ : std_logic;
signal \N__34610\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34601\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34592\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34586\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34583\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34577\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34550\ : std_logic;
signal \N__34547\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34522\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34514\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34496\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34483\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34475\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34469\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34460\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34451\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34405\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34315\ : std_logic;
signal \N__34312\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34297\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34287\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34222\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34199\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34160\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34064\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34061\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34033\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33992\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33974\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33958\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33907\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33899\ : std_logic;
signal \N__33896\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33873\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33824\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33794\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33773\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33740\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33728\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33713\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33667\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33663\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33660\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33652\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33602\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33590\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33446\ : std_logic;
signal \N__33443\ : std_logic;
signal \N__33440\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33434\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33404\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33386\ : std_logic;
signal \N__33377\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33371\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33368\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33308\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33302\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33253\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33218\ : std_logic;
signal \N__33215\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33182\ : std_logic;
signal \N__33179\ : std_logic;
signal \N__33176\ : std_logic;
signal \N__33173\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33160\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33146\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33125\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33101\ : std_logic;
signal \N__33098\ : std_logic;
signal \N__33095\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33073\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33065\ : std_logic;
signal \N__33062\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33056\ : std_logic;
signal \N__33053\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33035\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33002\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32985\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32960\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32926\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32891\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32882\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32853\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32849\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32845\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32823\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32813\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32780\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32769\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32742\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32710\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32690\ : std_logic;
signal \N__32687\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32676\ : std_logic;
signal \N__32675\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32655\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32649\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32598\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32525\ : std_logic;
signal \N__32524\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32484\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32480\ : std_logic;
signal \N__32477\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32434\ : std_logic;
signal \N__32431\ : std_logic;
signal \N__32428\ : std_logic;
signal \N__32425\ : std_logic;
signal \N__32420\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32408\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32402\ : std_logic;
signal \N__32399\ : std_logic;
signal \N__32396\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32378\ : std_logic;
signal \N__32377\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32375\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32356\ : std_logic;
signal \N__32353\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32309\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32270\ : std_logic;
signal \N__32267\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32251\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32237\ : std_logic;
signal \N__32234\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32192\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32153\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32063\ : std_logic;
signal \N__32062\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32041\ : std_logic;
signal \N__32030\ : std_logic;
signal \N__32027\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32018\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32014\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31991\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31967\ : std_logic;
signal \N__31964\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31955\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31916\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31903\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31868\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31864\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31826\ : std_logic;
signal \N__31825\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31822\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31814\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31807\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31799\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31778\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31676\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31646\ : std_logic;
signal \N__31643\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31631\ : std_logic;
signal \N__31628\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31601\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31574\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31550\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31508\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31486\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31421\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31412\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31409\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31406\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31403\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31400\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31334\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31319\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31295\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31276\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31253\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31242\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31144\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31112\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31107\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31046\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31025\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31019\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31016\ : std_logic;
signal \N__31011\ : std_logic;
signal \N__31008\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__30998\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30955\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30914\ : std_logic;
signal \N__30911\ : std_logic;
signal \N__30908\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30900\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30809\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30799\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30779\ : std_logic;
signal \N__30776\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30746\ : std_logic;
signal \N__30743\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30716\ : std_logic;
signal \N__30713\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30704\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30658\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30641\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30602\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30586\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30578\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30575\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30544\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30539\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30526\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30520\ : std_logic;
signal \N__30517\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30503\ : std_logic;
signal \N__30500\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30467\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30440\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30434\ : std_logic;
signal \N__30431\ : std_logic;
signal \N__30428\ : std_logic;
signal \N__30425\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30401\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30364\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30310\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30304\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30290\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30257\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30201\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30196\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30191\ : std_logic;
signal \N__30188\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30135\ : std_logic;
signal \N__30132\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30107\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30059\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30044\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30016\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29960\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29925\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29919\ : std_logic;
signal \N__29916\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29894\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29853\ : std_logic;
signal \N__29850\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29777\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29735\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29729\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29720\ : std_logic;
signal \N__29717\ : std_logic;
signal \N__29714\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29704\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29698\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29630\ : std_logic;
signal \N__29627\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29600\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29563\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29461\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29452\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29443\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29423\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29413\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29403\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29386\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29370\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29352\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29309\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29188\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29182\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29160\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28961\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28854\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28700\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28675\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28619\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28603\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28568\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28535\ : std_logic;
signal \N__28532\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28526\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28511\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28496\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28490\ : std_logic;
signal \N__28487\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28463\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28409\ : std_logic;
signal \N__28406\ : std_logic;
signal \N__28403\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28349\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28316\ : std_logic;
signal \N__28313\ : std_logic;
signal \N__28310\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28304\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28274\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28271\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28262\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28241\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28214\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28184\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28179\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28094\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__27998\ : std_logic;
signal \N__27995\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27944\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27868\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27846\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27731\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27677\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27593\ : std_logic;
signal \N__27590\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27518\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27491\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27473\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27467\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27422\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27416\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27329\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27317\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27266\ : std_logic;
signal \N__27263\ : std_logic;
signal \N__27260\ : std_logic;
signal \N__27257\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27206\ : std_logic;
signal \N__27203\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27170\ : std_logic;
signal \N__27167\ : std_logic;
signal \N__27164\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27155\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27122\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27113\ : std_logic;
signal \N__27110\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27095\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27086\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27071\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27043\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27017\ : std_logic;
signal \N__27014\ : std_logic;
signal \N__27011\ : std_logic;
signal \N__27008\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26945\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26921\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26907\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26901\ : std_logic;
signal \N__26898\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26849\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26821\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26783\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26749\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26729\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26711\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26707\ : std_logic;
signal \N__26704\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26696\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26543\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26453\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26407\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25724\ : std_logic;
signal \N__25721\ : std_logic;
signal \N__25718\ : std_logic;
signal \N__25715\ : std_logic;
signal \N__25712\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25709\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25631\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25592\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25562\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25538\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25529\ : std_logic;
signal \N__25526\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25406\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25281\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25195\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25052\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25040\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25016\ : std_logic;
signal \N__25013\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24701\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24668\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24656\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24617\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24599\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24380\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24244\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23873\ : std_logic;
signal \N__23870\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23399\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23006\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22910\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22772\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22715\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22628\ : std_logic;
signal \N__22625\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22142\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22133\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21758\ : std_logic;
signal \N__21755\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21216\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20885\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20747\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20720\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20447\ : std_logic;
signal \N__20444\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20390\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20330\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20126\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20117\ : std_logic;
signal \N__20114\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20105\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20048\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20027\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19949\ : std_logic;
signal \N__19940\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19934\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19442\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18978\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18923\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18589\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18583\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18539\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18362\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17534\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17309\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17246\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16892\ : std_logic;
signal \N__16889\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16799\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16571\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16565\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16265\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15747\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14912\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14495\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \VCCG0\ : std_logic;
signal \N_428_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.m14_i_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \HDA_STRAP.N_16_cascade_\ : std_logic;
signal \HDA_STRAP.HDA_SDO_ATP_3_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal \HDA_STRAP.un4_count_9_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_12\ : std_logic;
signal \HDA_STRAP.un4_count_11\ : std_logic;
signal \HDA_STRAP.un4_count_13_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_10\ : std_logic;
signal \HDA_STRAP.un4_count_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_5\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_4_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_10\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_13\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_1\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \POWERLED.g1_i_a4_0_1_cascade_\ : std_logic;
signal \POWERLED.N_12\ : std_logic;
signal \POWERLED.N_5_cascade_\ : std_logic;
signal \POWERLED.pwm_out_en_cascade_\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.N_11\ : std_logic;
signal \POWERLED.g0_2_1\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal \POWERLED.N_2360_i_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_11_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_9\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_8\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \bfn_2_1_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_1\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_3\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7\ : std_logic;
signal \HDA_STRAP.countZ0Z_8\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_9\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_13\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_15\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \HDA_STRAP.curr_state_RNIH91AZ0Z_0\ : std_logic;
signal \HDA_STRAP.un4_count\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_16\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_rst_7\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_7\ : std_logic;
signal \PCH_PWRGD.count_rst_3\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_4_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_5_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_3_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_6_0\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2226_i_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_state_7_0\ : std_logic;
signal \PCH_PWRGD.N_386_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_1_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_2_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_11_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_11_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_12_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_2\ : std_logic;
signal \PCH_PWRGD.count_rst_14\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_0_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_10\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.curr_state_0_0\ : std_logic;
signal \PCH_PWRGD.N_2244_i\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.N_2244_i_cascade_\ : std_logic;
signal \PCH_PWRGD.N_655_cascade_\ : std_logic;
signal \PCH_PWRGD.m6_i_i_a2\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.N_386\ : std_logic;
signal \PCH_PWRGD.N_2226_i\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.N_655\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \N_626_cascade_\ : std_logic;
signal \POWERLED.G_30Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ_un6_count\ : std_logic;
signal \G_30_cascade_\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_4_l_fx\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.count_1_5_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.count_1_5\ : std_logic;
signal \POWERLED.un79_clk_100khzlto6_0_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khz\ : std_logic;
signal \POWERLED.un79_clk_100khz_cascade_\ : std_logic;
signal \POWERLED.N_2360_i\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \VPP_VDDQ.N_64_i\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \bfn_2_14_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.N_92_0\ : std_logic;
signal \G_30\ : std_logic;
signal \VPP_VDDQ.count_2_1_8_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.count_2_1_9_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.count_2_1_14_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_4_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_4\ : std_logic;
signal \VPP_VDDQ.count_2_0_5\ : std_logic;
signal \VPP_VDDQ.count_2_1_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_12_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \VPP_VDDQ_curr_state_0\ : std_logic;
signal \VPP_VDDQ_curr_state_1\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\ : std_logic;
signal \N_626\ : std_logic;
signal \PCH_PWRGD.curr_state_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.N_38_f0\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \VPP_VDDQ.count_2_0_10\ : std_logic;
signal \VPP_VDDQ.count_2_1_10_cascade_\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_4_7_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \POWERLED.N_4842_i\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.count_i_3\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \POWERLED.count_RNIGTVS_1Z0Z_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.count_i_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.N_4841_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.count_i_8\ : std_logic;
signal \bfn_4_10_0_\ : std_logic;
signal \POWERLED.N_4849_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.count_i_10\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.count_i_11\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.N_4851_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.N_4855_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.N_4856_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.N_437_cascade_\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.curr_state_1_0\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_8\ : std_logic;
signal \POWERLED.count_RNIAKSS_0Z0Z_2\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.un79_clk_100khzlto4_0_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlt6\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_8\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.count_RNIJEFE_0Z0Z_4\ : std_logic;
signal \POWERLED.mult1_un159_sum_i_8\ : std_logic;
signal \POWERLED.count_RNIUGSJ_0Z0Z_1\ : std_logic;
signal \POWERLED.N_660\ : std_logic;
signal \POWERLED.count_0_sqmuxa_cascade_\ : std_logic;
signal \POWERLED.count_1_0_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_1_1\ : std_logic;
signal \POWERLED.count_1_1_cascade_\ : std_logic;
signal \POWERLED.un1_count_axb_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.countZ0Z_14_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5\ : std_logic;
signal \POWERLED.g1_i_o4_4\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \VPP_VDDQ.count_2_0_2\ : std_logic;
signal \VPP_VDDQ.count_2_1_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\ : std_logic;
signal \VPP_VDDQ.count_2_1_13\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \PCH_PWRGD.N_670\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal vccst_en : std_logic;
signal \G_12\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_8\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.un1_count_axb_1\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \POWERLED.un1_count_axb_2\ : std_logic;
signal \POWERLED.count_1_2\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_cry_2_c_RNICZ0Z419\ : std_logic;
signal \POWERLED.un1_count_cry_2\ : std_logic;
signal \POWERLED.un1_count_axb_4\ : std_logic;
signal \POWERLED.count_1_4\ : std_logic;
signal \POWERLED.un1_count_cry_3\ : std_logic;
signal \POWERLED.un1_count_axb_5\ : std_logic;
signal \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\ : std_logic;
signal \POWERLED.un1_count_cry_4\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.count_1_11\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.un1_count_cry_11\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.count_1_14\ : std_logic;
signal \POWERLED.un1_count_cry_13\ : std_logic;
signal \POWERLED.count_0_sqmuxa\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\ : std_logic;
signal \POWERLED.un1_count_axb_12\ : std_logic;
signal \POWERLED.count_1_9\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.count_1_10\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.count_1_6\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \POWERLED.count_1_8\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.count_2_1_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_ok_cascade_\ : std_logic;
signal vccst_pwrgd : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_9\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_0_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\ : std_logic;
signal \VPP_VDDQ.N_1_i_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_6_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_6\ : std_logic;
signal v1p8a_ok : std_logic;
signal v5a_ok : std_logic;
signal v33a_ok : std_logic;
signal slp_susn : std_logic;
signal v33a_enn : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_1_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2_1_11_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.N_60_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.N_60\ : std_logic;
signal \VPP_VDDQ.N_60_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \G_2161\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un166_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_8\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_8\ : std_logic;
signal \POWERLED.count_RNICOIT_0Z0Z_12\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \POWERLED.count_1_13\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.countZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.count_1_12\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_3_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_6\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_3\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.g1_i_o4_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.count_1_7\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.N_6\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \bfn_6_15_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \VPP_VDDQ.N_53_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.N_664_cascade_\ : std_logic;
signal \VPP_VDDQ.m4_0_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIZ0Z_1\ : std_logic;
signal vddq_ok : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_664\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.N_53\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal \N_557_g\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12_cascade_\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_cascade_\ : std_logic;
signal \POWERLED.dutycycle_1_0_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_0_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_1_cascade_\ : std_logic;
signal \dutycycle_RNII6848_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_1\ : std_logic;
signal \POWERLED.dutycycle_eena_0_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.N_15\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_\ : std_logic;
signal \POWERLED.N_672_cascade_\ : std_logic;
signal \dutycycle_RNI_1_5\ : std_logic;
signal \POWERLED_un1_dutycycle_172_m1\ : std_logic;
signal \dutycycle_RNI_3_1_cascade_\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_4_1\ : std_logic;
signal \POWERLED.g0_7_a2_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_0\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0_a2_0_4_cascade_\ : std_logic;
signal \POWERLED.N_604\ : std_logic;
signal \POWERLED.func_state_RNI1O2V5Z0Z_1\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.N_9_i_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_32_and_i_0_a2_0_0_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0_a2_0_3\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_0\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_0\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_2\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_2\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_3\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_11\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_12\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_28\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_axb_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \POWERLED.N_413_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.N_413_N\ : std_logic;
signal \POWERLED.N_430_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_1\ : std_logic;
signal \SUSWARN_N_fast\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m0\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m1_ns_1_cascade_\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m1\ : std_logic;
signal \COUNTER.tmp_0_fast_RNI0RLUZ0Z1\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_10Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.N_676_cascade_\ : std_logic;
signal \G_11_i_a10_0_1_cascade_\ : std_logic;
signal \G_11_i_2\ : std_logic;
signal \N_9_2_cascade_\ : std_logic;
signal \N_8_3\ : std_logic;
signal \G_11_i_a10_0_1\ : std_logic;
signal \N_8_3_cascade_\ : std_logic;
signal \POWERLED.N_10_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_1\ : std_logic;
signal \POWERLED.dutycycle_0_5\ : std_logic;
signal \POWERLED.g0_i_o4_2\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5_cascade_\ : std_logic;
signal \POWERLED.N_546\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_5\ : std_logic;
signal \POWERLED.N_612\ : std_logic;
signal \N_16_0\ : std_logic;
signal \POWERLED.g0_0_1\ : std_logic;
signal \POWERLED.N_598_cascade_\ : std_logic;
signal \POWERLED.N_450_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI5FJ65Z0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI5FJ65Z0Z_13_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11_cascade_\ : std_logic;
signal \POWERLED.N_2336_i\ : std_logic;
signal \POWERLED.N_449\ : std_logic;
signal \POWERLED.un1_m2_e_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_56_a1_2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNIT70K5Z0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_8_cascade_\ : std_logic;
signal \POWERLED.N_6_3_cascade_\ : std_logic;
signal \POWERLED.g0_9_1_0\ : std_logic;
signal \POWERLED.N_9_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_15Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.N_4_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_12_1_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ1Z_14\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_15\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.N_492\ : std_logic;
signal \POWERLED.count_clk_en_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \bfn_8_16_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_axb_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11\ : std_logic;
signal \POWERLED.count_clk_1_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12_cZ0\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.count_clk_1_15\ : std_logic;
signal \POWERLED.un1_count_clk_2_axb_14\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11\ : std_logic;
signal \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_264_i\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.N_662\ : std_logic;
signal \RSMRST_PWRGD.N_555_cascade_\ : std_logic;
signal \RSMRST_PWRGD.G_14\ : std_logic;
signal \N_92_g\ : std_logic;
signal \RSMRST_PWRGD.G_14_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_92_1\ : std_logic;
signal \POWERLED.N_423_0_cascade_\ : std_logic;
signal \POWERLED.g1_cascade_\ : std_logic;
signal \POWERLED.g0_0_0\ : std_logic;
signal \POWERLED.N_8_0_0\ : std_logic;
signal \POWERLED.g0_0_2_cascade_\ : std_logic;
signal \POWERLED.N_541_cascade_\ : std_logic;
signal \POWERLED.N_542\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \POWERLED.g2\ : std_logic;
signal \POWERLED.g0_0_5\ : std_logic;
signal \POWERLED.g2_0\ : std_logic;
signal \POWERLED.g2_cascade_\ : std_logic;
signal \POWERLED.N_13_0_0_0\ : std_logic;
signal \POWERLED.func_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_0\ : std_logic;
signal suswarn_n : std_logic;
signal \POWERLED.N_8_0_cascade_\ : std_logic;
signal \POWERLED.N_16_2\ : std_logic;
signal \POWERLED.dutycycle_e_N_3L4_0_1_cascade_\ : std_logic;
signal \POWERLED.g0_8Z0Z_0\ : std_logic;
signal \POWERLED.N_435_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_0\ : std_logic;
signal \POWERLED.func_state_1_m2s2_i_0_0\ : std_logic;
signal \POWERLED.N_423_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_10Z0Z_0\ : std_logic;
signal \POWERLED.N_613\ : std_logic;
signal \POWERLED.un1_clk_100khz_51_and_i_3_1_cascade_\ : std_logic;
signal \POWERLED.N_252_N\ : std_logic;
signal \POWERLED.dutycycle_eena_13_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_13_cascade_\ : std_logic;
signal \POWERLED.N_452\ : std_logic;
signal \POWERLED.dutycycle_set_1\ : std_logic;
signal \POWERLED.func_state_RNI12ASZ0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI12ASZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3\ : std_logic;
signal \POWERLED.dutycycle_eena_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_13Z0Z_0\ : std_logic;
signal \POWERLED.N_2363_0_cascade_\ : std_logic;
signal \POWERLED.N_12_3_0\ : std_logic;
signal \G_11_i_a10_2_1_cascade_\ : std_logic;
signal \POWERLED.g2_3\ : std_logic;
signal \N_28\ : std_logic;
signal \N_7\ : std_logic;
signal \N_50\ : std_logic;
signal \N_7_cascade_\ : std_logic;
signal \POWERLED.N_2363_0\ : std_logic;
signal \POWERLED.g1_0_1_cascade_\ : std_logic;
signal \N_43\ : std_logic;
signal \POWERLED.g2_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_7_l_fx\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \N_428\ : std_logic;
signal pch_pwrok : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \dutycycle_RNII6848_0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_cZ0\ : std_logic;
signal \POWERLED.N_435_i\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_53_59_a0_0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_56_a1_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_0\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.G_7_i_a5_1_1_cascade_\ : std_logic;
signal \POWERLED.N_11_1\ : std_logic;
signal \POWERLED.N_16_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.g0_9_1\ : std_logic;
signal \POWERLED.g0_9_1_1_0\ : std_logic;
signal \POWERLED.dutycycle_RNIHDMC5Z0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI6SKJ1Z0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNIHDMC5Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_41_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\ : std_logic;
signal \POWERLED.dutycycle_RNIHDMC5Z0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.N_17_cascade_\ : std_logic;
signal \POWERLED.N_8_2\ : std_logic;
signal \POWERLED.G_7_i_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.N_625\ : std_logic;
signal \POWERLED.N_625_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNINSEUC_0Z0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.count_clk_1_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_0\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_2_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNINSEUCZ0Z_10\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_o2_1_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.count_clk_1_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_axb_12\ : std_logic;
signal \POWERLED.count_clk_1_14\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.count_off_0_9\ : std_logic;
signal \POWERLED.count_offZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_off_1_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.count_off_1_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.N_627\ : std_logic;
signal \POWERLED.N_688\ : std_logic;
signal \POWERLED.N_74\ : std_logic;
signal \POWERLED.N_6_1_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_1_cascade_\ : std_logic;
signal \POWERLED.func_state_cascade_\ : std_logic;
signal \POWERLED.N_426_i\ : std_logic;
signal \POWERLED.N_562\ : std_logic;
signal \POWERLED.func_state_enZ0\ : std_logic;
signal \POWERLED.func_state_1_m2_1\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\ : std_logic;
signal \POWERLED.count_off_0_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_offZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.un34_clk_100khz_11\ : std_logic;
signal \POWERLED.un34_clk_100khz_8_cascade_\ : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10_cascade_\ : std_logic;
signal \POWERLED.count_off_RNI8AQHZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m2_ns_1_1\ : std_logic;
signal \POWERLED.N_494\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_i_m2_1_6_cascade_\ : std_logic;
signal \POWERLED.N_453\ : std_logic;
signal \POWERLED.N_133\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0\ : std_logic;
signal \POWERLED.N_490\ : std_logic;
signal \POWERLED.g1_0_2\ : std_logic;
signal \POWERLED.func_state_RNI2MQDZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_13_1_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_a2_d\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\ : std_logic;
signal \POWERLED.dutycycle_e_1_4\ : std_logic;
signal \POWERLED.dutycycle_e_1_4_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIJ17U4Z0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\ : std_logic;
signal \POWERLED.dutycycle_e_1_7\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.dutycycle_e_1_7_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI9S7D5Z0Z_1\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_25_0_tz_1_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_4\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI2MQDZ0Z_1\ : std_logic;
signal \POWERLED.func_state_RNI2MQDZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI_8Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.func_state_RNIMQ0F_0Z0Z_1\ : std_logic;
signal \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d\ : std_logic;
signal \POWERLED.func_state_RNIMQ0F_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI2MQDZ0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNIEBSB1Z0Z_7\ : std_logic;
signal \POWERLED.N_545\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\ : std_logic;
signal \POWERLED.N_71\ : std_logic;
signal \POWERLED.N_2075_tz_tz\ : std_logic;
signal \POWERLED.N_600\ : std_logic;
signal \POWERLED.count_clk_en_0\ : std_logic;
signal \POWERLED.N_443\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_1\ : std_logic;
signal \POWERLED.N_443_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNINSEUCZ0Z_7\ : std_logic;
signal \POWERLED.N_668\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_2\ : std_logic;
signal \N_247\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_0\ : std_logic;
signal \RSMRSTn_rep1\ : std_logic;
signal \POWERLED.N_506_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_10\ : std_logic;
signal \POWERLED.g0_i_0_1\ : std_logic;
signal \POWERLED.N_514_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIHDMC5Z0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.N_508\ : std_logic;
signal \POWERLED.N_512_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_11\ : std_logic;
signal \POWERLED.N_526_cascade_\ : std_logic;
signal \POWERLED.un1_clk_100khz_47_and_i_1\ : std_logic;
signal \POWERLED.dutycycle_en_11\ : std_logic;
signal \POWERLED.N_518_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNIE3861_0Z0Z_12\ : std_logic;
signal \POWERLED.N_520_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIPK9V4Z0Z_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNIN405GZ0\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \POWERLED.count_off_RNI8AQHZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_0_0_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.count_off_1_14\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.count_off_0_7\ : std_logic;
signal \POWERLED.count_off_1_8\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.count_off_0_2\ : std_logic;
signal \POWERLED.count_off_1_5\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_0_6\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_offZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_9\ : std_logic;
signal \POWERLED.count_off_0_11\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_off_1_13\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_offZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.un34_clk_100khz_10\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \POWERLED.count_off_1_0_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_offZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1\ : std_logic;
signal \POWERLED.N_123\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_a6_1_0_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_4\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_0_2_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_5_cascade_\ : std_logic;
signal \POWERLED.N_421\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_0_2_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI31IBHZ0Z_0\ : std_logic;
signal \POWERLED.N_6_2\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.func_state_RNIBVNSZ0Z_0\ : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.func_state_RNI_3Z0Z_1\ : std_logic;
signal \POWERLED.func_state_RNIBVNSZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m0_1_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_7_2\ : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal v5s_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_1_cascade_\ : std_logic;
signal v33s_ok : std_logic;
signal vccin_en : std_logic;
signal \POWERLED.N_253\ : std_logic;
signal \POWERLED.func_state_RNI_6Z0Z_1\ : std_logic;
signal \POWERLED.g1_1\ : std_logic;
signal \POWERLED.func_state_RNI_6Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_2361_0_cascade_\ : std_logic;
signal \N_6_0\ : std_logic;
signal \POWERLED.dutycycle_e_N_6L11_1\ : std_logic;
signal \POWERLED.dutycycle_RNI2MQDZ0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIOGRSZ0Z_4\ : std_logic;
signal \POWERLED.G_11_i_o10_1_0\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \N_9_0\ : std_logic;
signal \RSMRSTn_rep2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.N_488\ : std_logic;
signal \POWERLED.N_540_1\ : std_logic;
signal \POWERLED_un1_dutycycle_172_m0_0\ : std_logic;
signal \POWERLED.N_435\ : std_logic;
signal \POWERLED.func_state_RNI_4Z0Z_1\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m0_ns_1_0\ : std_logic;
signal \POWERLED.func_state_RNI_4Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI5DLRZ0Z_5\ : std_logic;
signal \SUSWARN_N_rep1\ : std_logic;
signal \POWERLED.dutycycle_RNI7ABC3Z0Z_5_cascade_\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \POWERLED.g2_1_1\ : std_logic;
signal \POWERLED.g1_1cf0\ : std_logic;
signal \POWERLED.dutycycleZ1Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \POWERLED.un1_clk_100khz_32_and_i_0cf0_cascade_\ : std_logic;
signal \RSMRSTn_fast\ : std_logic;
signal \POWERLED.un1_clk_100khz_32_and_i_0\ : std_logic;
signal v5s_enn : std_logic;
signal \POWERLED.N_2291_i\ : std_logic;
signal \POWERLED.N_676\ : std_logic;
signal \POWERLED.dutycycle_RNI6SKJ1Z0Z_3\ : std_logic;
signal \POWERLED.func_state_RNILP0FZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_523\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIHDMC5Z0Z_3\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\ : std_logic;
signal \POWERLED.dutycycleZ1Z_3\ : std_logic;
signal \POWERLED.N_430_iZ0\ : std_logic;
signal \POWERLED.N_5_0_cascade_\ : std_logic;
signal \POWERLED.N_12_2\ : std_logic;
signal \POWERLED.g0_7_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.i2_mux\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.N_2341_i_cascade_\ : std_logic;
signal \POWERLED.N_430\ : std_logic;
signal \POWERLED.N_529_cascade_\ : std_logic;
signal \G_141\ : std_logic;
signal \POWERLED.dutycycle_en_12\ : std_logic;
signal \POWERLED.func_state_RNILP0FZ0Z_1\ : std_logic;
signal \POWERLED.func_state\ : std_logic;
signal \POWERLED.N_527\ : std_logic;
signal \POWERLED.N_2341_i\ : std_logic;
signal \POWERLED.un1_clk_100khz_48_and_i_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_8\ : std_logic;
signal \POWERLED.g0_i_0_0_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal vpp_en : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.G_7_i_o5_0\ : std_logic;
signal slp_s4n : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_e_N_3L4_1\ : std_logic;
signal \POWERLED.func_state_RNI_8Z0Z_1\ : std_logic;
signal \VCCST_EN_i_1\ : std_logic;
signal \POWERLED.N_203\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.N_505\ : std_logic;
signal \count_clk_RNINSEUC_0_6\ : std_logic;
signal \POWERLED.N_412_i\ : std_logic;
signal slp_s3n : std_logic;
signal \POWERLED.N_251\ : std_logic;
signal rsmrstn : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.N_524\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.func_state_RNIUQMRH_0_1\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal fpga_osc : std_logic;
signal \POWERLED.count_clk_en\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    SLP_S0n <= \SLP_S0n_wire\;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__36183\,
            DIN => \N__36182\,
            DOUT => \N__36181\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36183\,
            PADOUT => \N__36182\,
            PADIN => \N__36181\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36174\,
            DIN => \N__36173\,
            DOUT => \N__36172\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36174\,
            PADOUT => \N__36173\,
            PADIN => \N__36172\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19646\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36165\,
            DIN => \N__36164\,
            DOUT => \N__36163\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36165\,
            PADOUT => \N__36164\,
            PADIN => \N__36163\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19710\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36156\,
            DIN => \N__36155\,
            DOUT => \N__36154\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36156\,
            PADOUT => \N__36155\,
            PADIN => \N__36154\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14906\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36147\,
            DIN => \N__36146\,
            DOUT => \N__36145\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36147\,
            PADOUT => \N__36146\,
            PADIN => \N__36145\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36138\,
            DIN => \N__36137\,
            DOUT => \N__36136\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36138\,
            PADOUT => \N__36137\,
            PADIN => \N__36136\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36129\,
            DIN => \N__36128\,
            DOUT => \N__36127\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36129\,
            PADOUT => \N__36128\,
            PADIN => \N__36127\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36120\,
            DIN => \N__36119\,
            DOUT => \N__36118\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36120\,
            PADOUT => \N__36119\,
            PADIN => \N__36118\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36111\,
            DIN => \N__36110\,
            DOUT => \N__36109\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36111\,
            PADOUT => \N__36110\,
            PADIN => \N__36109\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30817\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__36102\,
            DIN => \N__36101\,
            DOUT => \N__36100\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36102\,
            PADOUT => \N__36101\,
            PADIN => \N__36100\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36093\,
            DIN => \N__36092\,
            DOUT => \N__36091\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36093\,
            PADOUT => \N__36092\,
            PADIN => \N__36091\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36084\,
            DIN => \N__36083\,
            DOUT => \N__36082\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36084\,
            PADOUT => \N__36083\,
            PADIN => \N__36082\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14630\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36075\,
            DIN => \N__36074\,
            DOUT => \N__36073\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36075\,
            PADOUT => \N__36074\,
            PADIN => \N__36073\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36066\,
            DIN => \N__36065\,
            DOUT => \N__36064\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36066\,
            PADOUT => \N__36065\,
            PADIN => \N__36064\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__36057\,
            DIN => \N__36056\,
            DOUT => \N__36055\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36057\,
            PADOUT => \N__36056\,
            PADIN => \N__36055\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36048\,
            DIN => \N__36047\,
            DOUT => \N__36046\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36048\,
            PADOUT => \N__36047\,
            PADIN => \N__36046\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36039\,
            DIN => \N__36038\,
            DOUT => \N__36037\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36039\,
            PADOUT => \N__36038\,
            PADIN => \N__36037\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__18557\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__36030\,
            DIN => \N__36029\,
            DOUT => \N__36028\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36030\,
            PADOUT => \N__36029\,
            PADIN => \N__36028\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36021\,
            DIN => \N__36020\,
            DOUT => \N__36019\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36021\,
            PADOUT => \N__36020\,
            PADIN => \N__36019\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36012\,
            DIN => \N__36011\,
            DOUT => \N__36010\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36012\,
            PADOUT => \N__36011\,
            PADIN => \N__36010\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24697\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36003\,
            DIN => \N__36002\,
            DOUT => \N__36001\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__36003\,
            PADOUT => \N__36002\,
            PADIN => \N__36001\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35994\,
            DIN => \N__35993\,
            DOUT => \N__35992\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35994\,
            PADOUT => \N__35993\,
            PADIN => \N__35992\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35985\,
            DIN => \N__35984\,
            DOUT => \N__35983\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35985\,
            PADOUT => \N__35984\,
            PADIN => \N__35983\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35976\,
            DIN => \N__35975\,
            DOUT => \N__35974\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35976\,
            PADOUT => \N__35975\,
            PADIN => \N__35974\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35967\,
            DIN => \N__35966\,
            DOUT => \N__35965\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35967\,
            PADOUT => \N__35966\,
            PADIN => \N__35965\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__35152\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35958\,
            DIN => \N__35957\,
            DOUT => \N__35956\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35958\,
            PADOUT => \N__35957\,
            PADIN => \N__35956\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35949\,
            DIN => \N__35948\,
            DOUT => \N__35947\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35949\,
            PADOUT => \N__35948\,
            PADIN => \N__35947\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19532\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35940\,
            DIN => \N__35939\,
            DOUT => \N__35938\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35940\,
            PADOUT => \N__35939\,
            PADIN => \N__35938\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25084\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35931\,
            DIN => \N__35930\,
            DOUT => \N__35929\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35931\,
            PADOUT => \N__35930\,
            PADIN => \N__35929\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35922\,
            DIN => \N__35921\,
            DOUT => \N__35920\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35922\,
            PADOUT => \N__35921\,
            PADIN => \N__35920\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35913\,
            DIN => \N__35912\,
            DOUT => \N__35911\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35913\,
            PADOUT => \N__35912\,
            PADIN => \N__35911\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35904\,
            DIN => \N__35903\,
            DOUT => \N__35902\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35904\,
            PADOUT => \N__35903\,
            PADIN => \N__35902\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35895\,
            DIN => \N__35894\,
            DOUT => \N__35893\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35895\,
            PADOUT => \N__35894\,
            PADIN => \N__35893\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35886\,
            DIN => \N__35885\,
            DOUT => \N__35884\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35886\,
            PADOUT => \N__35885\,
            PADIN => \N__35884\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14039\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35877\,
            DIN => \N__35876\,
            DOUT => \N__35875\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35877\,
            PADOUT => \N__35876\,
            PADIN => \N__35875\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35868\,
            DIN => \N__35867\,
            DOUT => \N__35866\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35868\,
            PADOUT => \N__35867\,
            PADIN => \N__35866\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32867\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35859\,
            DIN => \N__35858\,
            DOUT => \N__35857\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35859\,
            PADOUT => \N__35858\,
            PADIN => \N__35857\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35850\,
            DIN => \N__35849\,
            DOUT => \N__35848\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35850\,
            PADOUT => \N__35849\,
            PADIN => \N__35848\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35841\,
            DIN => \N__35840\,
            DOUT => \N__35839\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35841\,
            PADOUT => \N__35840\,
            PADIN => \N__35839\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35832\,
            DIN => \N__35831\,
            DOUT => \N__35830\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35832\,
            PADOUT => \N__35831\,
            PADIN => \N__35830\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35823\,
            DIN => \N__35822\,
            DOUT => \N__35821\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35823\,
            PADOUT => \N__35822\,
            PADIN => \N__35821\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19769\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35814\,
            DIN => \N__35813\,
            DOUT => \N__35812\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35814\,
            PADOUT => \N__35813\,
            PADIN => \N__35812\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35805\,
            DIN => \N__35804\,
            DOUT => \N__35803\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35805\,
            PADOUT => \N__35804\,
            PADIN => \N__35803\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30818\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35796\,
            DIN => \N__35795\,
            DOUT => \N__35794\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35796\,
            PADOUT => \N__35795\,
            PADIN => \N__35794\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35787\,
            DIN => \N__35786\,
            DOUT => \N__35785\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35787\,
            PADOUT => \N__35786\,
            PADIN => \N__35785\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23135\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35778\,
            DIN => \N__35777\,
            DOUT => \N__35776\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35778\,
            PADOUT => \N__35777\,
            PADIN => \N__35776\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19724\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35769\,
            DIN => \N__35768\,
            DOUT => \N__35767\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35769\,
            PADOUT => \N__35768\,
            PADIN => \N__35767\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35760\,
            DIN => \N__35759\,
            DOUT => \N__35758\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35760\,
            PADOUT => \N__35759\,
            PADIN => \N__35758\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__35751\,
            DIN => \N__35750\,
            DOUT => \N__35749\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35751\,
            PADOUT => \N__35750\,
            PADIN => \N__35749\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35742\,
            DIN => \N__35741\,
            DOUT => \N__35740\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35742\,
            PADOUT => \N__35741\,
            PADIN => \N__35740\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35733\,
            DIN => \N__35732\,
            DOUT => \N__35731\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35733\,
            PADOUT => \N__35732\,
            PADIN => \N__35731\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29732\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35724\,
            DIN => \N__35723\,
            DOUT => \N__35722\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35724\,
            PADOUT => \N__35723\,
            PADIN => \N__35722\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35715\,
            DIN => \N__35714\,
            DOUT => \N__35713\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35715\,
            PADOUT => \N__35714\,
            PADIN => \N__35713\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35706\,
            DIN => \N__35705\,
            DOUT => \N__35704\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35706\,
            PADOUT => \N__35705\,
            PADIN => \N__35704\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35697\,
            DIN => \N__35696\,
            DOUT => \N__35695\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35697\,
            PADOUT => \N__35696\,
            PADIN => \N__35695\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35688\,
            DIN => \N__35687\,
            DOUT => \N__35686\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35688\,
            PADOUT => \N__35687\,
            PADIN => \N__35686\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35679\,
            DIN => \N__35678\,
            DOUT => \N__35677\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35679\,
            PADOUT => \N__35678\,
            PADIN => \N__35677\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35670\,
            DIN => \N__35669\,
            DOUT => \N__35668\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35670\,
            PADOUT => \N__35669\,
            PADIN => \N__35668\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25088\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__35661\,
            DIN => \N__35660\,
            DOUT => \N__35659\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__35661\,
            PADOUT => \N__35660\,
            PADIN => \N__35659\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__8387\ : InMux
    port map (
            O => \N__35642\,
            I => \N__35638\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__35641\,
            I => \N__35630\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__35638\,
            I => \N__35626\
        );

    \I__8384\ : InMux
    port map (
            O => \N__35637\,
            I => \N__35614\
        );

    \I__8383\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35614\
        );

    \I__8382\ : InMux
    port map (
            O => \N__35635\,
            I => \N__35614\
        );

    \I__8381\ : InMux
    port map (
            O => \N__35634\,
            I => \N__35614\
        );

    \I__8380\ : InMux
    port map (
            O => \N__35633\,
            I => \N__35614\
        );

    \I__8379\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35611\
        );

    \I__8378\ : InMux
    port map (
            O => \N__35629\,
            I => \N__35608\
        );

    \I__8377\ : Span4Mux_v
    port map (
            O => \N__35626\,
            I => \N__35605\
        );

    \I__8376\ : InMux
    port map (
            O => \N__35625\,
            I => \N__35602\
        );

    \I__8375\ : LocalMux
    port map (
            O => \N__35614\,
            I => \N__35597\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__35611\,
            I => \N__35597\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__35608\,
            I => \N__35594\
        );

    \I__8372\ : Span4Mux_v
    port map (
            O => \N__35605\,
            I => \N__35591\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__35602\,
            I => \N__35586\
        );

    \I__8370\ : Sp12to4
    port map (
            O => \N__35597\,
            I => \N__35586\
        );

    \I__8369\ : Span4Mux_s2_h
    port map (
            O => \N__35594\,
            I => \N__35583\
        );

    \I__8368\ : Odrv4
    port map (
            O => \N__35591\,
            I => \count_clk_RNINSEUC_0_6\
        );

    \I__8367\ : Odrv12
    port map (
            O => \N__35586\,
            I => \count_clk_RNINSEUC_0_6\
        );

    \I__8366\ : Odrv4
    port map (
            O => \N__35583\,
            I => \count_clk_RNINSEUC_0_6\
        );

    \I__8365\ : InMux
    port map (
            O => \N__35576\,
            I => \N__35572\
        );

    \I__8364\ : CascadeMux
    port map (
            O => \N__35575\,
            I => \N__35569\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__35572\,
            I => \N__35565\
        );

    \I__8362\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35562\
        );

    \I__8361\ : CascadeMux
    port map (
            O => \N__35568\,
            I => \N__35558\
        );

    \I__8360\ : Span4Mux_v
    port map (
            O => \N__35565\,
            I => \N__35552\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__35562\,
            I => \N__35552\
        );

    \I__8358\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35548\
        );

    \I__8357\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35545\
        );

    \I__8356\ : InMux
    port map (
            O => \N__35557\,
            I => \N__35542\
        );

    \I__8355\ : Span4Mux_h
    port map (
            O => \N__35552\,
            I => \N__35537\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__35551\,
            I => \N__35534\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__35548\,
            I => \N__35526\
        );

    \I__8352\ : LocalMux
    port map (
            O => \N__35545\,
            I => \N__35526\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__35542\,
            I => \N__35526\
        );

    \I__8350\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35523\
        );

    \I__8349\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35520\
        );

    \I__8348\ : Span4Mux_v
    port map (
            O => \N__35537\,
            I => \N__35517\
        );

    \I__8347\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35512\
        );

    \I__8346\ : InMux
    port map (
            O => \N__35533\,
            I => \N__35512\
        );

    \I__8345\ : Span4Mux_v
    port map (
            O => \N__35526\,
            I => \N__35507\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__35523\,
            I => \N__35507\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35504\
        );

    \I__8342\ : Odrv4
    port map (
            O => \N__35517\,
            I => \POWERLED.N_412_i\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__35512\,
            I => \POWERLED.N_412_i\
        );

    \I__8340\ : Odrv4
    port map (
            O => \N__35507\,
            I => \POWERLED.N_412_i\
        );

    \I__8339\ : Odrv12
    port map (
            O => \N__35504\,
            I => \POWERLED.N_412_i\
        );

    \I__8338\ : CascadeMux
    port map (
            O => \N__35495\,
            I => \N__35492\
        );

    \I__8337\ : InMux
    port map (
            O => \N__35492\,
            I => \N__35485\
        );

    \I__8336\ : InMux
    port map (
            O => \N__35491\,
            I => \N__35485\
        );

    \I__8335\ : CascadeMux
    port map (
            O => \N__35490\,
            I => \N__35482\
        );

    \I__8334\ : LocalMux
    port map (
            O => \N__35485\,
            I => \N__35477\
        );

    \I__8333\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35467\
        );

    \I__8332\ : InMux
    port map (
            O => \N__35481\,
            I => \N__35462\
        );

    \I__8331\ : InMux
    port map (
            O => \N__35480\,
            I => \N__35462\
        );

    \I__8330\ : Span4Mux_v
    port map (
            O => \N__35477\,
            I => \N__35459\
        );

    \I__8329\ : CascadeMux
    port map (
            O => \N__35476\,
            I => \N__35454\
        );

    \I__8328\ : CascadeMux
    port map (
            O => \N__35475\,
            I => \N__35451\
        );

    \I__8327\ : InMux
    port map (
            O => \N__35474\,
            I => \N__35439\
        );

    \I__8326\ : InMux
    port map (
            O => \N__35473\,
            I => \N__35430\
        );

    \I__8325\ : InMux
    port map (
            O => \N__35472\,
            I => \N__35430\
        );

    \I__8324\ : InMux
    port map (
            O => \N__35471\,
            I => \N__35430\
        );

    \I__8323\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35430\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__35467\,
            I => \N__35425\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__35462\,
            I => \N__35425\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__35459\,
            I => \N__35422\
        );

    \I__8319\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35419\
        );

    \I__8318\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35416\
        );

    \I__8317\ : InMux
    port map (
            O => \N__35454\,
            I => \N__35413\
        );

    \I__8316\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35410\
        );

    \I__8315\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35404\
        );

    \I__8314\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35404\
        );

    \I__8313\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35394\
        );

    \I__8312\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35394\
        );

    \I__8311\ : InMux
    port map (
            O => \N__35446\,
            I => \N__35394\
        );

    \I__8310\ : InMux
    port map (
            O => \N__35445\,
            I => \N__35394\
        );

    \I__8309\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35391\
        );

    \I__8308\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35385\
        );

    \I__8307\ : InMux
    port map (
            O => \N__35442\,
            I => \N__35385\
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__35439\,
            I => \N__35380\
        );

    \I__8305\ : LocalMux
    port map (
            O => \N__35430\,
            I => \N__35380\
        );

    \I__8304\ : Span4Mux_v
    port map (
            O => \N__35425\,
            I => \N__35374\
        );

    \I__8303\ : Span4Mux_h
    port map (
            O => \N__35422\,
            I => \N__35369\
        );

    \I__8302\ : LocalMux
    port map (
            O => \N__35419\,
            I => \N__35369\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__35416\,
            I => \N__35366\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__35413\,
            I => \N__35361\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__35410\,
            I => \N__35361\
        );

    \I__8298\ : InMux
    port map (
            O => \N__35409\,
            I => \N__35358\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__35404\,
            I => \N__35355\
        );

    \I__8296\ : InMux
    port map (
            O => \N__35403\,
            I => \N__35352\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__35394\,
            I => \N__35346\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__35391\,
            I => \N__35346\
        );

    \I__8293\ : CascadeMux
    port map (
            O => \N__35390\,
            I => \N__35341\
        );

    \I__8292\ : LocalMux
    port map (
            O => \N__35385\,
            I => \N__35337\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__35380\,
            I => \N__35334\
        );

    \I__8290\ : InMux
    port map (
            O => \N__35379\,
            I => \N__35331\
        );

    \I__8289\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35326\
        );

    \I__8288\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35326\
        );

    \I__8287\ : IoSpan4Mux
    port map (
            O => \N__35374\,
            I => \N__35321\
        );

    \I__8286\ : Span4Mux_v
    port map (
            O => \N__35369\,
            I => \N__35318\
        );

    \I__8285\ : Span4Mux_v
    port map (
            O => \N__35366\,
            I => \N__35311\
        );

    \I__8284\ : Span4Mux_v
    port map (
            O => \N__35361\,
            I => \N__35311\
        );

    \I__8283\ : LocalMux
    port map (
            O => \N__35358\,
            I => \N__35311\
        );

    \I__8282\ : Span4Mux_h
    port map (
            O => \N__35355\,
            I => \N__35308\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__35352\,
            I => \N__35305\
        );

    \I__8280\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35302\
        );

    \I__8279\ : Span4Mux_s1_h
    port map (
            O => \N__35346\,
            I => \N__35299\
        );

    \I__8278\ : InMux
    port map (
            O => \N__35345\,
            I => \N__35294\
        );

    \I__8277\ : InMux
    port map (
            O => \N__35344\,
            I => \N__35294\
        );

    \I__8276\ : InMux
    port map (
            O => \N__35341\,
            I => \N__35289\
        );

    \I__8275\ : InMux
    port map (
            O => \N__35340\,
            I => \N__35289\
        );

    \I__8274\ : Span4Mux_v
    port map (
            O => \N__35337\,
            I => \N__35286\
        );

    \I__8273\ : Span4Mux_v
    port map (
            O => \N__35334\,
            I => \N__35279\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__35331\,
            I => \N__35279\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__35326\,
            I => \N__35279\
        );

    \I__8270\ : InMux
    port map (
            O => \N__35325\,
            I => \N__35276\
        );

    \I__8269\ : InMux
    port map (
            O => \N__35324\,
            I => \N__35273\
        );

    \I__8268\ : IoSpan4Mux
    port map (
            O => \N__35321\,
            I => \N__35269\
        );

    \I__8267\ : Span4Mux_s2_v
    port map (
            O => \N__35318\,
            I => \N__35264\
        );

    \I__8266\ : Span4Mux_v
    port map (
            O => \N__35311\,
            I => \N__35264\
        );

    \I__8265\ : Span4Mux_v
    port map (
            O => \N__35308\,
            I => \N__35259\
        );

    \I__8264\ : Span4Mux_s1_h
    port map (
            O => \N__35305\,
            I => \N__35259\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__35302\,
            I => \N__35256\
        );

    \I__8262\ : Span4Mux_v
    port map (
            O => \N__35299\,
            I => \N__35249\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__35294\,
            I => \N__35249\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__35289\,
            I => \N__35249\
        );

    \I__8259\ : Span4Mux_h
    port map (
            O => \N__35286\,
            I => \N__35240\
        );

    \I__8258\ : Span4Mux_v
    port map (
            O => \N__35279\,
            I => \N__35240\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__35276\,
            I => \N__35240\
        );

    \I__8256\ : LocalMux
    port map (
            O => \N__35273\,
            I => \N__35240\
        );

    \I__8255\ : InMux
    port map (
            O => \N__35272\,
            I => \N__35237\
        );

    \I__8254\ : IoSpan4Mux
    port map (
            O => \N__35269\,
            I => \N__35232\
        );

    \I__8253\ : IoSpan4Mux
    port map (
            O => \N__35264\,
            I => \N__35232\
        );

    \I__8252\ : Span4Mux_v
    port map (
            O => \N__35259\,
            I => \N__35225\
        );

    \I__8251\ : Span4Mux_s1_h
    port map (
            O => \N__35256\,
            I => \N__35225\
        );

    \I__8250\ : Span4Mux_v
    port map (
            O => \N__35249\,
            I => \N__35225\
        );

    \I__8249\ : Span4Mux_v
    port map (
            O => \N__35240\,
            I => \N__35220\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__35237\,
            I => \N__35220\
        );

    \I__8247\ : Odrv4
    port map (
            O => \N__35232\,
            I => slp_s3n
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__35225\,
            I => slp_s3n
        );

    \I__8245\ : Odrv4
    port map (
            O => \N__35220\,
            I => slp_s3n
        );

    \I__8244\ : InMux
    port map (
            O => \N__35213\,
            I => \N__35210\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__35210\,
            I => \N__35203\
        );

    \I__8242\ : InMux
    port map (
            O => \N__35209\,
            I => \N__35200\
        );

    \I__8241\ : InMux
    port map (
            O => \N__35208\,
            I => \N__35195\
        );

    \I__8240\ : InMux
    port map (
            O => \N__35207\,
            I => \N__35195\
        );

    \I__8239\ : CascadeMux
    port map (
            O => \N__35206\,
            I => \N__35191\
        );

    \I__8238\ : Span4Mux_v
    port map (
            O => \N__35203\,
            I => \N__35188\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__35200\,
            I => \N__35183\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__35195\,
            I => \N__35183\
        );

    \I__8235\ : InMux
    port map (
            O => \N__35194\,
            I => \N__35180\
        );

    \I__8234\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35177\
        );

    \I__8233\ : Span4Mux_v
    port map (
            O => \N__35188\,
            I => \N__35172\
        );

    \I__8232\ : Sp12to4
    port map (
            O => \N__35183\,
            I => \N__35165\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__35180\,
            I => \N__35165\
        );

    \I__8230\ : LocalMux
    port map (
            O => \N__35177\,
            I => \N__35165\
        );

    \I__8229\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35160\
        );

    \I__8228\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35160\
        );

    \I__8227\ : Odrv4
    port map (
            O => \N__35172\,
            I => \POWERLED.N_251\
        );

    \I__8226\ : Odrv12
    port map (
            O => \N__35165\,
            I => \POWERLED.N_251\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__35160\,
            I => \POWERLED.N_251\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__35153\,
            I => \N__35149\
        );

    \I__8223\ : IoInMux
    port map (
            O => \N__35152\,
            I => \N__35145\
        );

    \I__8222\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35139\
        );

    \I__8221\ : CascadeMux
    port map (
            O => \N__35148\,
            I => \N__35136\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__35145\,
            I => \N__35132\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__35144\,
            I => \N__35128\
        );

    \I__8218\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35123\
        );

    \I__8217\ : InMux
    port map (
            O => \N__35142\,
            I => \N__35120\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__35139\,
            I => \N__35115\
        );

    \I__8215\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35112\
        );

    \I__8214\ : CascadeMux
    port map (
            O => \N__35135\,
            I => \N__35107\
        );

    \I__8213\ : Span4Mux_s3_v
    port map (
            O => \N__35132\,
            I => \N__35104\
        );

    \I__8212\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35101\
        );

    \I__8211\ : InMux
    port map (
            O => \N__35128\,
            I => \N__35098\
        );

    \I__8210\ : InMux
    port map (
            O => \N__35127\,
            I => \N__35094\
        );

    \I__8209\ : InMux
    port map (
            O => \N__35126\,
            I => \N__35091\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__35123\,
            I => \N__35086\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__35120\,
            I => \N__35086\
        );

    \I__8206\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35082\
        );

    \I__8205\ : InMux
    port map (
            O => \N__35118\,
            I => \N__35079\
        );

    \I__8204\ : Span4Mux_s1_h
    port map (
            O => \N__35115\,
            I => \N__35074\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__35112\,
            I => \N__35074\
        );

    \I__8202\ : InMux
    port map (
            O => \N__35111\,
            I => \N__35071\
        );

    \I__8201\ : InMux
    port map (
            O => \N__35110\,
            I => \N__35068\
        );

    \I__8200\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35065\
        );

    \I__8199\ : Span4Mux_v
    port map (
            O => \N__35104\,
            I => \N__35060\
        );

    \I__8198\ : LocalMux
    port map (
            O => \N__35101\,
            I => \N__35060\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__35098\,
            I => \N__35057\
        );

    \I__8196\ : InMux
    port map (
            O => \N__35097\,
            I => \N__35054\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__35094\,
            I => \N__35051\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__35091\,
            I => \N__35044\
        );

    \I__8193\ : Span4Mux_s3_h
    port map (
            O => \N__35086\,
            I => \N__35044\
        );

    \I__8192\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35041\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__35082\,
            I => \N__35036\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__35079\,
            I => \N__35036\
        );

    \I__8189\ : Span4Mux_v
    port map (
            O => \N__35074\,
            I => \N__35031\
        );

    \I__8188\ : LocalMux
    port map (
            O => \N__35071\,
            I => \N__35031\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__35068\,
            I => \N__35028\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__35065\,
            I => \N__35025\
        );

    \I__8185\ : Span4Mux_h
    port map (
            O => \N__35060\,
            I => \N__35018\
        );

    \I__8184\ : Span4Mux_h
    port map (
            O => \N__35057\,
            I => \N__35018\
        );

    \I__8183\ : LocalMux
    port map (
            O => \N__35054\,
            I => \N__35018\
        );

    \I__8182\ : Span4Mux_s3_h
    port map (
            O => \N__35051\,
            I => \N__35015\
        );

    \I__8181\ : InMux
    port map (
            O => \N__35050\,
            I => \N__35012\
        );

    \I__8180\ : InMux
    port map (
            O => \N__35049\,
            I => \N__35009\
        );

    \I__8179\ : Span4Mux_v
    port map (
            O => \N__35044\,
            I => \N__35004\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__35041\,
            I => \N__35004\
        );

    \I__8177\ : Span4Mux_v
    port map (
            O => \N__35036\,
            I => \N__34995\
        );

    \I__8176\ : Span4Mux_v
    port map (
            O => \N__35031\,
            I => \N__34995\
        );

    \I__8175\ : Span4Mux_s1_h
    port map (
            O => \N__35028\,
            I => \N__34995\
        );

    \I__8174\ : Span4Mux_s1_h
    port map (
            O => \N__35025\,
            I => \N__34995\
        );

    \I__8173\ : Span4Mux_v
    port map (
            O => \N__35018\,
            I => \N__34992\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__35015\,
            I => \N__34987\
        );

    \I__8171\ : LocalMux
    port map (
            O => \N__35012\,
            I => \N__34987\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__35009\,
            I => \N__34982\
        );

    \I__8169\ : Span4Mux_v
    port map (
            O => \N__35004\,
            I => \N__34982\
        );

    \I__8168\ : Span4Mux_v
    port map (
            O => \N__34995\,
            I => \N__34977\
        );

    \I__8167\ : Span4Mux_v
    port map (
            O => \N__34992\,
            I => \N__34977\
        );

    \I__8166\ : Odrv4
    port map (
            O => \N__34987\,
            I => rsmrstn
        );

    \I__8165\ : Odrv4
    port map (
            O => \N__34982\,
            I => rsmrstn
        );

    \I__8164\ : Odrv4
    port map (
            O => \N__34977\,
            I => rsmrstn
        );

    \I__8163\ : CascadeMux
    port map (
            O => \N__34970\,
            I => \N__34964\
        );

    \I__8162\ : InMux
    port map (
            O => \N__34969\,
            I => \N__34961\
        );

    \I__8161\ : CascadeMux
    port map (
            O => \N__34968\,
            I => \N__34956\
        );

    \I__8160\ : CascadeMux
    port map (
            O => \N__34967\,
            I => \N__34953\
        );

    \I__8159\ : InMux
    port map (
            O => \N__34964\,
            I => \N__34950\
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__34961\,
            I => \N__34947\
        );

    \I__8157\ : InMux
    port map (
            O => \N__34960\,
            I => \N__34944\
        );

    \I__8156\ : InMux
    port map (
            O => \N__34959\,
            I => \N__34941\
        );

    \I__8155\ : InMux
    port map (
            O => \N__34956\,
            I => \N__34938\
        );

    \I__8154\ : InMux
    port map (
            O => \N__34953\,
            I => \N__34931\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__34950\,
            I => \N__34928\
        );

    \I__8152\ : Span4Mux_v
    port map (
            O => \N__34947\,
            I => \N__34925\
        );

    \I__8151\ : LocalMux
    port map (
            O => \N__34944\,
            I => \N__34918\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__34941\,
            I => \N__34918\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__34938\,
            I => \N__34918\
        );

    \I__8148\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34915\
        );

    \I__8147\ : InMux
    port map (
            O => \N__34936\,
            I => \N__34912\
        );

    \I__8146\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34909\
        );

    \I__8145\ : InMux
    port map (
            O => \N__34934\,
            I => \N__34906\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__34931\,
            I => \N__34901\
        );

    \I__8143\ : Span4Mux_s3_h
    port map (
            O => \N__34928\,
            I => \N__34901\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__34925\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8141\ : Odrv12
    port map (
            O => \N__34918\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8140\ : LocalMux
    port map (
            O => \N__34915\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__34912\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8138\ : LocalMux
    port map (
            O => \N__34909\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__34906\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__34901\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__8135\ : InMux
    port map (
            O => \N__34886\,
            I => \N__34883\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__34883\,
            I => \POWERLED.N_524\
        );

    \I__8133\ : CascadeMux
    port map (
            O => \N__34880\,
            I => \N__34876\
        );

    \I__8132\ : CascadeMux
    port map (
            O => \N__34879\,
            I => \N__34873\
        );

    \I__8131\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34869\
        );

    \I__8130\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34866\
        );

    \I__8129\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34861\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__34869\,
            I => \N__34858\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__34866\,
            I => \N__34855\
        );

    \I__8126\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34850\
        );

    \I__8125\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34850\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34847\
        );

    \I__8123\ : Span4Mux_h
    port map (
            O => \N__34858\,
            I => \N__34844\
        );

    \I__8122\ : Odrv4
    port map (
            O => \N__34855\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__8121\ : LocalMux
    port map (
            O => \N__34850\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__8120\ : Odrv4
    port map (
            O => \N__34847\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__34844\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__8118\ : InMux
    port map (
            O => \N__34835\,
            I => \N__34821\
        );

    \I__8117\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34821\
        );

    \I__8116\ : InMux
    port map (
            O => \N__34833\,
            I => \N__34821\
        );

    \I__8115\ : InMux
    port map (
            O => \N__34832\,
            I => \N__34821\
        );

    \I__8114\ : InMux
    port map (
            O => \N__34831\,
            I => \N__34816\
        );

    \I__8113\ : InMux
    port map (
            O => \N__34830\,
            I => \N__34816\
        );

    \I__8112\ : LocalMux
    port map (
            O => \N__34821\,
            I => \N__34803\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__34816\,
            I => \N__34803\
        );

    \I__8110\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34794\
        );

    \I__8109\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34794\
        );

    \I__8108\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34794\
        );

    \I__8107\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34794\
        );

    \I__8106\ : InMux
    port map (
            O => \N__34811\,
            I => \N__34787\
        );

    \I__8105\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34787\
        );

    \I__8104\ : InMux
    port map (
            O => \N__34809\,
            I => \N__34787\
        );

    \I__8103\ : InMux
    port map (
            O => \N__34808\,
            I => \N__34779\
        );

    \I__8102\ : Span4Mux_s1_v
    port map (
            O => \N__34803\,
            I => \N__34772\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__34794\,
            I => \N__34772\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__34787\,
            I => \N__34772\
        );

    \I__8099\ : InMux
    port map (
            O => \N__34786\,
            I => \N__34761\
        );

    \I__8098\ : InMux
    port map (
            O => \N__34785\,
            I => \N__34761\
        );

    \I__8097\ : InMux
    port map (
            O => \N__34784\,
            I => \N__34761\
        );

    \I__8096\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34761\
        );

    \I__8095\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34761\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__34779\,
            I => \POWERLED.func_state_RNIUQMRH_0_1\
        );

    \I__8093\ : Odrv4
    port map (
            O => \N__34772\,
            I => \POWERLED.func_state_RNIUQMRH_0_1\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__34761\,
            I => \POWERLED.func_state_RNIUQMRH_0_1\
        );

    \I__8091\ : InMux
    port map (
            O => \N__34754\,
            I => \N__34751\
        );

    \I__8090\ : LocalMux
    port map (
            O => \N__34751\,
            I => \N__34748\
        );

    \I__8089\ : Span4Mux_s2_v
    port map (
            O => \N__34748\,
            I => \N__34745\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__34745\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__8087\ : ClkMux
    port map (
            O => \N__34742\,
            I => \N__34734\
        );

    \I__8086\ : ClkMux
    port map (
            O => \N__34741\,
            I => \N__34731\
        );

    \I__8085\ : ClkMux
    port map (
            O => \N__34740\,
            I => \N__34728\
        );

    \I__8084\ : ClkMux
    port map (
            O => \N__34739\,
            I => \N__34721\
        );

    \I__8083\ : ClkMux
    port map (
            O => \N__34738\,
            I => \N__34712\
        );

    \I__8082\ : ClkMux
    port map (
            O => \N__34737\,
            I => \N__34709\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__34734\,
            I => \N__34705\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__34731\,
            I => \N__34702\
        );

    \I__8079\ : LocalMux
    port map (
            O => \N__34728\,
            I => \N__34696\
        );

    \I__8078\ : ClkMux
    port map (
            O => \N__34727\,
            I => \N__34693\
        );

    \I__8077\ : ClkMux
    port map (
            O => \N__34726\,
            I => \N__34690\
        );

    \I__8076\ : ClkMux
    port map (
            O => \N__34725\,
            I => \N__34687\
        );

    \I__8075\ : ClkMux
    port map (
            O => \N__34724\,
            I => \N__34682\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__34721\,
            I => \N__34673\
        );

    \I__8073\ : ClkMux
    port map (
            O => \N__34720\,
            I => \N__34670\
        );

    \I__8072\ : ClkMux
    port map (
            O => \N__34719\,
            I => \N__34667\
        );

    \I__8071\ : ClkMux
    port map (
            O => \N__34718\,
            I => \N__34664\
        );

    \I__8070\ : ClkMux
    port map (
            O => \N__34717\,
            I => \N__34661\
        );

    \I__8069\ : ClkMux
    port map (
            O => \N__34716\,
            I => \N__34657\
        );

    \I__8068\ : ClkMux
    port map (
            O => \N__34715\,
            I => \N__34652\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__34712\,
            I => \N__34645\
        );

    \I__8066\ : LocalMux
    port map (
            O => \N__34709\,
            I => \N__34645\
        );

    \I__8065\ : ClkMux
    port map (
            O => \N__34708\,
            I => \N__34642\
        );

    \I__8064\ : Span4Mux_v
    port map (
            O => \N__34705\,
            I => \N__34639\
        );

    \I__8063\ : Span4Mux_s3_h
    port map (
            O => \N__34702\,
            I => \N__34636\
        );

    \I__8062\ : ClkMux
    port map (
            O => \N__34701\,
            I => \N__34633\
        );

    \I__8061\ : ClkMux
    port map (
            O => \N__34700\,
            I => \N__34630\
        );

    \I__8060\ : ClkMux
    port map (
            O => \N__34699\,
            I => \N__34627\
        );

    \I__8059\ : Span4Mux_v
    port map (
            O => \N__34696\,
            I => \N__34622\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__34693\,
            I => \N__34622\
        );

    \I__8057\ : LocalMux
    port map (
            O => \N__34690\,
            I => \N__34616\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__34687\,
            I => \N__34616\
        );

    \I__8055\ : ClkMux
    port map (
            O => \N__34686\,
            I => \N__34613\
        );

    \I__8054\ : ClkMux
    port map (
            O => \N__34685\,
            I => \N__34610\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__34682\,
            I => \N__34607\
        );

    \I__8052\ : ClkMux
    port map (
            O => \N__34681\,
            I => \N__34604\
        );

    \I__8051\ : ClkMux
    port map (
            O => \N__34680\,
            I => \N__34601\
        );

    \I__8050\ : ClkMux
    port map (
            O => \N__34679\,
            I => \N__34597\
        );

    \I__8049\ : ClkMux
    port map (
            O => \N__34678\,
            I => \N__34593\
        );

    \I__8048\ : ClkMux
    port map (
            O => \N__34677\,
            I => \N__34589\
        );

    \I__8047\ : ClkMux
    port map (
            O => \N__34676\,
            I => \N__34586\
        );

    \I__8046\ : Span4Mux_s2_v
    port map (
            O => \N__34673\,
            I => \N__34577\
        );

    \I__8045\ : LocalMux
    port map (
            O => \N__34670\,
            I => \N__34577\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__34667\,
            I => \N__34574\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__34664\,
            I => \N__34570\
        );

    \I__8042\ : LocalMux
    port map (
            O => \N__34661\,
            I => \N__34567\
        );

    \I__8041\ : ClkMux
    port map (
            O => \N__34660\,
            I => \N__34564\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__34657\,
            I => \N__34561\
        );

    \I__8039\ : ClkMux
    port map (
            O => \N__34656\,
            I => \N__34558\
        );

    \I__8038\ : ClkMux
    port map (
            O => \N__34655\,
            I => \N__34554\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__34652\,
            I => \N__34547\
        );

    \I__8036\ : ClkMux
    port map (
            O => \N__34651\,
            I => \N__34544\
        );

    \I__8035\ : ClkMux
    port map (
            O => \N__34650\,
            I => \N__34541\
        );

    \I__8034\ : Span4Mux_s3_v
    port map (
            O => \N__34645\,
            I => \N__34534\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__34642\,
            I => \N__34534\
        );

    \I__8032\ : Span4Mux_h
    port map (
            O => \N__34639\,
            I => \N__34525\
        );

    \I__8031\ : Span4Mux_h
    port map (
            O => \N__34636\,
            I => \N__34525\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__34633\,
            I => \N__34525\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__34630\,
            I => \N__34522\
        );

    \I__8028\ : LocalMux
    port map (
            O => \N__34627\,
            I => \N__34517\
        );

    \I__8027\ : Span4Mux_v
    port map (
            O => \N__34622\,
            I => \N__34517\
        );

    \I__8026\ : ClkMux
    port map (
            O => \N__34621\,
            I => \N__34514\
        );

    \I__8025\ : Span4Mux_h
    port map (
            O => \N__34616\,
            I => \N__34506\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__34613\,
            I => \N__34506\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__34610\,
            I => \N__34506\
        );

    \I__8022\ : Span4Mux_s1_v
    port map (
            O => \N__34607\,
            I => \N__34499\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__34604\,
            I => \N__34499\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__34601\,
            I => \N__34499\
        );

    \I__8019\ : ClkMux
    port map (
            O => \N__34600\,
            I => \N__34496\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__34597\,
            I => \N__34492\
        );

    \I__8017\ : ClkMux
    port map (
            O => \N__34596\,
            I => \N__34486\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__34593\,
            I => \N__34483\
        );

    \I__8015\ : ClkMux
    port map (
            O => \N__34592\,
            I => \N__34480\
        );

    \I__8014\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34475\
        );

    \I__8013\ : LocalMux
    port map (
            O => \N__34586\,
            I => \N__34475\
        );

    \I__8012\ : ClkMux
    port map (
            O => \N__34585\,
            I => \N__34472\
        );

    \I__8011\ : ClkMux
    port map (
            O => \N__34584\,
            I => \N__34469\
        );

    \I__8010\ : ClkMux
    port map (
            O => \N__34583\,
            I => \N__34466\
        );

    \I__8009\ : ClkMux
    port map (
            O => \N__34582\,
            I => \N__34460\
        );

    \I__8008\ : Span4Mux_v
    port map (
            O => \N__34577\,
            I => \N__34455\
        );

    \I__8007\ : Span4Mux_s1_h
    port map (
            O => \N__34574\,
            I => \N__34455\
        );

    \I__8006\ : ClkMux
    port map (
            O => \N__34573\,
            I => \N__34452\
        );

    \I__8005\ : Span4Mux_s2_v
    port map (
            O => \N__34570\,
            I => \N__34444\
        );

    \I__8004\ : Span4Mux_s2_h
    port map (
            O => \N__34567\,
            I => \N__34444\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__34564\,
            I => \N__34444\
        );

    \I__8002\ : Span4Mux_s1_h
    port map (
            O => \N__34561\,
            I => \N__34439\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__34558\,
            I => \N__34439\
        );

    \I__8000\ : ClkMux
    port map (
            O => \N__34557\,
            I => \N__34436\
        );

    \I__7999\ : LocalMux
    port map (
            O => \N__34554\,
            I => \N__34433\
        );

    \I__7998\ : ClkMux
    port map (
            O => \N__34553\,
            I => \N__34430\
        );

    \I__7997\ : ClkMux
    port map (
            O => \N__34552\,
            I => \N__34427\
        );

    \I__7996\ : ClkMux
    port map (
            O => \N__34551\,
            I => \N__34420\
        );

    \I__7995\ : ClkMux
    port map (
            O => \N__34550\,
            I => \N__34417\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__34547\,
            I => \N__34409\
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34409\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34409\
        );

    \I__7991\ : ClkMux
    port map (
            O => \N__34540\,
            I => \N__34406\
        );

    \I__7990\ : ClkMux
    port map (
            O => \N__34539\,
            I => \N__34400\
        );

    \I__7989\ : Span4Mux_v
    port map (
            O => \N__34534\,
            I => \N__34395\
        );

    \I__7988\ : ClkMux
    port map (
            O => \N__34533\,
            I => \N__34392\
        );

    \I__7987\ : ClkMux
    port map (
            O => \N__34532\,
            I => \N__34389\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__34525\,
            I => \N__34380\
        );

    \I__7985\ : Span4Mux_h
    port map (
            O => \N__34522\,
            I => \N__34380\
        );

    \I__7984\ : Span4Mux_h
    port map (
            O => \N__34517\,
            I => \N__34380\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__34514\,
            I => \N__34380\
        );

    \I__7982\ : ClkMux
    port map (
            O => \N__34513\,
            I => \N__34377\
        );

    \I__7981\ : Span4Mux_v
    port map (
            O => \N__34506\,
            I => \N__34370\
        );

    \I__7980\ : Span4Mux_v
    port map (
            O => \N__34499\,
            I => \N__34370\
        );

    \I__7979\ : LocalMux
    port map (
            O => \N__34496\,
            I => \N__34370\
        );

    \I__7978\ : ClkMux
    port map (
            O => \N__34495\,
            I => \N__34367\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__34492\,
            I => \N__34364\
        );

    \I__7976\ : ClkMux
    port map (
            O => \N__34491\,
            I => \N__34361\
        );

    \I__7975\ : ClkMux
    port map (
            O => \N__34490\,
            I => \N__34358\
        );

    \I__7974\ : ClkMux
    port map (
            O => \N__34489\,
            I => \N__34355\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__34486\,
            I => \N__34347\
        );

    \I__7972\ : Span4Mux_h
    port map (
            O => \N__34483\,
            I => \N__34347\
        );

    \I__7971\ : LocalMux
    port map (
            O => \N__34480\,
            I => \N__34347\
        );

    \I__7970\ : Span4Mux_v
    port map (
            O => \N__34475\,
            I => \N__34340\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__34472\,
            I => \N__34340\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__34469\,
            I => \N__34340\
        );

    \I__7967\ : LocalMux
    port map (
            O => \N__34466\,
            I => \N__34337\
        );

    \I__7966\ : ClkMux
    port map (
            O => \N__34465\,
            I => \N__34334\
        );

    \I__7965\ : ClkMux
    port map (
            O => \N__34464\,
            I => \N__34330\
        );

    \I__7964\ : ClkMux
    port map (
            O => \N__34463\,
            I => \N__34327\
        );

    \I__7963\ : LocalMux
    port map (
            O => \N__34460\,
            I => \N__34323\
        );

    \I__7962\ : Span4Mux_v
    port map (
            O => \N__34455\,
            I => \N__34318\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__34452\,
            I => \N__34318\
        );

    \I__7960\ : ClkMux
    port map (
            O => \N__34451\,
            I => \N__34315\
        );

    \I__7959\ : Span4Mux_v
    port map (
            O => \N__34444\,
            I => \N__34312\
        );

    \I__7958\ : Span4Mux_h
    port map (
            O => \N__34439\,
            I => \N__34307\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__34436\,
            I => \N__34307\
        );

    \I__7956\ : Span4Mux_s2_v
    port map (
            O => \N__34433\,
            I => \N__34300\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__34430\,
            I => \N__34300\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__34427\,
            I => \N__34300\
        );

    \I__7953\ : ClkMux
    port map (
            O => \N__34426\,
            I => \N__34297\
        );

    \I__7952\ : ClkMux
    port map (
            O => \N__34425\,
            I => \N__34294\
        );

    \I__7951\ : ClkMux
    port map (
            O => \N__34424\,
            I => \N__34290\
        );

    \I__7950\ : ClkMux
    port map (
            O => \N__34423\,
            I => \N__34287\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34283\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__34417\,
            I => \N__34280\
        );

    \I__7947\ : ClkMux
    port map (
            O => \N__34416\,
            I => \N__34277\
        );

    \I__7946\ : Span4Mux_v
    port map (
            O => \N__34409\,
            I => \N__34272\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__34406\,
            I => \N__34272\
        );

    \I__7944\ : ClkMux
    port map (
            O => \N__34405\,
            I => \N__34269\
        );

    \I__7943\ : ClkMux
    port map (
            O => \N__34404\,
            I => \N__34266\
        );

    \I__7942\ : ClkMux
    port map (
            O => \N__34403\,
            I => \N__34261\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__34400\,
            I => \N__34258\
        );

    \I__7940\ : ClkMux
    port map (
            O => \N__34399\,
            I => \N__34255\
        );

    \I__7939\ : ClkMux
    port map (
            O => \N__34398\,
            I => \N__34251\
        );

    \I__7938\ : Span4Mux_v
    port map (
            O => \N__34395\,
            I => \N__34246\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__34392\,
            I => \N__34246\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__34389\,
            I => \N__34242\
        );

    \I__7935\ : Span4Mux_v
    port map (
            O => \N__34380\,
            I => \N__34239\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__34377\,
            I => \N__34236\
        );

    \I__7933\ : Span4Mux_v
    port map (
            O => \N__34370\,
            I => \N__34227\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__34367\,
            I => \N__34227\
        );

    \I__7931\ : Span4Mux_s2_v
    port map (
            O => \N__34364\,
            I => \N__34227\
        );

    \I__7930\ : LocalMux
    port map (
            O => \N__34361\,
            I => \N__34227\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__34358\,
            I => \N__34222\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__34355\,
            I => \N__34222\
        );

    \I__7927\ : ClkMux
    port map (
            O => \N__34354\,
            I => \N__34219\
        );

    \I__7926\ : Span4Mux_v
    port map (
            O => \N__34347\,
            I => \N__34210\
        );

    \I__7925\ : Span4Mux_v
    port map (
            O => \N__34340\,
            I => \N__34210\
        );

    \I__7924\ : Span4Mux_s3_h
    port map (
            O => \N__34337\,
            I => \N__34210\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__34334\,
            I => \N__34210\
        );

    \I__7922\ : ClkMux
    port map (
            O => \N__34333\,
            I => \N__34207\
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34202\
        );

    \I__7920\ : LocalMux
    port map (
            O => \N__34327\,
            I => \N__34202\
        );

    \I__7919\ : ClkMux
    port map (
            O => \N__34326\,
            I => \N__34199\
        );

    \I__7918\ : Span4Mux_h
    port map (
            O => \N__34323\,
            I => \N__34195\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__34318\,
            I => \N__34190\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__34315\,
            I => \N__34190\
        );

    \I__7915\ : Span4Mux_h
    port map (
            O => \N__34312\,
            I => \N__34179\
        );

    \I__7914\ : Span4Mux_v
    port map (
            O => \N__34307\,
            I => \N__34179\
        );

    \I__7913\ : Span4Mux_v
    port map (
            O => \N__34300\,
            I => \N__34179\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__34297\,
            I => \N__34179\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__34294\,
            I => \N__34179\
        );

    \I__7910\ : ClkMux
    port map (
            O => \N__34293\,
            I => \N__34176\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__34290\,
            I => \N__34173\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__34287\,
            I => \N__34170\
        );

    \I__7907\ : ClkMux
    port map (
            O => \N__34286\,
            I => \N__34167\
        );

    \I__7906\ : Span4Mux_v
    port map (
            O => \N__34283\,
            I => \N__34160\
        );

    \I__7905\ : Span4Mux_h
    port map (
            O => \N__34280\,
            I => \N__34160\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34160\
        );

    \I__7903\ : Span4Mux_v
    port map (
            O => \N__34272\,
            I => \N__34155\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__34269\,
            I => \N__34155\
        );

    \I__7901\ : LocalMux
    port map (
            O => \N__34266\,
            I => \N__34152\
        );

    \I__7900\ : ClkMux
    port map (
            O => \N__34265\,
            I => \N__34149\
        );

    \I__7899\ : ClkMux
    port map (
            O => \N__34264\,
            I => \N__34146\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__34261\,
            I => \N__34143\
        );

    \I__7897\ : Span4Mux_h
    port map (
            O => \N__34258\,
            I => \N__34138\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34138\
        );

    \I__7895\ : ClkMux
    port map (
            O => \N__34254\,
            I => \N__34135\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__34251\,
            I => \N__34130\
        );

    \I__7893\ : Sp12to4
    port map (
            O => \N__34246\,
            I => \N__34130\
        );

    \I__7892\ : ClkMux
    port map (
            O => \N__34245\,
            I => \N__34127\
        );

    \I__7891\ : IoSpan4Mux
    port map (
            O => \N__34242\,
            I => \N__34124\
        );

    \I__7890\ : Span4Mux_h
    port map (
            O => \N__34239\,
            I => \N__34121\
        );

    \I__7889\ : Span4Mux_h
    port map (
            O => \N__34236\,
            I => \N__34112\
        );

    \I__7888\ : Span4Mux_v
    port map (
            O => \N__34227\,
            I => \N__34112\
        );

    \I__7887\ : Span4Mux_v
    port map (
            O => \N__34222\,
            I => \N__34112\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__34219\,
            I => \N__34112\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__34210\,
            I => \N__34107\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__34207\,
            I => \N__34107\
        );

    \I__7883\ : Span4Mux_s2_v
    port map (
            O => \N__34202\,
            I => \N__34104\
        );

    \I__7882\ : LocalMux
    port map (
            O => \N__34199\,
            I => \N__34101\
        );

    \I__7881\ : ClkMux
    port map (
            O => \N__34198\,
            I => \N__34098\
        );

    \I__7880\ : Span4Mux_v
    port map (
            O => \N__34195\,
            I => \N__34089\
        );

    \I__7879\ : Span4Mux_h
    port map (
            O => \N__34190\,
            I => \N__34089\
        );

    \I__7878\ : Span4Mux_v
    port map (
            O => \N__34179\,
            I => \N__34089\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__34176\,
            I => \N__34089\
        );

    \I__7876\ : Span4Mux_s1_h
    port map (
            O => \N__34173\,
            I => \N__34082\
        );

    \I__7875\ : Span4Mux_s1_h
    port map (
            O => \N__34170\,
            I => \N__34082\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34082\
        );

    \I__7873\ : Span4Mux_v
    port map (
            O => \N__34160\,
            I => \N__34071\
        );

    \I__7872\ : Span4Mux_s2_h
    port map (
            O => \N__34155\,
            I => \N__34071\
        );

    \I__7871\ : Span4Mux_s2_h
    port map (
            O => \N__34152\,
            I => \N__34071\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__34149\,
            I => \N__34071\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__34146\,
            I => \N__34071\
        );

    \I__7868\ : Span4Mux_s2_h
    port map (
            O => \N__34143\,
            I => \N__34064\
        );

    \I__7867\ : Span4Mux_h
    port map (
            O => \N__34138\,
            I => \N__34064\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__34135\,
            I => \N__34064\
        );

    \I__7865\ : Span12Mux_s5_h
    port map (
            O => \N__34130\,
            I => \N__34056\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__34127\,
            I => \N__34056\
        );

    \I__7863\ : IoSpan4Mux
    port map (
            O => \N__34124\,
            I => \N__34047\
        );

    \I__7862\ : IoSpan4Mux
    port map (
            O => \N__34121\,
            I => \N__34047\
        );

    \I__7861\ : IoSpan4Mux
    port map (
            O => \N__34112\,
            I => \N__34047\
        );

    \I__7860\ : IoSpan4Mux
    port map (
            O => \N__34107\,
            I => \N__34047\
        );

    \I__7859\ : Span4Mux_h
    port map (
            O => \N__34104\,
            I => \N__34040\
        );

    \I__7858\ : Span4Mux_h
    port map (
            O => \N__34101\,
            I => \N__34040\
        );

    \I__7857\ : LocalMux
    port map (
            O => \N__34098\,
            I => \N__34040\
        );

    \I__7856\ : Span4Mux_v
    port map (
            O => \N__34089\,
            I => \N__34033\
        );

    \I__7855\ : Span4Mux_h
    port map (
            O => \N__34082\,
            I => \N__34033\
        );

    \I__7854\ : Span4Mux_h
    port map (
            O => \N__34071\,
            I => \N__34033\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__34064\,
            I => \N__34030\
        );

    \I__7852\ : ClkMux
    port map (
            O => \N__34063\,
            I => \N__34027\
        );

    \I__7851\ : ClkMux
    port map (
            O => \N__34062\,
            I => \N__34024\
        );

    \I__7850\ : ClkMux
    port map (
            O => \N__34061\,
            I => \N__34021\
        );

    \I__7849\ : Odrv12
    port map (
            O => \N__34056\,
            I => fpga_osc
        );

    \I__7848\ : Odrv4
    port map (
            O => \N__34047\,
            I => fpga_osc
        );

    \I__7847\ : Odrv4
    port map (
            O => \N__34040\,
            I => fpga_osc
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__34033\,
            I => fpga_osc
        );

    \I__7845\ : Odrv4
    port map (
            O => \N__34030\,
            I => fpga_osc
        );

    \I__7844\ : LocalMux
    port map (
            O => \N__34027\,
            I => fpga_osc
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__34024\,
            I => fpga_osc
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__34021\,
            I => fpga_osc
        );

    \I__7841\ : CEMux
    port map (
            O => \N__34004\,
            I => \N__33999\
        );

    \I__7840\ : CEMux
    port map (
            O => \N__34003\,
            I => \N__33993\
        );

    \I__7839\ : CEMux
    port map (
            O => \N__34002\,
            I => \N__33989\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__33999\,
            I => \N__33979\
        );

    \I__7837\ : CascadeMux
    port map (
            O => \N__33998\,
            I => \N__33974\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__33997\,
            I => \N__33971\
        );

    \I__7835\ : CEMux
    port map (
            O => \N__33996\,
            I => \N__33967\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__33993\,
            I => \N__33964\
        );

    \I__7833\ : CEMux
    port map (
            O => \N__33992\,
            I => \N__33961\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__33989\,
            I => \N__33958\
        );

    \I__7831\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33948\
        );

    \I__7830\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33948\
        );

    \I__7829\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33948\
        );

    \I__7828\ : CascadeMux
    port map (
            O => \N__33985\,
            I => \N__33945\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33937\
        );

    \I__7826\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33937\
        );

    \I__7825\ : InMux
    port map (
            O => \N__33982\,
            I => \N__33937\
        );

    \I__7824\ : Span4Mux_s2_v
    port map (
            O => \N__33979\,
            I => \N__33930\
        );

    \I__7823\ : InMux
    port map (
            O => \N__33978\,
            I => \N__33927\
        );

    \I__7822\ : InMux
    port map (
            O => \N__33977\,
            I => \N__33918\
        );

    \I__7821\ : InMux
    port map (
            O => \N__33974\,
            I => \N__33918\
        );

    \I__7820\ : InMux
    port map (
            O => \N__33971\,
            I => \N__33918\
        );

    \I__7819\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33918\
        );

    \I__7818\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33910\
        );

    \I__7817\ : Span4Mux_s1_h
    port map (
            O => \N__33964\,
            I => \N__33910\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33907\
        );

    \I__7815\ : Span4Mux_v
    port map (
            O => \N__33958\,
            I => \N__33904\
        );

    \I__7814\ : InMux
    port map (
            O => \N__33957\,
            I => \N__33899\
        );

    \I__7813\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33899\
        );

    \I__7812\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33896\
        );

    \I__7811\ : LocalMux
    port map (
            O => \N__33948\,
            I => \N__33893\
        );

    \I__7810\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33888\
        );

    \I__7809\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33888\
        );

    \I__7808\ : LocalMux
    port map (
            O => \N__33937\,
            I => \N__33885\
        );

    \I__7807\ : CEMux
    port map (
            O => \N__33936\,
            I => \N__33882\
        );

    \I__7806\ : CEMux
    port map (
            O => \N__33935\,
            I => \N__33879\
        );

    \I__7805\ : CEMux
    port map (
            O => \N__33934\,
            I => \N__33876\
        );

    \I__7804\ : CEMux
    port map (
            O => \N__33933\,
            I => \N__33873\
        );

    \I__7803\ : Span4Mux_s3_h
    port map (
            O => \N__33930\,
            I => \N__33870\
        );

    \I__7802\ : LocalMux
    port map (
            O => \N__33927\,
            I => \N__33865\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__33918\,
            I => \N__33865\
        );

    \I__7800\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33858\
        );

    \I__7799\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33858\
        );

    \I__7798\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33858\
        );

    \I__7797\ : Span4Mux_s2_v
    port map (
            O => \N__33910\,
            I => \N__33841\
        );

    \I__7796\ : Span4Mux_s2_v
    port map (
            O => \N__33907\,
            I => \N__33841\
        );

    \I__7795\ : Span4Mux_v
    port map (
            O => \N__33904\,
            I => \N__33841\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__33899\,
            I => \N__33841\
        );

    \I__7793\ : LocalMux
    port map (
            O => \N__33896\,
            I => \N__33841\
        );

    \I__7792\ : Span4Mux_h
    port map (
            O => \N__33893\,
            I => \N__33841\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__33888\,
            I => \N__33841\
        );

    \I__7790\ : Span4Mux_s2_v
    port map (
            O => \N__33885\,
            I => \N__33841\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__33882\,
            I => \POWERLED.count_clk_en\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__33879\,
            I => \POWERLED.count_clk_en\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__33876\,
            I => \POWERLED.count_clk_en\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__33873\,
            I => \POWERLED.count_clk_en\
        );

    \I__7785\ : Odrv4
    port map (
            O => \N__33870\,
            I => \POWERLED.count_clk_en\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__33865\,
            I => \POWERLED.count_clk_en\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__33858\,
            I => \POWERLED.count_clk_en\
        );

    \I__7782\ : Odrv4
    port map (
            O => \N__33841\,
            I => \POWERLED.count_clk_en\
        );

    \I__7781\ : CascadeMux
    port map (
            O => \N__33824\,
            I => \POWERLED.N_2341_i_cascade_\
        );

    \I__7780\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33812\
        );

    \I__7779\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33812\
        );

    \I__7778\ : InMux
    port map (
            O => \N__33819\,
            I => \N__33808\
        );

    \I__7777\ : InMux
    port map (
            O => \N__33818\,
            I => \N__33805\
        );

    \I__7776\ : InMux
    port map (
            O => \N__33817\,
            I => \N__33799\
        );

    \I__7775\ : LocalMux
    port map (
            O => \N__33812\,
            I => \N__33796\
        );

    \I__7774\ : InMux
    port map (
            O => \N__33811\,
            I => \N__33790\
        );

    \I__7773\ : LocalMux
    port map (
            O => \N__33808\,
            I => \N__33786\
        );

    \I__7772\ : LocalMux
    port map (
            O => \N__33805\,
            I => \N__33783\
        );

    \I__7771\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33780\
        );

    \I__7770\ : InMux
    port map (
            O => \N__33803\,
            I => \N__33777\
        );

    \I__7769\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33773\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__33799\,
            I => \N__33768\
        );

    \I__7767\ : Span4Mux_h
    port map (
            O => \N__33796\,
            I => \N__33768\
        );

    \I__7766\ : InMux
    port map (
            O => \N__33795\,
            I => \N__33765\
        );

    \I__7765\ : InMux
    port map (
            O => \N__33794\,
            I => \N__33762\
        );

    \I__7764\ : InMux
    port map (
            O => \N__33793\,
            I => \N__33759\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__33790\,
            I => \N__33756\
        );

    \I__7762\ : InMux
    port map (
            O => \N__33789\,
            I => \N__33753\
        );

    \I__7761\ : Span4Mux_s3_h
    port map (
            O => \N__33786\,
            I => \N__33748\
        );

    \I__7760\ : Span4Mux_v
    port map (
            O => \N__33783\,
            I => \N__33748\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33743\
        );

    \I__7758\ : LocalMux
    port map (
            O => \N__33777\,
            I => \N__33743\
        );

    \I__7757\ : InMux
    port map (
            O => \N__33776\,
            I => \N__33740\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__33773\,
            I => \N__33728\
        );

    \I__7755\ : Span4Mux_v
    port map (
            O => \N__33768\,
            I => \N__33728\
        );

    \I__7754\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33728\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33725\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__33759\,
            I => \N__33718\
        );

    \I__7751\ : Span4Mux_v
    port map (
            O => \N__33756\,
            I => \N__33718\
        );

    \I__7750\ : LocalMux
    port map (
            O => \N__33753\,
            I => \N__33718\
        );

    \I__7749\ : Span4Mux_v
    port map (
            O => \N__33748\,
            I => \N__33713\
        );

    \I__7748\ : Span4Mux_s3_h
    port map (
            O => \N__33743\,
            I => \N__33713\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__33740\,
            I => \N__33710\
        );

    \I__7746\ : InMux
    port map (
            O => \N__33739\,
            I => \N__33707\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33738\,
            I => \N__33704\
        );

    \I__7744\ : InMux
    port map (
            O => \N__33737\,
            I => \N__33697\
        );

    \I__7743\ : InMux
    port map (
            O => \N__33736\,
            I => \N__33697\
        );

    \I__7742\ : InMux
    port map (
            O => \N__33735\,
            I => \N__33697\
        );

    \I__7741\ : Span4Mux_v
    port map (
            O => \N__33728\,
            I => \N__33690\
        );

    \I__7740\ : Span4Mux_s0_h
    port map (
            O => \N__33725\,
            I => \N__33690\
        );

    \I__7739\ : Span4Mux_v
    port map (
            O => \N__33718\,
            I => \N__33690\
        );

    \I__7738\ : Odrv4
    port map (
            O => \N__33713\,
            I => \POWERLED.N_430\
        );

    \I__7737\ : Odrv4
    port map (
            O => \N__33710\,
            I => \POWERLED.N_430\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__33707\,
            I => \POWERLED.N_430\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__33704\,
            I => \POWERLED.N_430\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__33697\,
            I => \POWERLED.N_430\
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__33690\,
            I => \POWERLED.N_430\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__33677\,
            I => \POWERLED.N_529_cascade_\
        );

    \I__7731\ : CascadeMux
    port map (
            O => \N__33674\,
            I => \N__33663\
        );

    \I__7730\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33652\
        );

    \I__7729\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33652\
        );

    \I__7728\ : CascadeMux
    port map (
            O => \N__33671\,
            I => \N__33648\
        );

    \I__7727\ : CascadeMux
    port map (
            O => \N__33670\,
            I => \N__33645\
        );

    \I__7726\ : CascadeMux
    port map (
            O => \N__33669\,
            I => \N__33639\
        );

    \I__7725\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33636\
        );

    \I__7724\ : InMux
    port map (
            O => \N__33667\,
            I => \N__33631\
        );

    \I__7723\ : InMux
    port map (
            O => \N__33666\,
            I => \N__33628\
        );

    \I__7722\ : InMux
    port map (
            O => \N__33663\,
            I => \N__33625\
        );

    \I__7721\ : InMux
    port map (
            O => \N__33662\,
            I => \N__33622\
        );

    \I__7720\ : InMux
    port map (
            O => \N__33661\,
            I => \N__33618\
        );

    \I__7719\ : InMux
    port map (
            O => \N__33660\,
            I => \N__33615\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33659\,
            I => \N__33612\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33658\,
            I => \N__33607\
        );

    \I__7716\ : InMux
    port map (
            O => \N__33657\,
            I => \N__33607\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__33652\,
            I => \N__33604\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33595\
        );

    \I__7713\ : InMux
    port map (
            O => \N__33648\,
            I => \N__33595\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33645\,
            I => \N__33590\
        );

    \I__7711\ : InMux
    port map (
            O => \N__33644\,
            I => \N__33590\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__33643\,
            I => \N__33586\
        );

    \I__7709\ : CascadeMux
    port map (
            O => \N__33642\,
            I => \N__33583\
        );

    \I__7708\ : InMux
    port map (
            O => \N__33639\,
            I => \N__33579\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__33636\,
            I => \N__33576\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33571\
        );

    \I__7705\ : InMux
    port map (
            O => \N__33634\,
            I => \N__33571\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33566\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33566\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__33625\,
            I => \N__33561\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__33622\,
            I => \N__33561\
        );

    \I__7700\ : IoInMux
    port map (
            O => \N__33621\,
            I => \N__33558\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__33618\,
            I => \N__33555\
        );

    \I__7698\ : LocalMux
    port map (
            O => \N__33615\,
            I => \N__33548\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__33612\,
            I => \N__33548\
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33548\
        );

    \I__7695\ : Span4Mux_h
    port map (
            O => \N__33604\,
            I => \N__33545\
        );

    \I__7694\ : InMux
    port map (
            O => \N__33603\,
            I => \N__33540\
        );

    \I__7693\ : InMux
    port map (
            O => \N__33602\,
            I => \N__33533\
        );

    \I__7692\ : InMux
    port map (
            O => \N__33601\,
            I => \N__33533\
        );

    \I__7691\ : InMux
    port map (
            O => \N__33600\,
            I => \N__33533\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__33595\,
            I => \N__33528\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__33590\,
            I => \N__33528\
        );

    \I__7688\ : InMux
    port map (
            O => \N__33589\,
            I => \N__33523\
        );

    \I__7687\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33523\
        );

    \I__7686\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33518\
        );

    \I__7685\ : InMux
    port map (
            O => \N__33582\,
            I => \N__33518\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__33579\,
            I => \N__33515\
        );

    \I__7683\ : Span4Mux_v
    port map (
            O => \N__33576\,
            I => \N__33510\
        );

    \I__7682\ : LocalMux
    port map (
            O => \N__33571\,
            I => \N__33510\
        );

    \I__7681\ : Span4Mux_v
    port map (
            O => \N__33566\,
            I => \N__33505\
        );

    \I__7680\ : Span4Mux_s0_h
    port map (
            O => \N__33561\,
            I => \N__33505\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__33558\,
            I => \N__33502\
        );

    \I__7678\ : Span4Mux_v
    port map (
            O => \N__33555\,
            I => \N__33497\
        );

    \I__7677\ : Span4Mux_v
    port map (
            O => \N__33548\,
            I => \N__33497\
        );

    \I__7676\ : Span4Mux_v
    port map (
            O => \N__33545\,
            I => \N__33494\
        );

    \I__7675\ : InMux
    port map (
            O => \N__33544\,
            I => \N__33489\
        );

    \I__7674\ : InMux
    port map (
            O => \N__33543\,
            I => \N__33489\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__33540\,
            I => \N__33484\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__33533\,
            I => \N__33484\
        );

    \I__7671\ : Span12Mux_s5_h
    port map (
            O => \N__33528\,
            I => \N__33479\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__33523\,
            I => \N__33479\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__33518\,
            I => \N__33470\
        );

    \I__7668\ : Span4Mux_v
    port map (
            O => \N__33515\,
            I => \N__33470\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__33510\,
            I => \N__33470\
        );

    \I__7666\ : Span4Mux_h
    port map (
            O => \N__33505\,
            I => \N__33470\
        );

    \I__7665\ : Odrv12
    port map (
            O => \N__33502\,
            I => \G_141\
        );

    \I__7664\ : Odrv4
    port map (
            O => \N__33497\,
            I => \G_141\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__33494\,
            I => \G_141\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__33489\,
            I => \G_141\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__33484\,
            I => \G_141\
        );

    \I__7660\ : Odrv12
    port map (
            O => \N__33479\,
            I => \G_141\
        );

    \I__7659\ : Odrv4
    port map (
            O => \N__33470\,
            I => \G_141\
        );

    \I__7658\ : CascadeMux
    port map (
            O => \N__33455\,
            I => \N__33452\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33446\
        );

    \I__7656\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33446\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__33446\,
            I => \N__33443\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__33443\,
            I => \N__33440\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__33440\,
            I => \POWERLED.dutycycle_en_12\
        );

    \I__7652\ : InMux
    port map (
            O => \N__33437\,
            I => \N__33429\
        );

    \I__7651\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33426\
        );

    \I__7650\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33423\
        );

    \I__7649\ : InMux
    port map (
            O => \N__33434\,
            I => \N__33418\
        );

    \I__7648\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33418\
        );

    \I__7647\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33415\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__33429\,
            I => \N__33412\
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__33426\,
            I => \N__33409\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__33423\,
            I => \N__33404\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__33418\,
            I => \N__33404\
        );

    \I__7642\ : LocalMux
    port map (
            O => \N__33415\,
            I => \N__33397\
        );

    \I__7641\ : Span4Mux_h
    port map (
            O => \N__33412\,
            I => \N__33397\
        );

    \I__7640\ : Span4Mux_v
    port map (
            O => \N__33409\,
            I => \N__33394\
        );

    \I__7639\ : Span4Mux_v
    port map (
            O => \N__33404\,
            I => \N__33391\
        );

    \I__7638\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33386\
        );

    \I__7637\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33386\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__33397\,
            I => \POWERLED.func_state_RNILP0FZ0Z_1\
        );

    \I__7635\ : Odrv4
    port map (
            O => \N__33394\,
            I => \POWERLED.func_state_RNILP0FZ0Z_1\
        );

    \I__7634\ : Odrv4
    port map (
            O => \N__33391\,
            I => \POWERLED.func_state_RNILP0FZ0Z_1\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33386\,
            I => \POWERLED.func_state_RNILP0FZ0Z_1\
        );

    \I__7632\ : CascadeMux
    port map (
            O => \N__33377\,
            I => \N__33373\
        );

    \I__7631\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33355\
        );

    \I__7630\ : InMux
    port map (
            O => \N__33373\,
            I => \N__33350\
        );

    \I__7629\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33350\
        );

    \I__7628\ : CascadeMux
    port map (
            O => \N__33371\,
            I => \N__33346\
        );

    \I__7627\ : InMux
    port map (
            O => \N__33370\,
            I => \N__33342\
        );

    \I__7626\ : InMux
    port map (
            O => \N__33369\,
            I => \N__33339\
        );

    \I__7625\ : InMux
    port map (
            O => \N__33368\,
            I => \N__33330\
        );

    \I__7624\ : InMux
    port map (
            O => \N__33367\,
            I => \N__33330\
        );

    \I__7623\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33330\
        );

    \I__7622\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33330\
        );

    \I__7621\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33327\
        );

    \I__7620\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33318\
        );

    \I__7619\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33318\
        );

    \I__7618\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33318\
        );

    \I__7617\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33318\
        );

    \I__7616\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33313\
        );

    \I__7615\ : InMux
    port map (
            O => \N__33358\,
            I => \N__33313\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__33355\,
            I => \N__33308\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__33350\,
            I => \N__33308\
        );

    \I__7612\ : InMux
    port map (
            O => \N__33349\,
            I => \N__33303\
        );

    \I__7611\ : InMux
    port map (
            O => \N__33346\,
            I => \N__33303\
        );

    \I__7610\ : InMux
    port map (
            O => \N__33345\,
            I => \N__33284\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__33342\,
            I => \N__33281\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__33339\,
            I => \N__33273\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__33330\,
            I => \N__33273\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__33327\,
            I => \N__33273\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__33318\,
            I => \N__33268\
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__33313\,
            I => \N__33268\
        );

    \I__7603\ : Span4Mux_s2_h
    port map (
            O => \N__33308\,
            I => \N__33263\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__33303\,
            I => \N__33263\
        );

    \I__7601\ : InMux
    port map (
            O => \N__33302\,
            I => \N__33258\
        );

    \I__7600\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33258\
        );

    \I__7599\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33253\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33253\
        );

    \I__7597\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33248\
        );

    \I__7596\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33248\
        );

    \I__7595\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33243\
        );

    \I__7594\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33243\
        );

    \I__7593\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33236\
        );

    \I__7592\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33236\
        );

    \I__7591\ : InMux
    port map (
            O => \N__33292\,
            I => \N__33236\
        );

    \I__7590\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33231\
        );

    \I__7589\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33231\
        );

    \I__7588\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33228\
        );

    \I__7587\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33223\
        );

    \I__7586\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33223\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__33284\,
            I => \N__33218\
        );

    \I__7584\ : Span4Mux_v
    port map (
            O => \N__33281\,
            I => \N__33218\
        );

    \I__7583\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33215\
        );

    \I__7582\ : Span4Mux_v
    port map (
            O => \N__33273\,
            I => \N__33208\
        );

    \I__7581\ : Span4Mux_h
    port map (
            O => \N__33268\,
            I => \N__33208\
        );

    \I__7580\ : Span4Mux_v
    port map (
            O => \N__33263\,
            I => \N__33208\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__33258\,
            I => \N__33193\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__33253\,
            I => \N__33193\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__33248\,
            I => \N__33193\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__33243\,
            I => \N__33193\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__33236\,
            I => \N__33193\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33193\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__33228\,
            I => \N__33193\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__33223\,
            I => \POWERLED.func_state\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__33218\,
            I => \POWERLED.func_state\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__33215\,
            I => \POWERLED.func_state\
        );

    \I__7569\ : Odrv4
    port map (
            O => \N__33208\,
            I => \POWERLED.func_state\
        );

    \I__7568\ : Odrv12
    port map (
            O => \N__33193\,
            I => \POWERLED.func_state\
        );

    \I__7567\ : CascadeMux
    port map (
            O => \N__33182\,
            I => \N__33179\
        );

    \I__7566\ : InMux
    port map (
            O => \N__33179\,
            I => \N__33176\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__33176\,
            I => \POWERLED.N_527\
        );

    \I__7564\ : InMux
    port map (
            O => \N__33173\,
            I => \N__33170\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__33170\,
            I => \N__33166\
        );

    \I__7562\ : InMux
    port map (
            O => \N__33169\,
            I => \N__33163\
        );

    \I__7561\ : Span4Mux_v
    port map (
            O => \N__33166\,
            I => \N__33160\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__33163\,
            I => \N__33155\
        );

    \I__7559\ : Span4Mux_h
    port map (
            O => \N__33160\,
            I => \N__33155\
        );

    \I__7558\ : Odrv4
    port map (
            O => \N__33155\,
            I => \POWERLED.N_2341_i\
        );

    \I__7557\ : InMux
    port map (
            O => \N__33152\,
            I => \N__33149\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__33149\,
            I => \POWERLED.un1_clk_100khz_48_and_i_1\
        );

    \I__7555\ : CascadeMux
    port map (
            O => \N__33146\,
            I => \N__33138\
        );

    \I__7554\ : CascadeMux
    port map (
            O => \N__33145\,
            I => \N__33129\
        );

    \I__7553\ : InMux
    port map (
            O => \N__33144\,
            I => \N__33125\
        );

    \I__7552\ : InMux
    port map (
            O => \N__33143\,
            I => \N__33119\
        );

    \I__7551\ : InMux
    port map (
            O => \N__33142\,
            I => \N__33116\
        );

    \I__7550\ : InMux
    port map (
            O => \N__33141\,
            I => \N__33112\
        );

    \I__7549\ : InMux
    port map (
            O => \N__33138\,
            I => \N__33109\
        );

    \I__7548\ : InMux
    port map (
            O => \N__33137\,
            I => \N__33101\
        );

    \I__7547\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33101\
        );

    \I__7546\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33098\
        );

    \I__7545\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33095\
        );

    \I__7544\ : InMux
    port map (
            O => \N__33133\,
            I => \N__33090\
        );

    \I__7543\ : InMux
    port map (
            O => \N__33132\,
            I => \N__33090\
        );

    \I__7542\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33082\
        );

    \I__7541\ : InMux
    port map (
            O => \N__33128\,
            I => \N__33082\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__33125\,
            I => \N__33079\
        );

    \I__7539\ : InMux
    port map (
            O => \N__33124\,
            I => \N__33076\
        );

    \I__7538\ : InMux
    port map (
            O => \N__33123\,
            I => \N__33073\
        );

    \I__7537\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33070\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__33119\,
            I => \N__33065\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__33116\,
            I => \N__33065\
        );

    \I__7534\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33062\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__33112\,
            I => \N__33057\
        );

    \I__7532\ : LocalMux
    port map (
            O => \N__33109\,
            I => \N__33057\
        );

    \I__7531\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33053\
        );

    \I__7530\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33048\
        );

    \I__7529\ : InMux
    port map (
            O => \N__33106\,
            I => \N__33045\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__33101\,
            I => \N__33042\
        );

    \I__7527\ : LocalMux
    port map (
            O => \N__33098\,
            I => \N__33035\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__33095\,
            I => \N__33035\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__33090\,
            I => \N__33035\
        );

    \I__7524\ : InMux
    port map (
            O => \N__33089\,
            I => \N__33028\
        );

    \I__7523\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33028\
        );

    \I__7522\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33028\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__33082\,
            I => \N__33019\
        );

    \I__7520\ : Span4Mux_h
    port map (
            O => \N__33079\,
            I => \N__33019\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__33076\,
            I => \N__33019\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__33073\,
            I => \N__33019\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__33070\,
            I => \N__33016\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__33065\,
            I => \N__33013\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__33062\,
            I => \N__33008\
        );

    \I__7514\ : Span4Mux_v
    port map (
            O => \N__33057\,
            I => \N__33008\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__33056\,
            I => \N__33005\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__33053\,
            I => \N__33002\
        );

    \I__7511\ : InMux
    port map (
            O => \N__33052\,
            I => \N__32997\
        );

    \I__7510\ : InMux
    port map (
            O => \N__33051\,
            I => \N__32997\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__33048\,
            I => \N__32994\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__32985\
        );

    \I__7507\ : Span4Mux_v
    port map (
            O => \N__33042\,
            I => \N__32985\
        );

    \I__7506\ : Span4Mux_v
    port map (
            O => \N__33035\,
            I => \N__32985\
        );

    \I__7505\ : LocalMux
    port map (
            O => \N__33028\,
            I => \N__32985\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__33019\,
            I => \N__32976\
        );

    \I__7503\ : Span4Mux_v
    port map (
            O => \N__33016\,
            I => \N__32976\
        );

    \I__7502\ : Span4Mux_s0_h
    port map (
            O => \N__33013\,
            I => \N__32976\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__33008\,
            I => \N__32976\
        );

    \I__7500\ : InMux
    port map (
            O => \N__33005\,
            I => \N__32973\
        );

    \I__7499\ : Odrv4
    port map (
            O => \N__33002\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__32997\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7497\ : Odrv12
    port map (
            O => \N__32994\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__32985\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7495\ : Odrv4
    port map (
            O => \N__32976\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7494\ : LocalMux
    port map (
            O => \N__32973\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__7493\ : InMux
    port map (
            O => \N__32960\,
            I => \N__32954\
        );

    \I__7492\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32950\
        );

    \I__7491\ : CascadeMux
    port map (
            O => \N__32958\,
            I => \N__32947\
        );

    \I__7490\ : CascadeMux
    port map (
            O => \N__32957\,
            I => \N__32943\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32937\
        );

    \I__7488\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32934\
        );

    \I__7487\ : LocalMux
    port map (
            O => \N__32950\,
            I => \N__32931\
        );

    \I__7486\ : InMux
    port map (
            O => \N__32947\,
            I => \N__32926\
        );

    \I__7485\ : InMux
    port map (
            O => \N__32946\,
            I => \N__32926\
        );

    \I__7484\ : InMux
    port map (
            O => \N__32943\,
            I => \N__32921\
        );

    \I__7483\ : InMux
    port map (
            O => \N__32942\,
            I => \N__32921\
        );

    \I__7482\ : InMux
    port map (
            O => \N__32941\,
            I => \N__32916\
        );

    \I__7481\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32916\
        );

    \I__7480\ : Span12Mux_s5_v
    port map (
            O => \N__32937\,
            I => \N__32911\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__32934\,
            I => \N__32911\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__32931\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__32926\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__7476\ : LocalMux
    port map (
            O => \N__32921\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__32916\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__7474\ : Odrv12
    port map (
            O => \N__32911\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8\
        );

    \I__7473\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32897\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__32897\,
            I => \POWERLED.g0_i_0_0_0\
        );

    \I__7471\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32891\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__32891\,
            I => \N__32888\
        );

    \I__7469\ : Span4Mux_v
    port map (
            O => \N__32888\,
            I => \N__32885\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__32885\,
            I => \N__32882\
        );

    \I__7467\ : Span4Mux_h
    port map (
            O => \N__32882\,
            I => \N__32877\
        );

    \I__7466\ : InMux
    port map (
            O => \N__32881\,
            I => \N__32872\
        );

    \I__7465\ : InMux
    port map (
            O => \N__32880\,
            I => \N__32872\
        );

    \I__7464\ : Odrv4
    port map (
            O => \N__32877\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__32872\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__7462\ : IoInMux
    port map (
            O => \N__32867\,
            I => \N__32864\
        );

    \I__7461\ : LocalMux
    port map (
            O => \N__32864\,
            I => \N__32861\
        );

    \I__7460\ : Span4Mux_s0_h
    port map (
            O => \N__32861\,
            I => \N__32858\
        );

    \I__7459\ : Odrv4
    port map (
            O => \N__32858\,
            I => vpp_en
        );

    \I__7458\ : CascadeMux
    port map (
            O => \N__32855\,
            I => \N__32841\
        );

    \I__7457\ : CascadeMux
    port map (
            O => \N__32854\,
            I => \N__32838\
        );

    \I__7456\ : CascadeMux
    port map (
            O => \N__32853\,
            I => \N__32833\
        );

    \I__7455\ : InMux
    port map (
            O => \N__32852\,
            I => \N__32823\
        );

    \I__7454\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32823\
        );

    \I__7453\ : InMux
    port map (
            O => \N__32850\,
            I => \N__32823\
        );

    \I__7452\ : InMux
    port map (
            O => \N__32849\,
            I => \N__32818\
        );

    \I__7451\ : InMux
    port map (
            O => \N__32848\,
            I => \N__32815\
        );

    \I__7450\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32807\
        );

    \I__7449\ : InMux
    port map (
            O => \N__32846\,
            I => \N__32807\
        );

    \I__7448\ : InMux
    port map (
            O => \N__32845\,
            I => \N__32802\
        );

    \I__7447\ : InMux
    port map (
            O => \N__32844\,
            I => \N__32802\
        );

    \I__7446\ : InMux
    port map (
            O => \N__32841\,
            I => \N__32797\
        );

    \I__7445\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32797\
        );

    \I__7444\ : InMux
    port map (
            O => \N__32837\,
            I => \N__32790\
        );

    \I__7443\ : InMux
    port map (
            O => \N__32836\,
            I => \N__32790\
        );

    \I__7442\ : InMux
    port map (
            O => \N__32833\,
            I => \N__32790\
        );

    \I__7441\ : InMux
    port map (
            O => \N__32832\,
            I => \N__32783\
        );

    \I__7440\ : InMux
    port map (
            O => \N__32831\,
            I => \N__32783\
        );

    \I__7439\ : InMux
    port map (
            O => \N__32830\,
            I => \N__32783\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__32823\,
            I => \N__32780\
        );

    \I__7437\ : CascadeMux
    port map (
            O => \N__32822\,
            I => \N__32777\
        );

    \I__7436\ : CascadeMux
    port map (
            O => \N__32821\,
            I => \N__32774\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__32818\,
            I => \N__32766\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32763\
        );

    \I__7433\ : InMux
    port map (
            O => \N__32814\,
            I => \N__32760\
        );

    \I__7432\ : InMux
    port map (
            O => \N__32813\,
            I => \N__32757\
        );

    \I__7431\ : InMux
    port map (
            O => \N__32812\,
            I => \N__32754\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32751\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__32802\,
            I => \N__32742\
        );

    \I__7428\ : LocalMux
    port map (
            O => \N__32797\,
            I => \N__32742\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32742\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__32783\,
            I => \N__32742\
        );

    \I__7425\ : Span4Mux_h
    port map (
            O => \N__32780\,
            I => \N__32739\
        );

    \I__7424\ : InMux
    port map (
            O => \N__32777\,
            I => \N__32736\
        );

    \I__7423\ : InMux
    port map (
            O => \N__32774\,
            I => \N__32731\
        );

    \I__7422\ : InMux
    port map (
            O => \N__32773\,
            I => \N__32731\
        );

    \I__7421\ : InMux
    port map (
            O => \N__32772\,
            I => \N__32728\
        );

    \I__7420\ : InMux
    port map (
            O => \N__32771\,
            I => \N__32721\
        );

    \I__7419\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32721\
        );

    \I__7418\ : InMux
    port map (
            O => \N__32769\,
            I => \N__32721\
        );

    \I__7417\ : Span4Mux_h
    port map (
            O => \N__32766\,
            I => \N__32710\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__32763\,
            I => \N__32710\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__32760\,
            I => \N__32710\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__32757\,
            I => \N__32710\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__32754\,
            I => \N__32710\
        );

    \I__7412\ : Span4Mux_h
    port map (
            O => \N__32751\,
            I => \N__32701\
        );

    \I__7411\ : Span4Mux_v
    port map (
            O => \N__32742\,
            I => \N__32701\
        );

    \I__7410\ : Span4Mux_v
    port map (
            O => \N__32739\,
            I => \N__32701\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__32736\,
            I => \N__32701\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__32731\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__32728\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__32721\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__32710\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__32701\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7403\ : InMux
    port map (
            O => \N__32690\,
            I => \N__32687\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__32687\,
            I => \N__32684\
        );

    \I__7401\ : Odrv12
    port map (
            O => \N__32684\,
            I => \POWERLED.G_7_i_o5_0\
        );

    \I__7400\ : CascadeMux
    port map (
            O => \N__32681\,
            I => \N__32677\
        );

    \I__7399\ : CascadeMux
    port map (
            O => \N__32680\,
            I => \N__32671\
        );

    \I__7398\ : InMux
    port map (
            O => \N__32677\,
            I => \N__32659\
        );

    \I__7397\ : InMux
    port map (
            O => \N__32676\,
            I => \N__32659\
        );

    \I__7396\ : InMux
    port map (
            O => \N__32675\,
            I => \N__32659\
        );

    \I__7395\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32659\
        );

    \I__7394\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32638\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32670\,
            I => \N__32638\
        );

    \I__7392\ : InMux
    port map (
            O => \N__32669\,
            I => \N__32638\
        );

    \I__7391\ : InMux
    port map (
            O => \N__32668\,
            I => \N__32635\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__32659\,
            I => \N__32630\
        );

    \I__7389\ : InMux
    port map (
            O => \N__32658\,
            I => \N__32625\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32625\
        );

    \I__7387\ : InMux
    port map (
            O => \N__32656\,
            I => \N__32622\
        );

    \I__7386\ : InMux
    port map (
            O => \N__32655\,
            I => \N__32615\
        );

    \I__7385\ : InMux
    port map (
            O => \N__32654\,
            I => \N__32615\
        );

    \I__7384\ : InMux
    port map (
            O => \N__32653\,
            I => \N__32615\
        );

    \I__7383\ : InMux
    port map (
            O => \N__32652\,
            I => \N__32612\
        );

    \I__7382\ : InMux
    port map (
            O => \N__32651\,
            I => \N__32609\
        );

    \I__7381\ : InMux
    port map (
            O => \N__32650\,
            I => \N__32602\
        );

    \I__7380\ : InMux
    port map (
            O => \N__32649\,
            I => \N__32602\
        );

    \I__7379\ : InMux
    port map (
            O => \N__32648\,
            I => \N__32602\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__32647\,
            I => \N__32599\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__32646\,
            I => \N__32595\
        );

    \I__7376\ : InMux
    port map (
            O => \N__32645\,
            I => \N__32592\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32585\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__32635\,
            I => \N__32585\
        );

    \I__7373\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32580\
        );

    \I__7372\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32580\
        );

    \I__7371\ : Span4Mux_s2_v
    port map (
            O => \N__32630\,
            I => \N__32573\
        );

    \I__7370\ : LocalMux
    port map (
            O => \N__32625\,
            I => \N__32573\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__32622\,
            I => \N__32570\
        );

    \I__7368\ : LocalMux
    port map (
            O => \N__32615\,
            I => \N__32567\
        );

    \I__7367\ : LocalMux
    port map (
            O => \N__32612\,
            I => \N__32560\
        );

    \I__7366\ : LocalMux
    port map (
            O => \N__32609\,
            I => \N__32560\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__32602\,
            I => \N__32560\
        );

    \I__7364\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32557\
        );

    \I__7363\ : InMux
    port map (
            O => \N__32598\,
            I => \N__32554\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32551\
        );

    \I__7361\ : LocalMux
    port map (
            O => \N__32592\,
            I => \N__32548\
        );

    \I__7360\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32545\
        );

    \I__7359\ : CascadeMux
    port map (
            O => \N__32590\,
            I => \N__32542\
        );

    \I__7358\ : Span4Mux_v
    port map (
            O => \N__32585\,
            I => \N__32535\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__32580\,
            I => \N__32535\
        );

    \I__7356\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32530\
        );

    \I__7355\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32530\
        );

    \I__7354\ : Span4Mux_v
    port map (
            O => \N__32573\,
            I => \N__32525\
        );

    \I__7353\ : Span4Mux_v
    port map (
            O => \N__32570\,
            I => \N__32518\
        );

    \I__7352\ : Span4Mux_h
    port map (
            O => \N__32567\,
            I => \N__32518\
        );

    \I__7351\ : Span4Mux_v
    port map (
            O => \N__32560\,
            I => \N__32513\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__32557\,
            I => \N__32513\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__32554\,
            I => \N__32510\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__32551\,
            I => \N__32503\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__32548\,
            I => \N__32503\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__32545\,
            I => \N__32503\
        );

    \I__7345\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32500\
        );

    \I__7344\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32497\
        );

    \I__7343\ : InMux
    port map (
            O => \N__32540\,
            I => \N__32494\
        );

    \I__7342\ : Span4Mux_h
    port map (
            O => \N__32535\,
            I => \N__32491\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__32530\,
            I => \N__32488\
        );

    \I__7340\ : InMux
    port map (
            O => \N__32529\,
            I => \N__32485\
        );

    \I__7339\ : InMux
    port map (
            O => \N__32528\,
            I => \N__32480\
        );

    \I__7338\ : Span4Mux_v
    port map (
            O => \N__32525\,
            I => \N__32477\
        );

    \I__7337\ : InMux
    port map (
            O => \N__32524\,
            I => \N__32472\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32523\,
            I => \N__32472\
        );

    \I__7335\ : Span4Mux_v
    port map (
            O => \N__32518\,
            I => \N__32457\
        );

    \I__7334\ : Span4Mux_h
    port map (
            O => \N__32513\,
            I => \N__32457\
        );

    \I__7333\ : Span4Mux_v
    port map (
            O => \N__32510\,
            I => \N__32457\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__32503\,
            I => \N__32457\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__32500\,
            I => \N__32457\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32497\,
            I => \N__32457\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32494\,
            I => \N__32457\
        );

    \I__7328\ : Span4Mux_v
    port map (
            O => \N__32491\,
            I => \N__32450\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__32488\,
            I => \N__32450\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__32485\,
            I => \N__32450\
        );

    \I__7325\ : InMux
    port map (
            O => \N__32484\,
            I => \N__32445\
        );

    \I__7324\ : InMux
    port map (
            O => \N__32483\,
            I => \N__32445\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__32480\,
            I => \N__32442\
        );

    \I__7322\ : Sp12to4
    port map (
            O => \N__32477\,
            I => \N__32437\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__32472\,
            I => \N__32437\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__32457\,
            I => \N__32434\
        );

    \I__7319\ : Span4Mux_h
    port map (
            O => \N__32450\,
            I => \N__32431\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__32445\,
            I => \N__32428\
        );

    \I__7317\ : Span12Mux_s8_h
    port map (
            O => \N__32442\,
            I => \N__32425\
        );

    \I__7316\ : Span12Mux_s8_h
    port map (
            O => \N__32437\,
            I => \N__32420\
        );

    \I__7315\ : Sp12to4
    port map (
            O => \N__32434\,
            I => \N__32420\
        );

    \I__7314\ : Span4Mux_v
    port map (
            O => \N__32431\,
            I => \N__32415\
        );

    \I__7313\ : Span4Mux_h
    port map (
            O => \N__32428\,
            I => \N__32415\
        );

    \I__7312\ : Odrv12
    port map (
            O => \N__32425\,
            I => slp_s4n
        );

    \I__7311\ : Odrv12
    port map (
            O => \N__32420\,
            I => slp_s4n
        );

    \I__7310\ : Odrv4
    port map (
            O => \N__32415\,
            I => slp_s4n
        );

    \I__7309\ : InMux
    port map (
            O => \N__32408\,
            I => \N__32403\
        );

    \I__7308\ : CascadeMux
    port map (
            O => \N__32407\,
            I => \N__32399\
        );

    \I__7307\ : CascadeMux
    port map (
            O => \N__32406\,
            I => \N__32396\
        );

    \I__7306\ : LocalMux
    port map (
            O => \N__32403\,
            I => \N__32391\
        );

    \I__7305\ : CascadeMux
    port map (
            O => \N__32402\,
            I => \N__32388\
        );

    \I__7304\ : InMux
    port map (
            O => \N__32399\,
            I => \N__32381\
        );

    \I__7303\ : InMux
    port map (
            O => \N__32396\,
            I => \N__32378\
        );

    \I__7302\ : InMux
    port map (
            O => \N__32395\,
            I => \N__32372\
        );

    \I__7301\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32369\
        );

    \I__7300\ : Span4Mux_v
    port map (
            O => \N__32391\,
            I => \N__32366\
        );

    \I__7299\ : InMux
    port map (
            O => \N__32388\,
            I => \N__32361\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32361\
        );

    \I__7297\ : InMux
    port map (
            O => \N__32386\,
            I => \N__32356\
        );

    \I__7296\ : InMux
    port map (
            O => \N__32385\,
            I => \N__32356\
        );

    \I__7295\ : CascadeMux
    port map (
            O => \N__32384\,
            I => \N__32353\
        );

    \I__7294\ : LocalMux
    port map (
            O => \N__32381\,
            I => \N__32347\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__32378\,
            I => \N__32347\
        );

    \I__7292\ : InMux
    port map (
            O => \N__32377\,
            I => \N__32344\
        );

    \I__7291\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32341\
        );

    \I__7290\ : InMux
    port map (
            O => \N__32375\,
            I => \N__32338\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__32372\,
            I => \N__32333\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32333\
        );

    \I__7287\ : Span4Mux_h
    port map (
            O => \N__32366\,
            I => \N__32328\
        );

    \I__7286\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32328\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__32356\,
            I => \N__32325\
        );

    \I__7284\ : InMux
    port map (
            O => \N__32353\,
            I => \N__32322\
        );

    \I__7283\ : InMux
    port map (
            O => \N__32352\,
            I => \N__32319\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__32347\,
            I => \N__32312\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__32344\,
            I => \N__32312\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__32341\,
            I => \N__32312\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__32338\,
            I => \N__32309\
        );

    \I__7278\ : Span4Mux_s3_v
    port map (
            O => \N__32333\,
            I => \N__32302\
        );

    \I__7277\ : Span4Mux_v
    port map (
            O => \N__32328\,
            I => \N__32302\
        );

    \I__7276\ : Span12Mux_v
    port map (
            O => \N__32325\,
            I => \N__32295\
        );

    \I__7275\ : LocalMux
    port map (
            O => \N__32322\,
            I => \N__32295\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__32319\,
            I => \N__32295\
        );

    \I__7273\ : Span4Mux_v
    port map (
            O => \N__32312\,
            I => \N__32290\
        );

    \I__7272\ : Span4Mux_v
    port map (
            O => \N__32309\,
            I => \N__32290\
        );

    \I__7271\ : InMux
    port map (
            O => \N__32308\,
            I => \N__32285\
        );

    \I__7270\ : InMux
    port map (
            O => \N__32307\,
            I => \N__32285\
        );

    \I__7269\ : Odrv4
    port map (
            O => \N__32302\,
            I => gpio_fpga_soc_4
        );

    \I__7268\ : Odrv12
    port map (
            O => \N__32295\,
            I => gpio_fpga_soc_4
        );

    \I__7267\ : Odrv4
    port map (
            O => \N__32290\,
            I => gpio_fpga_soc_4
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__32285\,
            I => gpio_fpga_soc_4
        );

    \I__7265\ : InMux
    port map (
            O => \N__32276\,
            I => \N__32267\
        );

    \I__7264\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32262\
        );

    \I__7263\ : InMux
    port map (
            O => \N__32274\,
            I => \N__32262\
        );

    \I__7262\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32259\
        );

    \I__7261\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32254\
        );

    \I__7260\ : CascadeMux
    port map (
            O => \N__32271\,
            I => \N__32251\
        );

    \I__7259\ : InMux
    port map (
            O => \N__32270\,
            I => \N__32245\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__32267\,
            I => \N__32241\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32238\
        );

    \I__7256\ : LocalMux
    port map (
            O => \N__32259\,
            I => \N__32234\
        );

    \I__7255\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32231\
        );

    \I__7254\ : InMux
    port map (
            O => \N__32257\,
            I => \N__32225\
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__32254\,
            I => \N__32222\
        );

    \I__7252\ : InMux
    port map (
            O => \N__32251\,
            I => \N__32219\
        );

    \I__7251\ : InMux
    port map (
            O => \N__32250\,
            I => \N__32216\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__32249\,
            I => \N__32212\
        );

    \I__7249\ : CascadeMux
    port map (
            O => \N__32248\,
            I => \N__32209\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__32245\,
            I => \N__32205\
        );

    \I__7247\ : InMux
    port map (
            O => \N__32244\,
            I => \N__32202\
        );

    \I__7246\ : Span4Mux_v
    port map (
            O => \N__32241\,
            I => \N__32197\
        );

    \I__7245\ : Span4Mux_v
    port map (
            O => \N__32238\,
            I => \N__32197\
        );

    \I__7244\ : CascadeMux
    port map (
            O => \N__32237\,
            I => \N__32194\
        );

    \I__7243\ : Span4Mux_v
    port map (
            O => \N__32234\,
            I => \N__32187\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__32231\,
            I => \N__32187\
        );

    \I__7241\ : InMux
    port map (
            O => \N__32230\,
            I => \N__32182\
        );

    \I__7240\ : InMux
    port map (
            O => \N__32229\,
            I => \N__32182\
        );

    \I__7239\ : InMux
    port map (
            O => \N__32228\,
            I => \N__32179\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__32225\,
            I => \N__32172\
        );

    \I__7237\ : Span4Mux_h
    port map (
            O => \N__32222\,
            I => \N__32172\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__32219\,
            I => \N__32172\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__32216\,
            I => \N__32169\
        );

    \I__7234\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32164\
        );

    \I__7233\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32164\
        );

    \I__7232\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32159\
        );

    \I__7231\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32159\
        );

    \I__7230\ : Span4Mux_v
    port map (
            O => \N__32205\,
            I => \N__32156\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__32202\,
            I => \N__32153\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__32197\,
            I => \N__32150\
        );

    \I__7227\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32147\
        );

    \I__7226\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32144\
        );

    \I__7225\ : InMux
    port map (
            O => \N__32192\,
            I => \N__32141\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__32187\,
            I => \N__32132\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__32182\,
            I => \N__32132\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__32179\,
            I => \N__32132\
        );

    \I__7221\ : Span4Mux_h
    port map (
            O => \N__32172\,
            I => \N__32132\
        );

    \I__7220\ : Span4Mux_v
    port map (
            O => \N__32169\,
            I => \N__32129\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32120\
        );

    \I__7218\ : LocalMux
    port map (
            O => \N__32159\,
            I => \N__32120\
        );

    \I__7217\ : Span4Mux_h
    port map (
            O => \N__32156\,
            I => \N__32120\
        );

    \I__7216\ : Span4Mux_s0_h
    port map (
            O => \N__32153\,
            I => \N__32120\
        );

    \I__7215\ : Odrv4
    port map (
            O => \N__32150\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__32147\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__32144\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7212\ : LocalMux
    port map (
            O => \N__32141\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7211\ : Odrv4
    port map (
            O => \N__32132\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7210\ : Odrv4
    port map (
            O => \N__32129\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7209\ : Odrv4
    port map (
            O => \N__32120\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__7208\ : InMux
    port map (
            O => \N__32105\,
            I => \N__32102\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__32102\,
            I => \N__32099\
        );

    \I__7206\ : Sp12to4
    port map (
            O => \N__32099\,
            I => \N__32096\
        );

    \I__7205\ : Odrv12
    port map (
            O => \N__32096\,
            I => \POWERLED.dutycycle_e_N_3L4_1\
        );

    \I__7204\ : CascadeMux
    port map (
            O => \N__32093\,
            I => \N__32089\
        );

    \I__7203\ : CascadeMux
    port map (
            O => \N__32092\,
            I => \N__32086\
        );

    \I__7202\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32076\
        );

    \I__7201\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32076\
        );

    \I__7200\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32071\
        );

    \I__7199\ : InMux
    port map (
            O => \N__32084\,
            I => \N__32071\
        );

    \I__7198\ : InMux
    port map (
            O => \N__32083\,
            I => \N__32068\
        );

    \I__7197\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32065\
        );

    \I__7196\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32059\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__32076\,
            I => \N__32052\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32071\,
            I => \N__32052\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__32068\,
            I => \N__32052\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__32065\,
            I => \N__32049\
        );

    \I__7191\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32046\
        );

    \I__7190\ : InMux
    port map (
            O => \N__32063\,
            I => \N__32041\
        );

    \I__7189\ : InMux
    port map (
            O => \N__32062\,
            I => \N__32041\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__32059\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__32052\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__7186\ : Odrv4
    port map (
            O => \N__32049\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__32046\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__32041\,
            I => \POWERLED.func_state_RNI_8Z0Z_1\
        );

    \I__7183\ : InMux
    port map (
            O => \N__32030\,
            I => \N__32027\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__32027\,
            I => \N__32022\
        );

    \I__7181\ : CascadeMux
    port map (
            O => \N__32026\,
            I => \N__32018\
        );

    \I__7180\ : CascadeMux
    port map (
            O => \N__32025\,
            I => \N__32015\
        );

    \I__7179\ : Span4Mux_s1_v
    port map (
            O => \N__32022\,
            I => \N__32009\
        );

    \I__7178\ : InMux
    port map (
            O => \N__32021\,
            I => \N__32004\
        );

    \I__7177\ : InMux
    port map (
            O => \N__32018\,
            I => \N__31998\
        );

    \I__7176\ : InMux
    port map (
            O => \N__32015\,
            I => \N__31998\
        );

    \I__7175\ : InMux
    port map (
            O => \N__32014\,
            I => \N__31991\
        );

    \I__7174\ : InMux
    port map (
            O => \N__32013\,
            I => \N__31991\
        );

    \I__7173\ : InMux
    port map (
            O => \N__32012\,
            I => \N__31988\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__32009\,
            I => \N__31984\
        );

    \I__7171\ : InMux
    port map (
            O => \N__32008\,
            I => \N__31979\
        );

    \I__7170\ : InMux
    port map (
            O => \N__32007\,
            I => \N__31979\
        );

    \I__7169\ : LocalMux
    port map (
            O => \N__32004\,
            I => \N__31976\
        );

    \I__7168\ : InMux
    port map (
            O => \N__32003\,
            I => \N__31973\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31970\
        );

    \I__7166\ : InMux
    port map (
            O => \N__31997\,
            I => \N__31967\
        );

    \I__7165\ : InMux
    port map (
            O => \N__31996\,
            I => \N__31964\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__31991\,
            I => \N__31959\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__31988\,
            I => \N__31959\
        );

    \I__7162\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31956\
        );

    \I__7161\ : Sp12to4
    port map (
            O => \N__31984\,
            I => \N__31950\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31947\
        );

    \I__7159\ : Span4Mux_v
    port map (
            O => \N__31976\,
            I => \N__31944\
        );

    \I__7158\ : LocalMux
    port map (
            O => \N__31973\,
            I => \N__31941\
        );

    \I__7157\ : Span4Mux_v
    port map (
            O => \N__31970\,
            I => \N__31932\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__31967\,
            I => \N__31932\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__31964\,
            I => \N__31932\
        );

    \I__7154\ : Span4Mux_v
    port map (
            O => \N__31959\,
            I => \N__31932\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__31956\,
            I => \N__31929\
        );

    \I__7152\ : InMux
    port map (
            O => \N__31955\,
            I => \N__31924\
        );

    \I__7151\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31924\
        );

    \I__7150\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31921\
        );

    \I__7149\ : Span12Mux_s8_h
    port map (
            O => \N__31950\,
            I => \N__31916\
        );

    \I__7148\ : Span12Mux_s3_h
    port map (
            O => \N__31947\,
            I => \N__31916\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__31944\,
            I => \N__31913\
        );

    \I__7146\ : Span4Mux_s1_v
    port map (
            O => \N__31941\,
            I => \N__31910\
        );

    \I__7145\ : Span4Mux_v
    port map (
            O => \N__31932\,
            I => \N__31903\
        );

    \I__7144\ : Span4Mux_s0_h
    port map (
            O => \N__31929\,
            I => \N__31903\
        );

    \I__7143\ : LocalMux
    port map (
            O => \N__31924\,
            I => \N__31903\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__31921\,
            I => \VCCST_EN_i_1\
        );

    \I__7141\ : Odrv12
    port map (
            O => \N__31916\,
            I => \VCCST_EN_i_1\
        );

    \I__7140\ : Odrv4
    port map (
            O => \N__31913\,
            I => \VCCST_EN_i_1\
        );

    \I__7139\ : Odrv4
    port map (
            O => \N__31910\,
            I => \VCCST_EN_i_1\
        );

    \I__7138\ : Odrv4
    port map (
            O => \N__31903\,
            I => \VCCST_EN_i_1\
        );

    \I__7137\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31888\
        );

    \I__7136\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31881\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31878\
        );

    \I__7134\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31875\
        );

    \I__7133\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31870\
        );

    \I__7132\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31870\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__31884\,
            I => \N__31865\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__31881\,
            I => \N__31861\
        );

    \I__7129\ : Span4Mux_v
    port map (
            O => \N__31878\,
            I => \N__31856\
        );

    \I__7128\ : LocalMux
    port map (
            O => \N__31875\,
            I => \N__31856\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__31870\,
            I => \N__31853\
        );

    \I__7126\ : InMux
    port map (
            O => \N__31869\,
            I => \N__31848\
        );

    \I__7125\ : InMux
    port map (
            O => \N__31868\,
            I => \N__31848\
        );

    \I__7124\ : InMux
    port map (
            O => \N__31865\,
            I => \N__31845\
        );

    \I__7123\ : InMux
    port map (
            O => \N__31864\,
            I => \N__31842\
        );

    \I__7122\ : Span4Mux_s1_h
    port map (
            O => \N__31861\,
            I => \N__31837\
        );

    \I__7121\ : Span4Mux_h
    port map (
            O => \N__31856\,
            I => \N__31837\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__31853\,
            I => \POWERLED.N_203\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__31848\,
            I => \POWERLED.N_203\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__31845\,
            I => \POWERLED.N_203\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__31842\,
            I => \POWERLED.N_203\
        );

    \I__7116\ : Odrv4
    port map (
            O => \N__31837\,
            I => \POWERLED.N_203\
        );

    \I__7115\ : CascadeMux
    port map (
            O => \N__31826\,
            I => \N__31817\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__31825\,
            I => \N__31814\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31824\,
            I => \N__31804\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31823\,
            I => \N__31799\
        );

    \I__7111\ : InMux
    port map (
            O => \N__31822\,
            I => \N__31799\
        );

    \I__7110\ : InMux
    port map (
            O => \N__31821\,
            I => \N__31789\
        );

    \I__7109\ : InMux
    port map (
            O => \N__31820\,
            I => \N__31789\
        );

    \I__7108\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31789\
        );

    \I__7107\ : InMux
    port map (
            O => \N__31814\,
            I => \N__31786\
        );

    \I__7106\ : InMux
    port map (
            O => \N__31813\,
            I => \N__31781\
        );

    \I__7105\ : InMux
    port map (
            O => \N__31812\,
            I => \N__31781\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31811\,
            I => \N__31778\
        );

    \I__7103\ : CascadeMux
    port map (
            O => \N__31810\,
            I => \N__31775\
        );

    \I__7102\ : CascadeMux
    port map (
            O => \N__31809\,
            I => \N__31770\
        );

    \I__7101\ : InMux
    port map (
            O => \N__31808\,
            I => \N__31766\
        );

    \I__7100\ : CascadeMux
    port map (
            O => \N__31807\,
            I => \N__31763\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__31804\,
            I => \N__31760\
        );

    \I__7098\ : LocalMux
    port map (
            O => \N__31799\,
            I => \N__31757\
        );

    \I__7097\ : CascadeMux
    port map (
            O => \N__31798\,
            I => \N__31753\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__31797\,
            I => \N__31747\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__31796\,
            I => \N__31743\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__31789\,
            I => \N__31739\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__31786\,
            I => \N__31736\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__31781\,
            I => \N__31733\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__31778\,
            I => \N__31730\
        );

    \I__7090\ : InMux
    port map (
            O => \N__31775\,
            I => \N__31723\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31774\,
            I => \N__31723\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31723\
        );

    \I__7087\ : InMux
    port map (
            O => \N__31770\,
            I => \N__31718\
        );

    \I__7086\ : InMux
    port map (
            O => \N__31769\,
            I => \N__31718\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31715\
        );

    \I__7084\ : InMux
    port map (
            O => \N__31763\,
            I => \N__31712\
        );

    \I__7083\ : Span4Mux_s2_h
    port map (
            O => \N__31760\,
            I => \N__31709\
        );

    \I__7082\ : Span12Mux_s5_v
    port map (
            O => \N__31757\,
            I => \N__31706\
        );

    \I__7081\ : InMux
    port map (
            O => \N__31756\,
            I => \N__31701\
        );

    \I__7080\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31701\
        );

    \I__7079\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31692\
        );

    \I__7078\ : InMux
    port map (
            O => \N__31751\,
            I => \N__31692\
        );

    \I__7077\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31692\
        );

    \I__7076\ : InMux
    port map (
            O => \N__31747\,
            I => \N__31692\
        );

    \I__7075\ : InMux
    port map (
            O => \N__31746\,
            I => \N__31685\
        );

    \I__7074\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31685\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31742\,
            I => \N__31685\
        );

    \I__7072\ : Span4Mux_v
    port map (
            O => \N__31739\,
            I => \N__31682\
        );

    \I__7071\ : Span4Mux_s2_h
    port map (
            O => \N__31736\,
            I => \N__31679\
        );

    \I__7070\ : Span12Mux_v
    port map (
            O => \N__31733\,
            I => \N__31676\
        );

    \I__7069\ : Span4Mux_v
    port map (
            O => \N__31730\,
            I => \N__31665\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31665\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__31718\,
            I => \N__31665\
        );

    \I__7066\ : Span4Mux_s3_h
    port map (
            O => \N__31715\,
            I => \N__31665\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__31712\,
            I => \N__31665\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__31709\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7063\ : Odrv12
    port map (
            O => \N__31706\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__31701\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7061\ : LocalMux
    port map (
            O => \N__31692\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7060\ : LocalMux
    port map (
            O => \N__31685\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7059\ : Odrv4
    port map (
            O => \N__31682\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7058\ : Odrv4
    port map (
            O => \N__31679\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7057\ : Odrv12
    port map (
            O => \N__31676\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7056\ : Odrv4
    port map (
            O => \N__31665\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__7055\ : CascadeMux
    port map (
            O => \N__31646\,
            I => \N__31643\
        );

    \I__7054\ : InMux
    port map (
            O => \N__31643\,
            I => \N__31640\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__31640\,
            I => \N__31637\
        );

    \I__7052\ : Span4Mux_v
    port map (
            O => \N__31637\,
            I => \N__31634\
        );

    \I__7051\ : Odrv4
    port map (
            O => \N__31634\,
            I => \POWERLED.N_505\
        );

    \I__7050\ : CascadeMux
    port map (
            O => \N__31631\,
            I => \POWERLED.dutycycleZ0Z_8_cascade_\
        );

    \I__7049\ : InMux
    port map (
            O => \N__31628\,
            I => \N__31622\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31627\,
            I => \N__31622\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__31622\,
            I => \POWERLED.dutycycle_RNIHDMC5Z0Z_3\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31619\,
            I => \N__31615\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31612\
        );

    \I__7044\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31607\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__31612\,
            I => \N__31607\
        );

    \I__7042\ : Span4Mux_s2_h
    port map (
            O => \N__31607\,
            I => \N__31604\
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__31604\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__7040\ : CascadeMux
    port map (
            O => \N__31601\,
            I => \N__31597\
        );

    \I__7039\ : InMux
    port map (
            O => \N__31600\,
            I => \N__31592\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31597\,
            I => \N__31592\
        );

    \I__7037\ : LocalMux
    port map (
            O => \N__31592\,
            I => \POWERLED.dutycycleZ1Z_3\
        );

    \I__7036\ : SRMux
    port map (
            O => \N__31589\,
            I => \N__31586\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__31586\,
            I => \N__31582\
        );

    \I__7034\ : SRMux
    port map (
            O => \N__31585\,
            I => \N__31577\
        );

    \I__7033\ : Span4Mux_h
    port map (
            O => \N__31582\,
            I => \N__31574\
        );

    \I__7032\ : SRMux
    port map (
            O => \N__31581\,
            I => \N__31571\
        );

    \I__7031\ : SRMux
    port map (
            O => \N__31580\,
            I => \N__31564\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__31577\,
            I => \N__31560\
        );

    \I__7029\ : IoSpan4Mux
    port map (
            O => \N__31574\,
            I => \N__31557\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__31571\,
            I => \N__31553\
        );

    \I__7027\ : SRMux
    port map (
            O => \N__31570\,
            I => \N__31550\
        );

    \I__7026\ : SRMux
    port map (
            O => \N__31569\,
            I => \N__31547\
        );

    \I__7025\ : SRMux
    port map (
            O => \N__31568\,
            I => \N__31544\
        );

    \I__7024\ : SRMux
    port map (
            O => \N__31567\,
            I => \N__31540\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__31564\,
            I => \N__31535\
        );

    \I__7022\ : SRMux
    port map (
            O => \N__31563\,
            I => \N__31532\
        );

    \I__7021\ : Span4Mux_h
    port map (
            O => \N__31560\,
            I => \N__31529\
        );

    \I__7020\ : IoSpan4Mux
    port map (
            O => \N__31557\,
            I => \N__31526\
        );

    \I__7019\ : SRMux
    port map (
            O => \N__31556\,
            I => \N__31523\
        );

    \I__7018\ : Span4Mux_s3_h
    port map (
            O => \N__31553\,
            I => \N__31514\
        );

    \I__7017\ : LocalMux
    port map (
            O => \N__31550\,
            I => \N__31514\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__31547\,
            I => \N__31514\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31514\
        );

    \I__7014\ : SRMux
    port map (
            O => \N__31543\,
            I => \N__31511\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__31540\,
            I => \N__31508\
        );

    \I__7012\ : SRMux
    port map (
            O => \N__31539\,
            I => \N__31505\
        );

    \I__7011\ : SRMux
    port map (
            O => \N__31538\,
            I => \N__31502\
        );

    \I__7010\ : Span4Mux_v
    port map (
            O => \N__31535\,
            I => \N__31499\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__31532\,
            I => \N__31494\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__31529\,
            I => \N__31494\
        );

    \I__7007\ : Span4Mux_s3_h
    port map (
            O => \N__31526\,
            I => \N__31491\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__31523\,
            I => \N__31486\
        );

    \I__7005\ : Span4Mux_v
    port map (
            O => \N__31514\,
            I => \N__31486\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31483\
        );

    \I__7003\ : Span4Mux_v
    port map (
            O => \N__31508\,
            I => \N__31480\
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__31505\,
            I => \N__31477\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31474\
        );

    \I__7000\ : Span4Mux_v
    port map (
            O => \N__31499\,
            I => \N__31471\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__31494\,
            I => \N__31468\
        );

    \I__6998\ : Sp12to4
    port map (
            O => \N__31491\,
            I => \N__31465\
        );

    \I__6997\ : Span4Mux_v
    port map (
            O => \N__31486\,
            I => \N__31462\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__31483\,
            I => \N__31455\
        );

    \I__6995\ : Span4Mux_v
    port map (
            O => \N__31480\,
            I => \N__31455\
        );

    \I__6994\ : Span4Mux_h
    port map (
            O => \N__31477\,
            I => \N__31455\
        );

    \I__6993\ : Span4Mux_h
    port map (
            O => \N__31474\,
            I => \N__31452\
        );

    \I__6992\ : Odrv4
    port map (
            O => \N__31471\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__31468\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__6990\ : Odrv12
    port map (
            O => \N__31465\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__6989\ : Odrv4
    port map (
            O => \N__31462\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__6988\ : Odrv4
    port map (
            O => \N__31455\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__6987\ : Odrv4
    port map (
            O => \N__31452\,
            I => \POWERLED.N_430_iZ0\
        );

    \I__6986\ : CascadeMux
    port map (
            O => \N__31439\,
            I => \POWERLED.N_5_0_cascade_\
        );

    \I__6985\ : InMux
    port map (
            O => \N__31436\,
            I => \N__31433\
        );

    \I__6984\ : LocalMux
    port map (
            O => \N__31433\,
            I => \POWERLED.N_12_2\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__31430\,
            I => \POWERLED.g0_7_1_cascade_\
        );

    \I__6982\ : InMux
    port map (
            O => \N__31427\,
            I => \N__31424\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__31424\,
            I => \N__31421\
        );

    \I__6980\ : Span4Mux_h
    port map (
            O => \N__31421\,
            I => \N__31418\
        );

    \I__6979\ : Odrv4
    port map (
            O => \N__31418\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_4\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31415\,
            I => \N__31395\
        );

    \I__6977\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31395\
        );

    \I__6976\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31388\
        );

    \I__6975\ : InMux
    port map (
            O => \N__31412\,
            I => \N__31388\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31388\
        );

    \I__6973\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31383\
        );

    \I__6972\ : InMux
    port map (
            O => \N__31409\,
            I => \N__31380\
        );

    \I__6971\ : InMux
    port map (
            O => \N__31408\,
            I => \N__31373\
        );

    \I__6970\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31373\
        );

    \I__6969\ : InMux
    port map (
            O => \N__31406\,
            I => \N__31373\
        );

    \I__6968\ : CascadeMux
    port map (
            O => \N__31405\,
            I => \N__31370\
        );

    \I__6967\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31367\
        );

    \I__6966\ : InMux
    port map (
            O => \N__31403\,
            I => \N__31364\
        );

    \I__6965\ : InMux
    port map (
            O => \N__31402\,
            I => \N__31359\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31359\
        );

    \I__6963\ : InMux
    port map (
            O => \N__31400\,
            I => \N__31356\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__31395\,
            I => \N__31353\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__31388\,
            I => \N__31349\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31342\
        );

    \I__6959\ : InMux
    port map (
            O => \N__31386\,
            I => \N__31337\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__31383\,
            I => \N__31334\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__31380\,
            I => \N__31329\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31329\
        );

    \I__6955\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31326\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__31367\,
            I => \N__31319\
        );

    \I__6953\ : LocalMux
    port map (
            O => \N__31364\,
            I => \N__31319\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__31359\,
            I => \N__31319\
        );

    \I__6951\ : LocalMux
    port map (
            O => \N__31356\,
            I => \N__31314\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__31353\,
            I => \N__31314\
        );

    \I__6949\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31311\
        );

    \I__6948\ : Span4Mux_s0_h
    port map (
            O => \N__31349\,
            I => \N__31308\
        );

    \I__6947\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31303\
        );

    \I__6946\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31303\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31298\
        );

    \I__6944\ : InMux
    port map (
            O => \N__31345\,
            I => \N__31298\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__31342\,
            I => \N__31295\
        );

    \I__6942\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31290\
        );

    \I__6941\ : InMux
    port map (
            O => \N__31340\,
            I => \N__31290\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__31337\,
            I => \N__31283\
        );

    \I__6939\ : Span12Mux_s7_v
    port map (
            O => \N__31334\,
            I => \N__31283\
        );

    \I__6938\ : Span12Mux_s8_v
    port map (
            O => \N__31329\,
            I => \N__31283\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__31326\,
            I => \N__31276\
        );

    \I__6936\ : Span4Mux_v
    port map (
            O => \N__31319\,
            I => \N__31276\
        );

    \I__6935\ : Span4Mux_h
    port map (
            O => \N__31314\,
            I => \N__31276\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__31311\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6933\ : Odrv4
    port map (
            O => \N__31308\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__31303\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6931\ : LocalMux
    port map (
            O => \N__31298\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6930\ : Odrv12
    port map (
            O => \N__31295\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__31290\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6928\ : Odrv12
    port map (
            O => \N__31283\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__31276\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6926\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31249\
        );

    \I__6925\ : CascadeMux
    port map (
            O => \N__31258\,
            I => \N__31246\
        );

    \I__6924\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31235\
        );

    \I__6923\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31235\
        );

    \I__6922\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31235\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__31254\,
            I => \N__31231\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__31253\,
            I => \N__31227\
        );

    \I__6919\ : CascadeMux
    port map (
            O => \N__31252\,
            I => \N__31221\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__31249\,
            I => \N__31212\
        );

    \I__6917\ : InMux
    port map (
            O => \N__31246\,
            I => \N__31207\
        );

    \I__6916\ : InMux
    port map (
            O => \N__31245\,
            I => \N__31207\
        );

    \I__6915\ : InMux
    port map (
            O => \N__31244\,
            I => \N__31204\
        );

    \I__6914\ : InMux
    port map (
            O => \N__31243\,
            I => \N__31199\
        );

    \I__6913\ : InMux
    port map (
            O => \N__31242\,
            I => \N__31199\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__31235\,
            I => \N__31196\
        );

    \I__6911\ : CascadeMux
    port map (
            O => \N__31234\,
            I => \N__31193\
        );

    \I__6910\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31188\
        );

    \I__6909\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31188\
        );

    \I__6908\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31183\
        );

    \I__6907\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31183\
        );

    \I__6906\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31176\
        );

    \I__6905\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31176\
        );

    \I__6904\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31176\
        );

    \I__6903\ : InMux
    port map (
            O => \N__31220\,
            I => \N__31173\
        );

    \I__6902\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31166\
        );

    \I__6901\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31166\
        );

    \I__6900\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31166\
        );

    \I__6899\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31163\
        );

    \I__6898\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31160\
        );

    \I__6897\ : Span4Mux_s3_h
    port map (
            O => \N__31212\,
            I => \N__31157\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__31207\,
            I => \N__31154\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__31204\,
            I => \N__31147\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__31199\,
            I => \N__31147\
        );

    \I__6893\ : Span4Mux_s3_h
    port map (
            O => \N__31196\,
            I => \N__31147\
        );

    \I__6892\ : InMux
    port map (
            O => \N__31193\,
            I => \N__31144\
        );

    \I__6891\ : LocalMux
    port map (
            O => \N__31188\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__31183\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__31176\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__31173\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__31166\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6886\ : LocalMux
    port map (
            O => \N__31163\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__31160\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6884\ : Odrv4
    port map (
            O => \N__31157\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__31154\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__31147\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__31144\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__6880\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31118\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__31118\,
            I => \N__31115\
        );

    \I__6878\ : Span4Mux_v
    port map (
            O => \N__31115\,
            I => \N__31112\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__31112\,
            I => \POWERLED.i2_mux\
        );

    \I__6876\ : InMux
    port map (
            O => \N__31109\,
            I => \N__31101\
        );

    \I__6875\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31098\
        );

    \I__6874\ : InMux
    port map (
            O => \N__31107\,
            I => \N__31095\
        );

    \I__6873\ : InMux
    port map (
            O => \N__31106\,
            I => \N__31090\
        );

    \I__6872\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31090\
        );

    \I__6871\ : InMux
    port map (
            O => \N__31104\,
            I => \N__31087\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__31101\,
            I => \N__31078\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__31098\,
            I => \N__31078\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31078\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__31090\,
            I => \N__31075\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__31087\,
            I => \N__31072\
        );

    \I__6865\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31069\
        );

    \I__6864\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31066\
        );

    \I__6863\ : Span4Mux_v
    port map (
            O => \N__31078\,
            I => \N__31061\
        );

    \I__6862\ : Span4Mux_s0_h
    port map (
            O => \N__31075\,
            I => \N__31061\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__31072\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__31069\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__31066\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__6858\ : Odrv4
    port map (
            O => \N__31061\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__6857\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31049\
        );

    \I__6856\ : LocalMux
    port map (
            O => \N__31049\,
            I => \POWERLED.g1_1cf0\
        );

    \I__6855\ : InMux
    port map (
            O => \N__31046\,
            I => \N__31041\
        );

    \I__6854\ : InMux
    port map (
            O => \N__31045\,
            I => \N__31036\
        );

    \I__6853\ : InMux
    port map (
            O => \N__31044\,
            I => \N__31036\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__31041\,
            I => \N__31032\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__31036\,
            I => \N__31029\
        );

    \I__6850\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31021\
        );

    \I__6849\ : Span4Mux_v
    port map (
            O => \N__31032\,
            I => \N__31011\
        );

    \I__6848\ : Span4Mux_s0_h
    port map (
            O => \N__31029\,
            I => \N__31011\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31008\
        );

    \I__6846\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31005\
        );

    \I__6845\ : InMux
    port map (
            O => \N__31026\,
            I => \N__30998\
        );

    \I__6844\ : InMux
    port map (
            O => \N__31025\,
            I => \N__30998\
        );

    \I__6843\ : InMux
    port map (
            O => \N__31024\,
            I => \N__30998\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__31021\,
            I => \N__30993\
        );

    \I__6841\ : InMux
    port map (
            O => \N__31020\,
            I => \N__30988\
        );

    \I__6840\ : InMux
    port map (
            O => \N__31019\,
            I => \N__30988\
        );

    \I__6839\ : InMux
    port map (
            O => \N__31018\,
            I => \N__30985\
        );

    \I__6838\ : InMux
    port map (
            O => \N__31017\,
            I => \N__30979\
        );

    \I__6837\ : InMux
    port map (
            O => \N__31016\,
            I => \N__30979\
        );

    \I__6836\ : Span4Mux_h
    port map (
            O => \N__31011\,
            I => \N__30972\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__31008\,
            I => \N__30972\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__31005\,
            I => \N__30972\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__30998\,
            I => \N__30969\
        );

    \I__6832\ : InMux
    port map (
            O => \N__30997\,
            I => \N__30966\
        );

    \I__6831\ : CascadeMux
    port map (
            O => \N__30996\,
            I => \N__30963\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__30993\,
            I => \N__30960\
        );

    \I__6829\ : LocalMux
    port map (
            O => \N__30988\,
            I => \N__30955\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__30985\,
            I => \N__30955\
        );

    \I__6827\ : InMux
    port map (
            O => \N__30984\,
            I => \N__30952\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__30979\,
            I => \N__30943\
        );

    \I__6825\ : Span4Mux_v
    port map (
            O => \N__30972\,
            I => \N__30943\
        );

    \I__6824\ : Span4Mux_v
    port map (
            O => \N__30969\,
            I => \N__30943\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30943\
        );

    \I__6822\ : InMux
    port map (
            O => \N__30963\,
            I => \N__30940\
        );

    \I__6821\ : Odrv4
    port map (
            O => \N__30960\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__6820\ : Odrv12
    port map (
            O => \N__30955\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__30952\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__30943\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__30940\,
            I => \POWERLED.dutycycleZ1Z_5\
        );

    \I__6816\ : CascadeMux
    port map (
            O => \N__30929\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_3_cascade_\
        );

    \I__6815\ : CascadeMux
    port map (
            O => \N__30926\,
            I => \N__30923\
        );

    \I__6814\ : InMux
    port map (
            O => \N__30923\,
            I => \N__30920\
        );

    \I__6813\ : LocalMux
    port map (
            O => \N__30920\,
            I => \N__30917\
        );

    \I__6812\ : Span4Mux_v
    port map (
            O => \N__30917\,
            I => \N__30914\
        );

    \I__6811\ : Span4Mux_h
    port map (
            O => \N__30914\,
            I => \N__30911\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__30911\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5\
        );

    \I__6809\ : CascadeMux
    port map (
            O => \N__30908\,
            I => \POWERLED.un1_clk_100khz_32_and_i_0cf0_cascade_\
        );

    \I__6808\ : CascadeMux
    port map (
            O => \N__30905\,
            I => \N__30902\
        );

    \I__6807\ : InMux
    port map (
            O => \N__30902\,
            I => \N__30895\
        );

    \I__6806\ : InMux
    port map (
            O => \N__30901\,
            I => \N__30892\
        );

    \I__6805\ : InMux
    port map (
            O => \N__30900\,
            I => \N__30889\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30899\,
            I => \N__30886\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30883\
        );

    \I__6802\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30879\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__30892\,
            I => \N__30874\
        );

    \I__6800\ : LocalMux
    port map (
            O => \N__30889\,
            I => \N__30874\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__30886\,
            I => \N__30869\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__30883\,
            I => \N__30869\
        );

    \I__6797\ : InMux
    port map (
            O => \N__30882\,
            I => \N__30866\
        );

    \I__6796\ : Span4Mux_s0_h
    port map (
            O => \N__30879\,
            I => \N__30863\
        );

    \I__6795\ : Span4Mux_v
    port map (
            O => \N__30874\,
            I => \N__30858\
        );

    \I__6794\ : Span4Mux_v
    port map (
            O => \N__30869\,
            I => \N__30858\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__30866\,
            I => \N__30855\
        );

    \I__6792\ : Span4Mux_h
    port map (
            O => \N__30863\,
            I => \N__30846\
        );

    \I__6791\ : Span4Mux_h
    port map (
            O => \N__30858\,
            I => \N__30846\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__30855\,
            I => \N__30846\
        );

    \I__6789\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30843\
        );

    \I__6788\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30840\
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__30846\,
            I => \RSMRSTn_fast\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__30843\,
            I => \RSMRSTn_fast\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__30840\,
            I => \RSMRSTn_fast\
        );

    \I__6784\ : CascadeMux
    port map (
            O => \N__30833\,
            I => \N__30829\
        );

    \I__6783\ : InMux
    port map (
            O => \N__30832\,
            I => \N__30824\
        );

    \I__6782\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30824\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__30824\,
            I => \N__30821\
        );

    \I__6780\ : Odrv12
    port map (
            O => \N__30821\,
            I => \POWERLED.un1_clk_100khz_32_and_i_0\
        );

    \I__6779\ : IoInMux
    port map (
            O => \N__30818\,
            I => \N__30814\
        );

    \I__6778\ : IoInMux
    port map (
            O => \N__30817\,
            I => \N__30811\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__30814\,
            I => \N__30804\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30804\
        );

    \I__6775\ : CascadeMux
    port map (
            O => \N__30810\,
            I => \N__30801\
        );

    \I__6774\ : InMux
    port map (
            O => \N__30809\,
            I => \N__30791\
        );

    \I__6773\ : IoSpan4Mux
    port map (
            O => \N__30804\,
            I => \N__30787\
        );

    \I__6772\ : InMux
    port map (
            O => \N__30801\,
            I => \N__30782\
        );

    \I__6771\ : InMux
    port map (
            O => \N__30800\,
            I => \N__30782\
        );

    \I__6770\ : InMux
    port map (
            O => \N__30799\,
            I => \N__30779\
        );

    \I__6769\ : CascadeMux
    port map (
            O => \N__30798\,
            I => \N__30776\
        );

    \I__6768\ : CascadeMux
    port map (
            O => \N__30797\,
            I => \N__30773\
        );

    \I__6767\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30770\
        );

    \I__6766\ : InMux
    port map (
            O => \N__30795\,
            I => \N__30767\
        );

    \I__6765\ : InMux
    port map (
            O => \N__30794\,
            I => \N__30764\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__30791\,
            I => \N__30761\
        );

    \I__6763\ : InMux
    port map (
            O => \N__30790\,
            I => \N__30758\
        );

    \I__6762\ : IoSpan4Mux
    port map (
            O => \N__30787\,
            I => \N__30755\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30782\,
            I => \N__30752\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__30779\,
            I => \N__30749\
        );

    \I__6759\ : InMux
    port map (
            O => \N__30776\,
            I => \N__30746\
        );

    \I__6758\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30743\
        );

    \I__6757\ : LocalMux
    port map (
            O => \N__30770\,
            I => \N__30739\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__30767\,
            I => \N__30730\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__30764\,
            I => \N__30730\
        );

    \I__6754\ : Span4Mux_v
    port map (
            O => \N__30761\,
            I => \N__30730\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30730\
        );

    \I__6752\ : Span4Mux_s2_h
    port map (
            O => \N__30755\,
            I => \N__30724\
        );

    \I__6751\ : Span4Mux_v
    port map (
            O => \N__30752\,
            I => \N__30724\
        );

    \I__6750\ : Span4Mux_h
    port map (
            O => \N__30749\,
            I => \N__30721\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__30746\,
            I => \N__30716\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__30743\,
            I => \N__30716\
        );

    \I__6747\ : InMux
    port map (
            O => \N__30742\,
            I => \N__30713\
        );

    \I__6746\ : Span4Mux_v
    port map (
            O => \N__30739\,
            I => \N__30704\
        );

    \I__6745\ : Span4Mux_v
    port map (
            O => \N__30730\,
            I => \N__30704\
        );

    \I__6744\ : InMux
    port map (
            O => \N__30729\,
            I => \N__30701\
        );

    \I__6743\ : Span4Mux_h
    port map (
            O => \N__30724\,
            I => \N__30698\
        );

    \I__6742\ : Span4Mux_h
    port map (
            O => \N__30721\,
            I => \N__30691\
        );

    \I__6741\ : Span4Mux_s3_h
    port map (
            O => \N__30716\,
            I => \N__30691\
        );

    \I__6740\ : LocalMux
    port map (
            O => \N__30713\,
            I => \N__30691\
        );

    \I__6739\ : InMux
    port map (
            O => \N__30712\,
            I => \N__30688\
        );

    \I__6738\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30681\
        );

    \I__6737\ : InMux
    port map (
            O => \N__30710\,
            I => \N__30681\
        );

    \I__6736\ : InMux
    port map (
            O => \N__30709\,
            I => \N__30681\
        );

    \I__6735\ : Span4Mux_h
    port map (
            O => \N__30704\,
            I => \N__30676\
        );

    \I__6734\ : LocalMux
    port map (
            O => \N__30701\,
            I => \N__30676\
        );

    \I__6733\ : Odrv4
    port map (
            O => \N__30698\,
            I => v5s_enn
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__30691\,
            I => v5s_enn
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__30688\,
            I => v5s_enn
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__30681\,
            I => v5s_enn
        );

    \I__6729\ : Odrv4
    port map (
            O => \N__30676\,
            I => v5s_enn
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__30665\,
            I => \N__30654\
        );

    \I__6727\ : CascadeMux
    port map (
            O => \N__30664\,
            I => \N__30651\
        );

    \I__6726\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30648\
        );

    \I__6725\ : InMux
    port map (
            O => \N__30662\,
            I => \N__30645\
        );

    \I__6724\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30641\
        );

    \I__6723\ : CascadeMux
    port map (
            O => \N__30660\,
            I => \N__30636\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__30659\,
            I => \N__30633\
        );

    \I__6721\ : CascadeMux
    port map (
            O => \N__30658\,
            I => \N__30626\
        );

    \I__6720\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30622\
        );

    \I__6719\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30617\
        );

    \I__6718\ : InMux
    port map (
            O => \N__30651\,
            I => \N__30617\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__30648\,
            I => \N__30611\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30645\,
            I => \N__30611\
        );

    \I__6715\ : CascadeMux
    port map (
            O => \N__30644\,
            I => \N__30608\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__30641\,
            I => \N__30605\
        );

    \I__6713\ : InMux
    port map (
            O => \N__30640\,
            I => \N__30602\
        );

    \I__6712\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30591\
        );

    \I__6711\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30591\
        );

    \I__6710\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30591\
        );

    \I__6709\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30591\
        );

    \I__6708\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30591\
        );

    \I__6707\ : InMux
    port map (
            O => \N__30630\,
            I => \N__30586\
        );

    \I__6706\ : InMux
    port map (
            O => \N__30629\,
            I => \N__30586\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30626\,
            I => \N__30581\
        );

    \I__6704\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30581\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__30622\,
            I => \N__30578\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__30617\,
            I => \N__30571\
        );

    \I__6701\ : InMux
    port map (
            O => \N__30616\,
            I => \N__30568\
        );

    \I__6700\ : Span4Mux_v
    port map (
            O => \N__30611\,
            I => \N__30565\
        );

    \I__6699\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30562\
        );

    \I__6698\ : Span4Mux_v
    port map (
            O => \N__30605\,
            I => \N__30552\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__30602\,
            I => \N__30552\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__30591\,
            I => \N__30552\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__30586\,
            I => \N__30547\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__30581\,
            I => \N__30547\
        );

    \I__6693\ : Span4Mux_s2_h
    port map (
            O => \N__30578\,
            I => \N__30544\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__30577\,
            I => \N__30541\
        );

    \I__6691\ : InMux
    port map (
            O => \N__30576\,
            I => \N__30532\
        );

    \I__6690\ : InMux
    port map (
            O => \N__30575\,
            I => \N__30532\
        );

    \I__6689\ : InMux
    port map (
            O => \N__30574\,
            I => \N__30532\
        );

    \I__6688\ : Span4Mux_s2_h
    port map (
            O => \N__30571\,
            I => \N__30529\
        );

    \I__6687\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30526\
        );

    \I__6686\ : Span4Mux_v
    port map (
            O => \N__30565\,
            I => \N__30523\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__30562\,
            I => \N__30520\
        );

    \I__6684\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30517\
        );

    \I__6683\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30514\
        );

    \I__6682\ : InMux
    port map (
            O => \N__30559\,
            I => \N__30511\
        );

    \I__6681\ : Span4Mux_v
    port map (
            O => \N__30552\,
            I => \N__30508\
        );

    \I__6680\ : Span4Mux_h
    port map (
            O => \N__30547\,
            I => \N__30503\
        );

    \I__6679\ : Span4Mux_v
    port map (
            O => \N__30544\,
            I => \N__30503\
        );

    \I__6678\ : InMux
    port map (
            O => \N__30541\,
            I => \N__30500\
        );

    \I__6677\ : InMux
    port map (
            O => \N__30540\,
            I => \N__30495\
        );

    \I__6676\ : InMux
    port map (
            O => \N__30539\,
            I => \N__30495\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__30532\,
            I => \N__30488\
        );

    \I__6674\ : Span4Mux_v
    port map (
            O => \N__30529\,
            I => \N__30488\
        );

    \I__6673\ : Span4Mux_s2_h
    port map (
            O => \N__30526\,
            I => \N__30488\
        );

    \I__6672\ : Odrv4
    port map (
            O => \N__30523\,
            I => \POWERLED.N_2291_i\
        );

    \I__6671\ : Odrv12
    port map (
            O => \N__30520\,
            I => \POWERLED.N_2291_i\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__30517\,
            I => \POWERLED.N_2291_i\
        );

    \I__6669\ : LocalMux
    port map (
            O => \N__30514\,
            I => \POWERLED.N_2291_i\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__30511\,
            I => \POWERLED.N_2291_i\
        );

    \I__6667\ : Odrv4
    port map (
            O => \N__30508\,
            I => \POWERLED.N_2291_i\
        );

    \I__6666\ : Odrv4
    port map (
            O => \N__30503\,
            I => \POWERLED.N_2291_i\
        );

    \I__6665\ : LocalMux
    port map (
            O => \N__30500\,
            I => \POWERLED.N_2291_i\
        );

    \I__6664\ : LocalMux
    port map (
            O => \N__30495\,
            I => \POWERLED.N_2291_i\
        );

    \I__6663\ : Odrv4
    port map (
            O => \N__30488\,
            I => \POWERLED.N_2291_i\
        );

    \I__6662\ : InMux
    port map (
            O => \N__30467\,
            I => \N__30458\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30458\
        );

    \I__6660\ : InMux
    port map (
            O => \N__30465\,
            I => \N__30458\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__30458\,
            I => \N__30455\
        );

    \I__6658\ : Span4Mux_s3_h
    port map (
            O => \N__30455\,
            I => \N__30452\
        );

    \I__6657\ : Odrv4
    port map (
            O => \N__30452\,
            I => \POWERLED.N_676\
        );

    \I__6656\ : InMux
    port map (
            O => \N__30449\,
            I => \N__30446\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__30446\,
            I => \POWERLED.dutycycle_RNI6SKJ1Z0Z_3\
        );

    \I__6654\ : CascadeMux
    port map (
            O => \N__30443\,
            I => \POWERLED.func_state_RNILP0FZ0Z_1_cascade_\
        );

    \I__6653\ : InMux
    port map (
            O => \N__30440\,
            I => \N__30437\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__30437\,
            I => \POWERLED.N_523\
        );

    \I__6651\ : CascadeMux
    port map (
            O => \N__30434\,
            I => \N__30431\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30431\,
            I => \N__30428\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__30428\,
            I => \POWERLED.G_11_i_o10_1_0\
        );

    \I__6648\ : InMux
    port map (
            O => \N__30425\,
            I => \N__30421\
        );

    \I__6647\ : CascadeMux
    port map (
            O => \N__30424\,
            I => \N__30412\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__30421\,
            I => \N__30409\
        );

    \I__6645\ : InMux
    port map (
            O => \N__30420\,
            I => \N__30406\
        );

    \I__6644\ : InMux
    port map (
            O => \N__30419\,
            I => \N__30401\
        );

    \I__6643\ : InMux
    port map (
            O => \N__30418\,
            I => \N__30401\
        );

    \I__6642\ : InMux
    port map (
            O => \N__30417\,
            I => \N__30397\
        );

    \I__6641\ : CascadeMux
    port map (
            O => \N__30416\,
            I => \N__30391\
        );

    \I__6640\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30387\
        );

    \I__6639\ : InMux
    port map (
            O => \N__30412\,
            I => \N__30384\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__30409\,
            I => \N__30381\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__30406\,
            I => \N__30378\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__30401\,
            I => \N__30375\
        );

    \I__6635\ : CascadeMux
    port map (
            O => \N__30400\,
            I => \N__30372\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__30397\,
            I => \N__30369\
        );

    \I__6633\ : InMux
    port map (
            O => \N__30396\,
            I => \N__30364\
        );

    \I__6632\ : InMux
    port map (
            O => \N__30395\,
            I => \N__30364\
        );

    \I__6631\ : InMux
    port map (
            O => \N__30394\,
            I => \N__30359\
        );

    \I__6630\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30359\
        );

    \I__6629\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30355\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__30387\,
            I => \N__30350\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__30384\,
            I => \N__30350\
        );

    \I__6626\ : Span4Mux_h
    port map (
            O => \N__30381\,
            I => \N__30345\
        );

    \I__6625\ : Span4Mux_v
    port map (
            O => \N__30378\,
            I => \N__30345\
        );

    \I__6624\ : Span4Mux_v
    port map (
            O => \N__30375\,
            I => \N__30342\
        );

    \I__6623\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30339\
        );

    \I__6622\ : Sp12to4
    port map (
            O => \N__30369\,
            I => \N__30332\
        );

    \I__6621\ : LocalMux
    port map (
            O => \N__30364\,
            I => \N__30332\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__30359\,
            I => \N__30332\
        );

    \I__6619\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30329\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__30355\,
            I => \N__30324\
        );

    \I__6617\ : Span4Mux_v
    port map (
            O => \N__30350\,
            I => \N__30324\
        );

    \I__6616\ : Odrv4
    port map (
            O => \N__30345\,
            I => \POWERLED.dutycycle\
        );

    \I__6615\ : Odrv4
    port map (
            O => \N__30342\,
            I => \POWERLED.dutycycle\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__30339\,
            I => \POWERLED.dutycycle\
        );

    \I__6613\ : Odrv12
    port map (
            O => \N__30332\,
            I => \POWERLED.dutycycle\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__30329\,
            I => \POWERLED.dutycycle\
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__30324\,
            I => \POWERLED.dutycycle\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30307\
        );

    \I__6609\ : InMux
    port map (
            O => \N__30310\,
            I => \N__30304\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__30307\,
            I => \N__30299\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__30304\,
            I => \N__30299\
        );

    \I__6606\ : Odrv4
    port map (
            O => \N__30299\,
            I => \N_9_0\
        );

    \I__6605\ : CascadeMux
    port map (
            O => \N__30296\,
            I => \N__30292\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30284\
        );

    \I__6603\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30284\
        );

    \I__6602\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30278\
        );

    \I__6601\ : InMux
    port map (
            O => \N__30290\,
            I => \N__30278\
        );

    \I__6600\ : InMux
    port map (
            O => \N__30289\,
            I => \N__30272\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__30284\,
            I => \N__30268\
        );

    \I__6598\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30265\
        );

    \I__6597\ : LocalMux
    port map (
            O => \N__30278\,
            I => \N__30261\
        );

    \I__6596\ : InMux
    port map (
            O => \N__30277\,
            I => \N__30257\
        );

    \I__6595\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30252\
        );

    \I__6594\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30252\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30249\
        );

    \I__6592\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30246\
        );

    \I__6591\ : Span4Mux_v
    port map (
            O => \N__30268\,
            I => \N__30241\
        );

    \I__6590\ : LocalMux
    port map (
            O => \N__30265\,
            I => \N__30241\
        );

    \I__6589\ : InMux
    port map (
            O => \N__30264\,
            I => \N__30238\
        );

    \I__6588\ : Span12Mux_v
    port map (
            O => \N__30261\,
            I => \N__30235\
        );

    \I__6587\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30232\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__30257\,
            I => \N__30229\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__30252\,
            I => \N__30224\
        );

    \I__6584\ : Span4Mux_s3_h
    port map (
            O => \N__30249\,
            I => \N__30224\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__30246\,
            I => \N__30219\
        );

    \I__6582\ : Span4Mux_v
    port map (
            O => \N__30241\,
            I => \N__30219\
        );

    \I__6581\ : LocalMux
    port map (
            O => \N__30238\,
            I => \RSMRSTn_rep2\
        );

    \I__6580\ : Odrv12
    port map (
            O => \N__30235\,
            I => \RSMRSTn_rep2\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__30232\,
            I => \RSMRSTn_rep2\
        );

    \I__6578\ : Odrv4
    port map (
            O => \N__30229\,
            I => \RSMRSTn_rep2\
        );

    \I__6577\ : Odrv4
    port map (
            O => \N__30224\,
            I => \RSMRSTn_rep2\
        );

    \I__6576\ : Odrv4
    port map (
            O => \N__30219\,
            I => \RSMRSTn_rep2\
        );

    \I__6575\ : CascadeMux
    port map (
            O => \N__30206\,
            I => \N__30201\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__30205\,
            I => \N__30198\
        );

    \I__6573\ : CascadeMux
    port map (
            O => \N__30204\,
            I => \N__30191\
        );

    \I__6572\ : InMux
    port map (
            O => \N__30201\,
            I => \N__30188\
        );

    \I__6571\ : InMux
    port map (
            O => \N__30198\,
            I => \N__30185\
        );

    \I__6570\ : InMux
    port map (
            O => \N__30197\,
            I => \N__30182\
        );

    \I__6569\ : InMux
    port map (
            O => \N__30196\,
            I => \N__30179\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__30195\,
            I => \N__30176\
        );

    \I__6567\ : InMux
    port map (
            O => \N__30194\,
            I => \N__30172\
        );

    \I__6566\ : InMux
    port map (
            O => \N__30191\,
            I => \N__30169\
        );

    \I__6565\ : LocalMux
    port map (
            O => \N__30188\,
            I => \N__30166\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__30185\,
            I => \N__30163\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30160\
        );

    \I__6562\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30157\
        );

    \I__6561\ : InMux
    port map (
            O => \N__30176\,
            I => \N__30154\
        );

    \I__6560\ : CascadeMux
    port map (
            O => \N__30175\,
            I => \N__30151\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__30172\,
            I => \N__30141\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__30169\,
            I => \N__30141\
        );

    \I__6557\ : Span4Mux_v
    port map (
            O => \N__30166\,
            I => \N__30141\
        );

    \I__6556\ : Span4Mux_h
    port map (
            O => \N__30163\,
            I => \N__30141\
        );

    \I__6555\ : Span4Mux_v
    port map (
            O => \N__30160\,
            I => \N__30135\
        );

    \I__6554\ : Span4Mux_v
    port map (
            O => \N__30157\,
            I => \N__30135\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30132\
        );

    \I__6552\ : InMux
    port map (
            O => \N__30151\,
            I => \N__30127\
        );

    \I__6551\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30127\
        );

    \I__6550\ : Span4Mux_v
    port map (
            O => \N__30141\,
            I => \N__30124\
        );

    \I__6549\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30121\
        );

    \I__6548\ : Span4Mux_h
    port map (
            O => \N__30135\,
            I => \N__30118\
        );

    \I__6547\ : Odrv12
    port map (
            O => \N__30132\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__30127\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__30124\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__30121\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6543\ : Odrv4
    port map (
            O => \N__30118\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__6542\ : InMux
    port map (
            O => \N__30107\,
            I => \N__30104\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__30104\,
            I => \POWERLED.N_488\
        );

    \I__6540\ : InMux
    port map (
            O => \N__30101\,
            I => \N__30098\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30095\
        );

    \I__6538\ : Sp12to4
    port map (
            O => \N__30095\,
            I => \N__30092\
        );

    \I__6537\ : Odrv12
    port map (
            O => \N__30092\,
            I => \POWERLED.N_540_1\
        );

    \I__6536\ : InMux
    port map (
            O => \N__30089\,
            I => \N__30086\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__30086\,
            I => \N__30083\
        );

    \I__6534\ : Span4Mux_h
    port map (
            O => \N__30083\,
            I => \N__30079\
        );

    \I__6533\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30076\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__30079\,
            I => \POWERLED_un1_dutycycle_172_m0_0\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__30076\,
            I => \POWERLED_un1_dutycycle_172_m0_0\
        );

    \I__6530\ : InMux
    port map (
            O => \N__30071\,
            I => \N__30065\
        );

    \I__6529\ : InMux
    port map (
            O => \N__30070\,
            I => \N__30062\
        );

    \I__6528\ : InMux
    port map (
            O => \N__30069\,
            I => \N__30059\
        );

    \I__6527\ : InMux
    port map (
            O => \N__30068\,
            I => \N__30056\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__30065\,
            I => \N__30047\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__30062\,
            I => \N__30047\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__30059\,
            I => \N__30044\
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__30056\,
            I => \N__30041\
        );

    \I__6522\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30034\
        );

    \I__6521\ : InMux
    port map (
            O => \N__30054\,
            I => \N__30034\
        );

    \I__6520\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30034\
        );

    \I__6519\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30030\
        );

    \I__6518\ : Span4Mux_v
    port map (
            O => \N__30047\,
            I => \N__30027\
        );

    \I__6517\ : Span4Mux_s2_h
    port map (
            O => \N__30044\,
            I => \N__30024\
        );

    \I__6516\ : Span4Mux_v
    port map (
            O => \N__30041\,
            I => \N__30019\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__30034\,
            I => \N__30019\
        );

    \I__6514\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30016\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__30013\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__30027\,
            I => \POWERLED.N_435\
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__30024\,
            I => \POWERLED.N_435\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__30019\,
            I => \POWERLED.N_435\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__30016\,
            I => \POWERLED.N_435\
        );

    \I__6508\ : Odrv12
    port map (
            O => \N__30013\,
            I => \POWERLED.N_435\
        );

    \I__6507\ : InMux
    port map (
            O => \N__30002\,
            I => \N__29999\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__29999\,
            I => \N__29996\
        );

    \I__6505\ : Span4Mux_v
    port map (
            O => \N__29996\,
            I => \N__29992\
        );

    \I__6504\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29989\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__29992\,
            I => \POWERLED.func_state_RNI_4Z0Z_1\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__29989\,
            I => \POWERLED.func_state_RNI_4Z0Z_1\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29981\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__29981\,
            I => \POWERLED.un1_dutycycle_172_m0_ns_1_0\
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__29978\,
            I => \POWERLED.func_state_RNI_4Z0Z_1_cascade_\
        );

    \I__6498\ : InMux
    port map (
            O => \N__29975\,
            I => \N__29972\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__29972\,
            I => \POWERLED.dutycycle_RNI5DLRZ0Z_5\
        );

    \I__6496\ : InMux
    port map (
            O => \N__29969\,
            I => \N__29965\
        );

    \I__6495\ : InMux
    port map (
            O => \N__29968\,
            I => \N__29962\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__29965\,
            I => \N__29955\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__29962\,
            I => \N__29952\
        );

    \I__6492\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29949\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29960\,
            I => \N__29946\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29940\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29940\
        );

    \I__6488\ : Span4Mux_v
    port map (
            O => \N__29955\,
            I => \N__29934\
        );

    \I__6487\ : Span4Mux_s1_h
    port map (
            O => \N__29952\,
            I => \N__29934\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__29949\,
            I => \N__29929\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__29946\,
            I => \N__29929\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__29945\,
            I => \N__29925\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__29940\,
            I => \N__29922\
        );

    \I__6482\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29919\
        );

    \I__6481\ : Span4Mux_h
    port map (
            O => \N__29934\,
            I => \N__29916\
        );

    \I__6480\ : Span12Mux_s7_v
    port map (
            O => \N__29929\,
            I => \N__29913\
        );

    \I__6479\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29908\
        );

    \I__6478\ : InMux
    port map (
            O => \N__29925\,
            I => \N__29908\
        );

    \I__6477\ : Odrv12
    port map (
            O => \N__29922\,
            I => \SUSWARN_N_rep1\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__29919\,
            I => \SUSWARN_N_rep1\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__29916\,
            I => \SUSWARN_N_rep1\
        );

    \I__6474\ : Odrv12
    port map (
            O => \N__29913\,
            I => \SUSWARN_N_rep1\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__29908\,
            I => \SUSWARN_N_rep1\
        );

    \I__6472\ : CascadeMux
    port map (
            O => \N__29897\,
            I => \POWERLED.dutycycle_RNI7ABC3Z0Z_5_cascade_\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__29894\,
            I => \N__29890\
        );

    \I__6470\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29880\
        );

    \I__6469\ : InMux
    port map (
            O => \N__29890\,
            I => \N__29880\
        );

    \I__6468\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29877\
        );

    \I__6467\ : CascadeMux
    port map (
            O => \N__29888\,
            I => \N__29874\
        );

    \I__6466\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29867\
        );

    \I__6465\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29867\
        );

    \I__6464\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29864\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29861\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__29877\,
            I => \N__29858\
        );

    \I__6461\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29853\
        );

    \I__6460\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29853\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__29872\,
            I => \N__29850\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__29867\,
            I => \N__29838\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__29864\,
            I => \N__29835\
        );

    \I__6456\ : Span4Mux_v
    port map (
            O => \N__29861\,
            I => \N__29832\
        );

    \I__6455\ : Span4Mux_h
    port map (
            O => \N__29858\,
            I => \N__29827\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__29853\,
            I => \N__29827\
        );

    \I__6453\ : InMux
    port map (
            O => \N__29850\,
            I => \N__29820\
        );

    \I__6452\ : InMux
    port map (
            O => \N__29849\,
            I => \N__29820\
        );

    \I__6451\ : InMux
    port map (
            O => \N__29848\,
            I => \N__29820\
        );

    \I__6450\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29817\
        );

    \I__6449\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29812\
        );

    \I__6448\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29812\
        );

    \I__6447\ : InMux
    port map (
            O => \N__29844\,
            I => \N__29803\
        );

    \I__6446\ : InMux
    port map (
            O => \N__29843\,
            I => \N__29803\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29803\
        );

    \I__6444\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29803\
        );

    \I__6443\ : Span4Mux_v
    port map (
            O => \N__29838\,
            I => \N__29798\
        );

    \I__6442\ : Span4Mux_h
    port map (
            O => \N__29835\,
            I => \N__29798\
        );

    \I__6441\ : Span4Mux_h
    port map (
            O => \N__29832\,
            I => \N__29793\
        );

    \I__6440\ : Span4Mux_v
    port map (
            O => \N__29827\,
            I => \N__29793\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29790\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__29817\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__29812\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__29803\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__6435\ : Odrv4
    port map (
            O => \N__29798\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__6434\ : Odrv4
    port map (
            O => \N__29793\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__6433\ : Odrv4
    port map (
            O => \N__29790\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__6432\ : InMux
    port map (
            O => \N__29777\,
            I => \N__29774\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__29774\,
            I => \N__29771\
        );

    \I__6430\ : Span4Mux_v
    port map (
            O => \N__29771\,
            I => \N__29768\
        );

    \I__6429\ : Odrv4
    port map (
            O => \N__29768\,
            I => \POWERLED.g2_1_1\
        );

    \I__6428\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29762\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__29762\,
            I => v5s_ok
        );

    \I__6426\ : InMux
    port map (
            O => \N__29759\,
            I => \N__29756\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__29756\,
            I => \N__29753\
        );

    \I__6424\ : Span4Mux_v
    port map (
            O => \N__29753\,
            I => \N__29750\
        );

    \I__6423\ : Odrv4
    port map (
            O => \N__29750\,
            I => vccst_cpu_ok
        );

    \I__6422\ : CascadeMux
    port map (
            O => \N__29747\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_1_cascade_\
        );

    \I__6421\ : InMux
    port map (
            O => \N__29744\,
            I => \N__29741\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__29741\,
            I => \N__29738\
        );

    \I__6419\ : Span12Mux_v
    port map (
            O => \N__29738\,
            I => \N__29735\
        );

    \I__6418\ : Odrv12
    port map (
            O => \N__29735\,
            I => v33s_ok
        );

    \I__6417\ : IoInMux
    port map (
            O => \N__29732\,
            I => \N__29729\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__29729\,
            I => \N__29726\
        );

    \I__6415\ : Span4Mux_s2_v
    port map (
            O => \N__29726\,
            I => \N__29723\
        );

    \I__6414\ : Span4Mux_v
    port map (
            O => \N__29723\,
            I => \N__29720\
        );

    \I__6413\ : Span4Mux_v
    port map (
            O => \N__29720\,
            I => \N__29717\
        );

    \I__6412\ : Odrv4
    port map (
            O => \N__29717\,
            I => vccin_en
        );

    \I__6411\ : InMux
    port map (
            O => \N__29714\,
            I => \N__29711\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__29711\,
            I => \N__29707\
        );

    \I__6409\ : InMux
    port map (
            O => \N__29710\,
            I => \N__29704\
        );

    \I__6408\ : Span4Mux_v
    port map (
            O => \N__29707\,
            I => \N__29698\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__29704\,
            I => \N__29698\
        );

    \I__6406\ : InMux
    port map (
            O => \N__29703\,
            I => \N__29694\
        );

    \I__6405\ : Span4Mux_h
    port map (
            O => \N__29698\,
            I => \N__29691\
        );

    \I__6404\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29688\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__29694\,
            I => \POWERLED.N_253\
        );

    \I__6402\ : Odrv4
    port map (
            O => \N__29691\,
            I => \POWERLED.N_253\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__29688\,
            I => \POWERLED.N_253\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__29681\,
            I => \N__29676\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__29680\,
            I => \N__29673\
        );

    \I__6398\ : InMux
    port map (
            O => \N__29679\,
            I => \N__29669\
        );

    \I__6397\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29664\
        );

    \I__6396\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29664\
        );

    \I__6395\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29661\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__29669\,
            I => \N__29658\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__29664\,
            I => \N__29653\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__29661\,
            I => \N__29653\
        );

    \I__6391\ : Span4Mux_h
    port map (
            O => \N__29658\,
            I => \N__29650\
        );

    \I__6390\ : Odrv12
    port map (
            O => \N__29653\,
            I => \POWERLED.func_state_RNI_6Z0Z_1\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__29650\,
            I => \POWERLED.func_state_RNI_6Z0Z_1\
        );

    \I__6388\ : InMux
    port map (
            O => \N__29645\,
            I => \N__29642\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__29642\,
            I => \N__29638\
        );

    \I__6386\ : InMux
    port map (
            O => \N__29641\,
            I => \N__29635\
        );

    \I__6385\ : Odrv12
    port map (
            O => \N__29638\,
            I => \POWERLED.g1_1\
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__29635\,
            I => \POWERLED.g1_1\
        );

    \I__6383\ : CascadeMux
    port map (
            O => \N__29630\,
            I => \POWERLED.func_state_RNI_6Z0Z_1_cascade_\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__29627\,
            I => \POWERLED.N_2361_0_cascade_\
        );

    \I__6381\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29618\
        );

    \I__6380\ : InMux
    port map (
            O => \N__29623\,
            I => \N__29618\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__29618\,
            I => \N__29615\
        );

    \I__6378\ : Odrv4
    port map (
            O => \N__29615\,
            I => \N_6_0\
        );

    \I__6377\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29609\
        );

    \I__6376\ : LocalMux
    port map (
            O => \N__29609\,
            I => \POWERLED.dutycycle_e_N_6L11_1\
        );

    \I__6375\ : CascadeMux
    port map (
            O => \N__29606\,
            I => \POWERLED.dutycycle_RNI2MQDZ0Z_4_cascade_\
        );

    \I__6374\ : CascadeMux
    port map (
            O => \N__29603\,
            I => \N__29600\
        );

    \I__6373\ : InMux
    port map (
            O => \N__29600\,
            I => \N__29597\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__29597\,
            I => \POWERLED.dutycycle_RNIOGRSZ0Z_4\
        );

    \I__6371\ : CascadeMux
    port map (
            O => \N__29594\,
            I => \POWERLED.un1_func_state25_6_0_0_a6_1_0_cascade_\
        );

    \I__6370\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29588\
        );

    \I__6369\ : LocalMux
    port map (
            O => \N__29588\,
            I => \N__29585\
        );

    \I__6368\ : Odrv12
    port map (
            O => \N__29585\,
            I => \POWERLED.un1_func_state25_6_0_o_N_4\
        );

    \I__6367\ : InMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__29579\,
            I => \POWERLED.un1_func_state25_6_0_0_0_2_1\
        );

    \I__6365\ : CascadeMux
    port map (
            O => \N__29576\,
            I => \POWERLED.un1_func_state25_6_0_o_N_5_cascade_\
        );

    \I__6364\ : InMux
    port map (
            O => \N__29573\,
            I => \N__29563\
        );

    \I__6363\ : CascadeMux
    port map (
            O => \N__29572\,
            I => \N__29560\
        );

    \I__6362\ : CascadeMux
    port map (
            O => \N__29571\,
            I => \N__29556\
        );

    \I__6361\ : InMux
    port map (
            O => \N__29570\,
            I => \N__29552\
        );

    \I__6360\ : InMux
    port map (
            O => \N__29569\,
            I => \N__29547\
        );

    \I__6359\ : InMux
    port map (
            O => \N__29568\,
            I => \N__29547\
        );

    \I__6358\ : InMux
    port map (
            O => \N__29567\,
            I => \N__29542\
        );

    \I__6357\ : InMux
    port map (
            O => \N__29566\,
            I => \N__29542\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__29563\,
            I => \N__29539\
        );

    \I__6355\ : InMux
    port map (
            O => \N__29560\,
            I => \N__29535\
        );

    \I__6354\ : InMux
    port map (
            O => \N__29559\,
            I => \N__29532\
        );

    \I__6353\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29525\
        );

    \I__6352\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29525\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__29552\,
            I => \N__29522\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__29547\,
            I => \N__29517\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__29542\,
            I => \N__29517\
        );

    \I__6348\ : Span4Mux_v
    port map (
            O => \N__29539\,
            I => \N__29514\
        );

    \I__6347\ : CascadeMux
    port map (
            O => \N__29538\,
            I => \N__29511\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__29535\,
            I => \N__29503\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__29532\,
            I => \N__29503\
        );

    \I__6344\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29498\
        );

    \I__6343\ : InMux
    port map (
            O => \N__29530\,
            I => \N__29498\
        );

    \I__6342\ : LocalMux
    port map (
            O => \N__29525\,
            I => \N__29495\
        );

    \I__6341\ : Span4Mux_h
    port map (
            O => \N__29522\,
            I => \N__29492\
        );

    \I__6340\ : Span4Mux_h
    port map (
            O => \N__29517\,
            I => \N__29487\
        );

    \I__6339\ : Span4Mux_h
    port map (
            O => \N__29514\,
            I => \N__29487\
        );

    \I__6338\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29478\
        );

    \I__6337\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29478\
        );

    \I__6336\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29478\
        );

    \I__6335\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29478\
        );

    \I__6334\ : Odrv12
    port map (
            O => \N__29503\,
            I => \POWERLED.N_421\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__29498\,
            I => \POWERLED.N_421\
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__29495\,
            I => \POWERLED.N_421\
        );

    \I__6331\ : Odrv4
    port map (
            O => \N__29492\,
            I => \POWERLED.N_421\
        );

    \I__6330\ : Odrv4
    port map (
            O => \N__29487\,
            I => \POWERLED.N_421\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__29478\,
            I => \POWERLED.N_421\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__29465\,
            I => \POWERLED.un1_func_state25_6_0_0_0_2_cascade_\
        );

    \I__6327\ : InMux
    port map (
            O => \N__29462\,
            I => \N__29453\
        );

    \I__6326\ : InMux
    port map (
            O => \N__29461\,
            I => \N__29453\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__29460\,
            I => \N__29449\
        );

    \I__6324\ : CEMux
    port map (
            O => \N__29459\,
            I => \N__29443\
        );

    \I__6323\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29440\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__29453\,
            I => \N__29437\
        );

    \I__6321\ : CEMux
    port map (
            O => \N__29452\,
            I => \N__29432\
        );

    \I__6320\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29423\
        );

    \I__6319\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29423\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29423\
        );

    \I__6317\ : InMux
    port map (
            O => \N__29446\,
            I => \N__29423\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__29443\,
            I => \N__29420\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__29440\,
            I => \N__29417\
        );

    \I__6314\ : Span4Mux_v
    port map (
            O => \N__29437\,
            I => \N__29414\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__29436\,
            I => \N__29408\
        );

    \I__6312\ : CascadeMux
    port map (
            O => \N__29435\,
            I => \N__29403\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__29432\,
            I => \N__29397\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__29423\,
            I => \N__29397\
        );

    \I__6309\ : Span4Mux_v
    port map (
            O => \N__29420\,
            I => \N__29390\
        );

    \I__6308\ : Span4Mux_v
    port map (
            O => \N__29417\,
            I => \N__29390\
        );

    \I__6307\ : Span4Mux_h
    port map (
            O => \N__29414\,
            I => \N__29390\
        );

    \I__6306\ : CascadeMux
    port map (
            O => \N__29413\,
            I => \N__29386\
        );

    \I__6305\ : CEMux
    port map (
            O => \N__29412\,
            I => \N__29382\
        );

    \I__6304\ : CEMux
    port map (
            O => \N__29411\,
            I => \N__29379\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29370\
        );

    \I__6302\ : InMux
    port map (
            O => \N__29407\,
            I => \N__29370\
        );

    \I__6301\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29370\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29403\,
            I => \N__29370\
        );

    \I__6299\ : InMux
    port map (
            O => \N__29402\,
            I => \N__29364\
        );

    \I__6298\ : Span4Mux_s3_v
    port map (
            O => \N__29397\,
            I => \N__29359\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__29390\,
            I => \N__29359\
        );

    \I__6296\ : CEMux
    port map (
            O => \N__29389\,
            I => \N__29352\
        );

    \I__6295\ : InMux
    port map (
            O => \N__29386\,
            I => \N__29352\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29352\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__29382\,
            I => \N__29345\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__29379\,
            I => \N__29345\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__29370\,
            I => \N__29345\
        );

    \I__6290\ : CEMux
    port map (
            O => \N__29369\,
            I => \N__29338\
        );

    \I__6289\ : InMux
    port map (
            O => \N__29368\,
            I => \N__29338\
        );

    \I__6288\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29338\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__29364\,
            I => \POWERLED.func_state_RNI31IBHZ0Z_0\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__29359\,
            I => \POWERLED.func_state_RNI31IBHZ0Z_0\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__29352\,
            I => \POWERLED.func_state_RNI31IBHZ0Z_0\
        );

    \I__6284\ : Odrv4
    port map (
            O => \N__29345\,
            I => \POWERLED.func_state_RNI31IBHZ0Z_0\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__29338\,
            I => \POWERLED.func_state_RNI31IBHZ0Z_0\
        );

    \I__6282\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29324\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__29324\,
            I => \N__29321\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__29321\,
            I => \POWERLED.N_6_2\
        );

    \I__6279\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29315\,
            I => \N__29311\
        );

    \I__6277\ : InMux
    port map (
            O => \N__29314\,
            I => \N__29306\
        );

    \I__6276\ : Span4Mux_v
    port map (
            O => \N__29311\,
            I => \N__29303\
        );

    \I__6275\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29298\
        );

    \I__6274\ : InMux
    port map (
            O => \N__29309\,
            I => \N__29298\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__29306\,
            I => \N__29295\
        );

    \I__6272\ : IoSpan4Mux
    port map (
            O => \N__29303\,
            I => \N__29289\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__29298\,
            I => \N__29289\
        );

    \I__6270\ : Span12Mux_v
    port map (
            O => \N__29295\,
            I => \N__29286\
        );

    \I__6269\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29283\
        );

    \I__6268\ : Span4Mux_s2_h
    port map (
            O => \N__29289\,
            I => \N__29280\
        );

    \I__6267\ : Odrv12
    port map (
            O => \N__29286\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__29283\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__6265\ : Odrv4
    port map (
            O => \N__29280\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__29273\,
            I => \N__29270\
        );

    \I__6263\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29267\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__29267\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0\
        );

    \I__6261\ : InMux
    port map (
            O => \N__29264\,
            I => \N__29257\
        );

    \I__6260\ : InMux
    port map (
            O => \N__29263\,
            I => \N__29254\
        );

    \I__6259\ : InMux
    port map (
            O => \N__29262\,
            I => \N__29251\
        );

    \I__6258\ : InMux
    port map (
            O => \N__29261\,
            I => \N__29248\
        );

    \I__6257\ : CascadeMux
    port map (
            O => \N__29260\,
            I => \N__29242\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29235\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__29254\,
            I => \N__29235\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__29251\,
            I => \N__29232\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__29248\,
            I => \N__29229\
        );

    \I__6252\ : InMux
    port map (
            O => \N__29247\,
            I => \N__29226\
        );

    \I__6251\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29221\
        );

    \I__6250\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29221\
        );

    \I__6249\ : InMux
    port map (
            O => \N__29242\,
            I => \N__29216\
        );

    \I__6248\ : InMux
    port map (
            O => \N__29241\,
            I => \N__29216\
        );

    \I__6247\ : InMux
    port map (
            O => \N__29240\,
            I => \N__29213\
        );

    \I__6246\ : Span4Mux_v
    port map (
            O => \N__29235\,
            I => \N__29208\
        );

    \I__6245\ : Span4Mux_h
    port map (
            O => \N__29232\,
            I => \N__29208\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__29229\,
            I => \N__29205\
        );

    \I__6243\ : LocalMux
    port map (
            O => \N__29226\,
            I => \N__29202\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__29221\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__29216\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__29213\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6239\ : Odrv4
    port map (
            O => \N__29208\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6238\ : Odrv4
    port map (
            O => \N__29205\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6237\ : Odrv12
    port map (
            O => \N__29202\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__6236\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29182\
        );

    \I__6235\ : InMux
    port map (
            O => \N__29188\,
            I => \N__29177\
        );

    \I__6234\ : InMux
    port map (
            O => \N__29187\,
            I => \N__29177\
        );

    \I__6233\ : InMux
    port map (
            O => \N__29186\,
            I => \N__29174\
        );

    \I__6232\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29171\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__29182\,
            I => \N__29168\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__29177\,
            I => \N__29165\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29160\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__29171\,
            I => \N__29160\
        );

    \I__6227\ : Span4Mux_v
    port map (
            O => \N__29168\,
            I => \N__29157\
        );

    \I__6226\ : Span12Mux_s7_v
    port map (
            O => \N__29165\,
            I => \N__29154\
        );

    \I__6225\ : Odrv12
    port map (
            O => \N__29160\,
            I => \POWERLED.func_state_RNI_3Z0Z_1\
        );

    \I__6224\ : Odrv4
    port map (
            O => \N__29157\,
            I => \POWERLED.func_state_RNI_3Z0Z_1\
        );

    \I__6223\ : Odrv12
    port map (
            O => \N__29154\,
            I => \POWERLED.func_state_RNI_3Z0Z_1\
        );

    \I__6222\ : CascadeMux
    port map (
            O => \N__29147\,
            I => \POWERLED.func_state_RNIBVNSZ0Z_0_cascade_\
        );

    \I__6221\ : InMux
    port map (
            O => \N__29144\,
            I => \N__29141\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__29141\,
            I => \POWERLED.func_state_1_m0_1_1\
        );

    \I__6219\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29135\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__29135\,
            I => \POWERLED.un1_func_state25_6_0_o_N_7_2\
        );

    \I__6217\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29127\
        );

    \I__6216\ : CascadeMux
    port map (
            O => \N__29131\,
            I => \N__29124\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__29130\,
            I => \N__29120\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__29127\,
            I => \N__29112\
        );

    \I__6213\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29103\
        );

    \I__6212\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29103\
        );

    \I__6211\ : InMux
    port map (
            O => \N__29120\,
            I => \N__29103\
        );

    \I__6210\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29103\
        );

    \I__6209\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29096\
        );

    \I__6208\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29096\
        );

    \I__6207\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29096\
        );

    \I__6206\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29093\
        );

    \I__6205\ : Span4Mux_v
    port map (
            O => \N__29112\,
            I => \N__29090\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29087\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29082\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__29093\,
            I => \N__29082\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__29090\,
            I => \N__29079\
        );

    \I__6200\ : Span4Mux_h
    port map (
            O => \N__29087\,
            I => \N__29076\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__29082\,
            I => \N__29073\
        );

    \I__6198\ : Odrv4
    port map (
            O => \N__29079\,
            I => rsmrst_pwrgd_signal
        );

    \I__6197\ : Odrv4
    port map (
            O => \N__29076\,
            I => rsmrst_pwrgd_signal
        );

    \I__6196\ : Odrv4
    port map (
            O => \N__29073\,
            I => rsmrst_pwrgd_signal
        );

    \I__6195\ : InMux
    port map (
            O => \N__29066\,
            I => \N__29063\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__29063\,
            I => \N__29060\
        );

    \I__6193\ : Odrv4
    port map (
            O => \N__29060\,
            I => \POWERLED.count_off_0_13\
        );

    \I__6192\ : InMux
    port map (
            O => \N__29057\,
            I => \N__29054\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__29054\,
            I => \N__29050\
        );

    \I__6190\ : InMux
    port map (
            O => \N__29053\,
            I => \N__29047\
        );

    \I__6189\ : Odrv4
    port map (
            O => \N__29050\,
            I => \POWERLED.count_off_1_13\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__29047\,
            I => \POWERLED.count_off_1_13\
        );

    \I__6187\ : CascadeMux
    port map (
            O => \N__29042\,
            I => \N__29039\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29036\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__29036\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__6184\ : CascadeMux
    port map (
            O => \N__29033\,
            I => \N__29029\
        );

    \I__6183\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29026\
        );

    \I__6182\ : InMux
    port map (
            O => \N__29029\,
            I => \N__29023\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__29026\,
            I => \N__29020\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__29023\,
            I => \N__29017\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__29020\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__29017\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__29012\,
            I => \POWERLED.count_offZ0Z_13_cascade_\
        );

    \I__6176\ : InMux
    port map (
            O => \N__29009\,
            I => \N__29005\
        );

    \I__6175\ : InMux
    port map (
            O => \N__29008\,
            I => \N__29002\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__29005\,
            I => \N__28999\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__29002\,
            I => \N__28996\
        );

    \I__6172\ : Span4Mux_v
    port map (
            O => \N__28999\,
            I => \N__28993\
        );

    \I__6171\ : Span4Mux_v
    port map (
            O => \N__28996\,
            I => \N__28990\
        );

    \I__6170\ : Span4Mux_v
    port map (
            O => \N__28993\,
            I => \N__28985\
        );

    \I__6169\ : Span4Mux_v
    port map (
            O => \N__28990\,
            I => \N__28985\
        );

    \I__6168\ : Odrv4
    port map (
            O => \N__28985\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__6167\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28979\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__28979\,
            I => \N__28976\
        );

    \I__6165\ : Odrv4
    port map (
            O => \N__28976\,
            I => \POWERLED.un34_clk_100khz_10\
        );

    \I__6164\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28970\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__28970\,
            I => \POWERLED.count_off_0_0\
        );

    \I__6162\ : CascadeMux
    port map (
            O => \N__28967\,
            I => \POWERLED.count_off_1_0_cascade_\
        );

    \I__6161\ : CascadeMux
    port map (
            O => \N__28964\,
            I => \N__28958\
        );

    \I__6160\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28951\
        );

    \I__6159\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28951\
        );

    \I__6158\ : InMux
    port map (
            O => \N__28961\,
            I => \N__28951\
        );

    \I__6157\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28948\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__28951\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__28948\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__6154\ : CascadeMux
    port map (
            O => \N__28943\,
            I => \POWERLED.count_offZ0Z_0_cascade_\
        );

    \I__6153\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28937\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__28937\,
            I => \POWERLED.count_off_RNIZ0Z_1\
        );

    \I__6151\ : CascadeMux
    port map (
            O => \N__28934\,
            I => \N__28912\
        );

    \I__6150\ : InMux
    port map (
            O => \N__28933\,
            I => \N__28905\
        );

    \I__6149\ : InMux
    port map (
            O => \N__28932\,
            I => \N__28905\
        );

    \I__6148\ : InMux
    port map (
            O => \N__28931\,
            I => \N__28905\
        );

    \I__6147\ : InMux
    port map (
            O => \N__28930\,
            I => \N__28900\
        );

    \I__6146\ : InMux
    port map (
            O => \N__28929\,
            I => \N__28900\
        );

    \I__6145\ : InMux
    port map (
            O => \N__28928\,
            I => \N__28893\
        );

    \I__6144\ : InMux
    port map (
            O => \N__28927\,
            I => \N__28893\
        );

    \I__6143\ : InMux
    port map (
            O => \N__28926\,
            I => \N__28893\
        );

    \I__6142\ : InMux
    port map (
            O => \N__28925\,
            I => \N__28884\
        );

    \I__6141\ : InMux
    port map (
            O => \N__28924\,
            I => \N__28884\
        );

    \I__6140\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28884\
        );

    \I__6139\ : InMux
    port map (
            O => \N__28922\,
            I => \N__28884\
        );

    \I__6138\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28875\
        );

    \I__6137\ : InMux
    port map (
            O => \N__28920\,
            I => \N__28875\
        );

    \I__6136\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28875\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28918\,
            I => \N__28875\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28866\
        );

    \I__6133\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28866\
        );

    \I__6132\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28866\
        );

    \I__6131\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28866\
        );

    \I__6130\ : LocalMux
    port map (
            O => \N__28905\,
            I => \N__28859\
        );

    \I__6129\ : LocalMux
    port map (
            O => \N__28900\,
            I => \N__28859\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__28893\,
            I => \N__28859\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__28884\,
            I => \N__28854\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__28875\,
            I => \N__28854\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__28866\,
            I => \POWERLED.N_123\
        );

    \I__6124\ : Odrv12
    port map (
            O => \N__28859\,
            I => \POWERLED.N_123\
        );

    \I__6123\ : Odrv4
    port map (
            O => \N__28854\,
            I => \POWERLED.N_123\
        );

    \I__6122\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28844\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__28844\,
            I => \POWERLED.count_off_0_1\
        );

    \I__6120\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \POWERLED.count_off_RNIZ0Z_1_cascade_\
        );

    \I__6119\ : InMux
    port map (
            O => \N__28838\,
            I => \N__28834\
        );

    \I__6118\ : InMux
    port map (
            O => \N__28837\,
            I => \N__28830\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28827\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28833\,
            I => \N__28824\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__28830\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__28827\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__6113\ : LocalMux
    port map (
            O => \N__28824\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__6112\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28811\
        );

    \I__6111\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28811\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__28811\,
            I => \POWERLED.count_off_1_2\
        );

    \I__6109\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28805\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__28805\,
            I => \POWERLED.count_off_0_2\
        );

    \I__6107\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28796\
        );

    \I__6106\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28796\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__28796\,
            I => \POWERLED.count_off_1_5\
        );

    \I__6104\ : InMux
    port map (
            O => \N__28793\,
            I => \N__28790\
        );

    \I__6103\ : LocalMux
    port map (
            O => \N__28790\,
            I => \POWERLED.count_off_0_5\
        );

    \I__6102\ : InMux
    port map (
            O => \N__28787\,
            I => \N__28784\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__28784\,
            I => \POWERLED.count_off_0_6\
        );

    \I__6100\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28775\
        );

    \I__6099\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28775\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__28775\,
            I => \POWERLED.count_off_1_6\
        );

    \I__6097\ : CascadeMux
    port map (
            O => \N__28772\,
            I => \N__28769\
        );

    \I__6096\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28766\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__28766\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__6094\ : CascadeMux
    port map (
            O => \N__28763\,
            I => \N__28759\
        );

    \I__6093\ : InMux
    port map (
            O => \N__28762\,
            I => \N__28756\
        );

    \I__6092\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28753\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__28756\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__28753\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__6089\ : CascadeMux
    port map (
            O => \N__28748\,
            I => \N__28744\
        );

    \I__6088\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28741\
        );

    \I__6087\ : InMux
    port map (
            O => \N__28744\,
            I => \N__28738\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__28741\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__28738\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__6084\ : CascadeMux
    port map (
            O => \N__28733\,
            I => \POWERLED.count_offZ0Z_6_cascade_\
        );

    \I__6083\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28727\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28724\
        );

    \I__6081\ : Odrv4
    port map (
            O => \N__28724\,
            I => \POWERLED.un34_clk_100khz_9\
        );

    \I__6080\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28718\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__28718\,
            I => \POWERLED.count_off_0_11\
        );

    \I__6078\ : InMux
    port map (
            O => \N__28715\,
            I => \N__28712\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__28712\,
            I => \N__28708\
        );

    \I__6076\ : InMux
    port map (
            O => \N__28711\,
            I => \N__28705\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__28708\,
            I => \POWERLED.count_off_1_11\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__28705\,
            I => \POWERLED.count_off_1_11\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__28700\,
            I => \N__28696\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28699\,
            I => \N__28693\
        );

    \I__6071\ : InMux
    port map (
            O => \N__28696\,
            I => \N__28690\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__28693\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__28690\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__28685\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\
        );

    \I__6067\ : CascadeMux
    port map (
            O => \N__28682\,
            I => \POWERLED.count_clkZ0Z_0_cascade_\
        );

    \I__6066\ : CascadeMux
    port map (
            O => \N__28679\,
            I => \POWERLED.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__6065\ : InMux
    port map (
            O => \N__28676\,
            I => \N__28671\
        );

    \I__6064\ : InMux
    port map (
            O => \N__28675\,
            I => \N__28666\
        );

    \I__6063\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28666\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__28671\,
            I => \N__28660\
        );

    \I__6061\ : LocalMux
    port map (
            O => \N__28666\,
            I => \N__28660\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28657\
        );

    \I__6059\ : Span4Mux_h
    port map (
            O => \N__28660\,
            I => \N__28654\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__28657\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__28654\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__6056\ : CascadeMux
    port map (
            O => \N__28649\,
            I => \POWERLED.count_clkZ0Z_1_cascade_\
        );

    \I__6055\ : InMux
    port map (
            O => \N__28646\,
            I => \N__28643\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__28643\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__6053\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28637\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__28637\,
            I => \N__28633\
        );

    \I__6051\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28630\
        );

    \I__6050\ : Span4Mux_s3_v
    port map (
            O => \N__28633\,
            I => \N__28627\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__28630\,
            I => \N__28624\
        );

    \I__6048\ : Odrv4
    port map (
            O => \N__28627\,
            I => \POWERLED.count_off_1_14\
        );

    \I__6047\ : Odrv4
    port map (
            O => \N__28624\,
            I => \POWERLED.count_off_1_14\
        );

    \I__6046\ : InMux
    port map (
            O => \N__28619\,
            I => \N__28616\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__28616\,
            I => \POWERLED.count_off_0_14\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28610\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__28610\,
            I => \N__28607\
        );

    \I__6042\ : Span4Mux_h
    port map (
            O => \N__28607\,
            I => \N__28604\
        );

    \I__6041\ : Span4Mux_v
    port map (
            O => \N__28604\,
            I => \N__28600\
        );

    \I__6040\ : InMux
    port map (
            O => \N__28603\,
            I => \N__28597\
        );

    \I__6039\ : Span4Mux_v
    port map (
            O => \N__28600\,
            I => \N__28594\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__28597\,
            I => \POWERLED.count_off_1_7\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__28594\,
            I => \POWERLED.count_off_1_7\
        );

    \I__6036\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28586\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__28586\,
            I => \N__28583\
        );

    \I__6034\ : Span12Mux_s7_h
    port map (
            O => \N__28583\,
            I => \N__28580\
        );

    \I__6033\ : Span12Mux_v
    port map (
            O => \N__28580\,
            I => \N__28577\
        );

    \I__6032\ : Odrv12
    port map (
            O => \N__28577\,
            I => \POWERLED.count_off_0_7\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28574\,
            I => \N__28571\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__28571\,
            I => \N__28568\
        );

    \I__6029\ : Span4Mux_h
    port map (
            O => \N__28568\,
            I => \N__28565\
        );

    \I__6028\ : Span4Mux_v
    port map (
            O => \N__28565\,
            I => \N__28561\
        );

    \I__6027\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28558\
        );

    \I__6026\ : Span4Mux_v
    port map (
            O => \N__28561\,
            I => \N__28555\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__28558\,
            I => \POWERLED.count_off_1_8\
        );

    \I__6024\ : Odrv4
    port map (
            O => \N__28555\,
            I => \POWERLED.count_off_1_8\
        );

    \I__6023\ : CascadeMux
    port map (
            O => \N__28550\,
            I => \N__28547\
        );

    \I__6022\ : InMux
    port map (
            O => \N__28547\,
            I => \N__28544\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__28544\,
            I => \N__28541\
        );

    \I__6020\ : Span12Mux_s8_h
    port map (
            O => \N__28541\,
            I => \N__28538\
        );

    \I__6019\ : Span12Mux_v
    port map (
            O => \N__28538\,
            I => \N__28535\
        );

    \I__6018\ : Odrv12
    port map (
            O => \N__28535\,
            I => \POWERLED.count_off_0_8\
        );

    \I__6017\ : CascadeMux
    port map (
            O => \N__28532\,
            I => \POWERLED.N_518_cascade_\
        );

    \I__6016\ : InMux
    port map (
            O => \N__28529\,
            I => \N__28522\
        );

    \I__6015\ : InMux
    port map (
            O => \N__28528\,
            I => \N__28515\
        );

    \I__6014\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28515\
        );

    \I__6013\ : InMux
    port map (
            O => \N__28526\,
            I => \N__28515\
        );

    \I__6012\ : CascadeMux
    port map (
            O => \N__28525\,
            I => \N__28512\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__28522\,
            I => \N__28505\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__28515\,
            I => \N__28502\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28499\
        );

    \I__6008\ : InMux
    port map (
            O => \N__28511\,
            I => \N__28496\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__28510\,
            I => \N__28492\
        );

    \I__6006\ : CascadeMux
    port map (
            O => \N__28509\,
            I => \N__28487\
        );

    \I__6005\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28484\
        );

    \I__6004\ : Span12Mux_s7_h
    port map (
            O => \N__28505\,
            I => \N__28481\
        );

    \I__6003\ : Span4Mux_h
    port map (
            O => \N__28502\,
            I => \N__28476\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__28499\,
            I => \N__28476\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__28496\,
            I => \N__28473\
        );

    \I__6000\ : InMux
    port map (
            O => \N__28495\,
            I => \N__28470\
        );

    \I__5999\ : InMux
    port map (
            O => \N__28492\,
            I => \N__28463\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28491\,
            I => \N__28463\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28490\,
            I => \N__28463\
        );

    \I__5996\ : InMux
    port map (
            O => \N__28487\,
            I => \N__28460\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__28484\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5994\ : Odrv12
    port map (
            O => \N__28481\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__28476\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5992\ : Odrv4
    port map (
            O => \N__28473\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__28470\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__28463\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__28460\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__5988\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28442\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__28442\,
            I => \POWERLED.dutycycle_RNIE3861_0Z0Z_12\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__28439\,
            I => \POWERLED.N_520_cascade_\
        );

    \I__5985\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28430\
        );

    \I__5984\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28430\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__28430\,
            I => \N__28427\
        );

    \I__5982\ : Span4Mux_h
    port map (
            O => \N__28427\,
            I => \N__28424\
        );

    \I__5981\ : Odrv4
    port map (
            O => \N__28424\,
            I => \POWERLED.dutycycle_RNIPK9V4Z0Z_12\
        );

    \I__5980\ : InMux
    port map (
            O => \N__28421\,
            I => \N__28417\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28414\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__28417\,
            I => \N__28409\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__28414\,
            I => \N__28409\
        );

    \I__5976\ : Span12Mux_s6_v
    port map (
            O => \N__28409\,
            I => \N__28406\
        );

    \I__5975\ : Odrv12
    port map (
            O => \N__28406\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIN405GZ0\
        );

    \I__5974\ : InMux
    port map (
            O => \N__28403\,
            I => \N__28400\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__28400\,
            I => \POWERLED.count_off_0_15\
        );

    \I__5972\ : CascadeMux
    port map (
            O => \N__28397\,
            I => \N__28394\
        );

    \I__5971\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28391\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__28391\,
            I => \N__28388\
        );

    \I__5969\ : Span4Mux_v
    port map (
            O => \N__28388\,
            I => \N__28385\
        );

    \I__5968\ : Span4Mux_v
    port map (
            O => \N__28385\,
            I => \N__28381\
        );

    \I__5967\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__28381\,
            I => \POWERLED.count_off_RNI8AQHZ0Z_10\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__28378\,
            I => \POWERLED.count_off_RNI8AQHZ0Z_10\
        );

    \I__5964\ : InMux
    port map (
            O => \N__28373\,
            I => \N__28370\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__28370\,
            I => \N__28367\
        );

    \I__5962\ : Odrv12
    port map (
            O => \N__28367\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_5\
        );

    \I__5961\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28360\
        );

    \I__5960\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28357\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__28360\,
            I => \N__28352\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__28357\,
            I => \N__28352\
        );

    \I__5957\ : Odrv12
    port map (
            O => \N__28352\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__5956\ : InMux
    port map (
            O => \N__28349\,
            I => \N__28343\
        );

    \I__5955\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28343\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__28343\,
            I => \N__28340\
        );

    \I__5953\ : Odrv12
    port map (
            O => \N__28340\,
            I => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__28337\,
            I => \N__28334\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28334\,
            I => \N__28331\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__28331\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__28328\,
            I => \POWERLED.N_514_cascade_\
        );

    \I__5948\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28319\
        );

    \I__5947\ : InMux
    port map (
            O => \N__28324\,
            I => \N__28319\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__28319\,
            I => \N__28316\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__28316\,
            I => \N__28313\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__28313\,
            I => \POWERLED.dutycycle_RNIHDMC5Z0Z_11\
        );

    \I__5943\ : InMux
    port map (
            O => \N__28310\,
            I => \N__28305\
        );

    \I__5942\ : InMux
    port map (
            O => \N__28309\,
            I => \N__28299\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__28308\,
            I => \N__28295\
        );

    \I__5940\ : LocalMux
    port map (
            O => \N__28305\,
            I => \N__28292\
        );

    \I__5939\ : InMux
    port map (
            O => \N__28304\,
            I => \N__28285\
        );

    \I__5938\ : InMux
    port map (
            O => \N__28303\,
            I => \N__28285\
        );

    \I__5937\ : InMux
    port map (
            O => \N__28302\,
            I => \N__28285\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__28299\,
            I => \N__28281\
        );

    \I__5935\ : CascadeMux
    port map (
            O => \N__28298\,
            I => \N__28275\
        );

    \I__5934\ : InMux
    port map (
            O => \N__28295\,
            I => \N__28268\
        );

    \I__5933\ : Span4Mux_v
    port map (
            O => \N__28292\,
            I => \N__28265\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__28285\,
            I => \N__28262\
        );

    \I__5931\ : InMux
    port map (
            O => \N__28284\,
            I => \N__28259\
        );

    \I__5930\ : Span4Mux_h
    port map (
            O => \N__28281\,
            I => \N__28256\
        );

    \I__5929\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28251\
        );

    \I__5928\ : InMux
    port map (
            O => \N__28279\,
            I => \N__28251\
        );

    \I__5927\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28246\
        );

    \I__5926\ : InMux
    port map (
            O => \N__28275\,
            I => \N__28246\
        );

    \I__5925\ : InMux
    port map (
            O => \N__28274\,
            I => \N__28241\
        );

    \I__5924\ : InMux
    port map (
            O => \N__28273\,
            I => \N__28241\
        );

    \I__5923\ : InMux
    port map (
            O => \N__28272\,
            I => \N__28236\
        );

    \I__5922\ : InMux
    port map (
            O => \N__28271\,
            I => \N__28236\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__28268\,
            I => \N__28233\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__28265\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5919\ : Odrv12
    port map (
            O => \N__28262\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__28259\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5917\ : Odrv4
    port map (
            O => \N__28256\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__28251\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__28246\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__28241\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__28236\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5912\ : Odrv4
    port map (
            O => \N__28233\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__5911\ : InMux
    port map (
            O => \N__28214\,
            I => \N__28211\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__28211\,
            I => \N__28208\
        );

    \I__5909\ : Odrv12
    port map (
            O => \N__28208\,
            I => \POWERLED.N_508\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__28205\,
            I => \POWERLED.N_512_cascade_\
        );

    \I__5907\ : InMux
    port map (
            O => \N__28202\,
            I => \N__28195\
        );

    \I__5906\ : InMux
    port map (
            O => \N__28201\,
            I => \N__28190\
        );

    \I__5905\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28190\
        );

    \I__5904\ : InMux
    port map (
            O => \N__28199\,
            I => \N__28187\
        );

    \I__5903\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28184\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__28195\,
            I => \N__28176\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28171\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__28187\,
            I => \N__28171\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__28184\,
            I => \N__28168\
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__28183\,
            I => \N__28159\
        );

    \I__5897\ : CascadeMux
    port map (
            O => \N__28182\,
            I => \N__28156\
        );

    \I__5896\ : InMux
    port map (
            O => \N__28181\,
            I => \N__28151\
        );

    \I__5895\ : InMux
    port map (
            O => \N__28180\,
            I => \N__28151\
        );

    \I__5894\ : CascadeMux
    port map (
            O => \N__28179\,
            I => \N__28148\
        );

    \I__5893\ : Span4Mux_v
    port map (
            O => \N__28176\,
            I => \N__28141\
        );

    \I__5892\ : Span4Mux_v
    port map (
            O => \N__28171\,
            I => \N__28141\
        );

    \I__5891\ : Span4Mux_v
    port map (
            O => \N__28168\,
            I => \N__28141\
        );

    \I__5890\ : InMux
    port map (
            O => \N__28167\,
            I => \N__28136\
        );

    \I__5889\ : InMux
    port map (
            O => \N__28166\,
            I => \N__28136\
        );

    \I__5888\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28131\
        );

    \I__5887\ : InMux
    port map (
            O => \N__28164\,
            I => \N__28131\
        );

    \I__5886\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28122\
        );

    \I__5885\ : InMux
    port map (
            O => \N__28162\,
            I => \N__28122\
        );

    \I__5884\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28122\
        );

    \I__5883\ : InMux
    port map (
            O => \N__28156\,
            I => \N__28122\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28119\
        );

    \I__5881\ : InMux
    port map (
            O => \N__28148\,
            I => \N__28116\
        );

    \I__5880\ : Odrv4
    port map (
            O => \N__28141\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__28136\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__28131\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__28122\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__28119\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__28116\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5874\ : InMux
    port map (
            O => \N__28103\,
            I => \N__28100\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__28100\,
            I => \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_11\
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__28097\,
            I => \POWERLED.N_526_cascade_\
        );

    \I__5871\ : InMux
    port map (
            O => \N__28094\,
            I => \N__28091\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__28091\,
            I => \POWERLED.un1_clk_100khz_47_and_i_1\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__28088\,
            I => \N__28084\
        );

    \I__5868\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28079\
        );

    \I__5867\ : InMux
    port map (
            O => \N__28084\,
            I => \N__28079\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__28076\
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__28076\,
            I => \POWERLED.dutycycle_en_11\
        );

    \I__5864\ : InMux
    port map (
            O => \N__28073\,
            I => \N__28070\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__28070\,
            I => \POWERLED.N_2075_tz_tz\
        );

    \I__5862\ : CascadeMux
    port map (
            O => \N__28067\,
            I => \N__28063\
        );

    \I__5861\ : InMux
    port map (
            O => \N__28066\,
            I => \N__28060\
        );

    \I__5860\ : InMux
    port map (
            O => \N__28063\,
            I => \N__28057\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__28060\,
            I => \N__28052\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28049\
        );

    \I__5857\ : InMux
    port map (
            O => \N__28056\,
            I => \N__28046\
        );

    \I__5856\ : InMux
    port map (
            O => \N__28055\,
            I => \N__28043\
        );

    \I__5855\ : Span4Mux_s1_h
    port map (
            O => \N__28052\,
            I => \N__28040\
        );

    \I__5854\ : Span4Mux_v
    port map (
            O => \N__28049\,
            I => \N__28033\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__28033\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28033\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__28040\,
            I => \N__28030\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__28033\,
            I => \N__28027\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__28030\,
            I => \POWERLED.N_600\
        );

    \I__5848\ : Odrv4
    port map (
            O => \N__28027\,
            I => \POWERLED.N_600\
        );

    \I__5847\ : InMux
    port map (
            O => \N__28022\,
            I => \N__28019\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__28019\,
            I => \N__28016\
        );

    \I__5845\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__28013\
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__28013\,
            I => \POWERLED.count_clk_en_0\
        );

    \I__5843\ : CascadeMux
    port map (
            O => \N__28010\,
            I => \N__28007\
        );

    \I__5842\ : InMux
    port map (
            O => \N__28007\,
            I => \N__28004\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__28004\,
            I => \N__28001\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__28001\,
            I => \POWERLED.N_443\
        );

    \I__5839\ : InMux
    port map (
            O => \N__27998\,
            I => \N__27995\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__27995\,
            I => \N__27992\
        );

    \I__5837\ : Odrv12
    port map (
            O => \N__27992\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_1\
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__27989\,
            I => \POWERLED.N_443_cascade_\
        );

    \I__5835\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27982\
        );

    \I__5834\ : InMux
    port map (
            O => \N__27985\,
            I => \N__27978\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__27982\,
            I => \N__27975\
        );

    \I__5832\ : CascadeMux
    port map (
            O => \N__27981\,
            I => \N__27972\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__27978\,
            I => \N__27969\
        );

    \I__5830\ : Span4Mux_v
    port map (
            O => \N__27975\,
            I => \N__27966\
        );

    \I__5829\ : InMux
    port map (
            O => \N__27972\,
            I => \N__27963\
        );

    \I__5828\ : Span4Mux_v
    port map (
            O => \N__27969\,
            I => \N__27960\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__27966\,
            I => \N__27955\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__27963\,
            I => \N__27955\
        );

    \I__5825\ : Span4Mux_v
    port map (
            O => \N__27960\,
            I => \N__27952\
        );

    \I__5824\ : Span4Mux_v
    port map (
            O => \N__27955\,
            I => \N__27949\
        );

    \I__5823\ : Odrv4
    port map (
            O => \N__27952\,
            I => \POWERLED.count_clk_RNINSEUCZ0Z_7\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__27949\,
            I => \POWERLED.count_clk_RNINSEUCZ0Z_7\
        );

    \I__5821\ : InMux
    port map (
            O => \N__27944\,
            I => \N__27940\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__27943\,
            I => \N__27937\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__27940\,
            I => \N__27934\
        );

    \I__5818\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27931\
        );

    \I__5817\ : Span4Mux_v
    port map (
            O => \N__27934\,
            I => \N__27928\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__27931\,
            I => \N__27924\
        );

    \I__5815\ : Span4Mux_v
    port map (
            O => \N__27928\,
            I => \N__27921\
        );

    \I__5814\ : InMux
    port map (
            O => \N__27927\,
            I => \N__27918\
        );

    \I__5813\ : Span4Mux_s2_h
    port map (
            O => \N__27924\,
            I => \N__27915\
        );

    \I__5812\ : IoSpan4Mux
    port map (
            O => \N__27921\,
            I => \N__27910\
        );

    \I__5811\ : LocalMux
    port map (
            O => \N__27918\,
            I => \N__27910\
        );

    \I__5810\ : Span4Mux_v
    port map (
            O => \N__27915\,
            I => \N__27905\
        );

    \I__5809\ : Span4Mux_s2_h
    port map (
            O => \N__27910\,
            I => \N__27905\
        );

    \I__5808\ : Odrv4
    port map (
            O => \N__27905\,
            I => \POWERLED.N_668\
        );

    \I__5807\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27899\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__27899\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_2\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__27896\,
            I => \N__27892\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__27895\,
            I => \N__27887\
        );

    \I__5803\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27883\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27891\,
            I => \N__27878\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27890\,
            I => \N__27878\
        );

    \I__5800\ : InMux
    port map (
            O => \N__27887\,
            I => \N__27875\
        );

    \I__5799\ : CascadeMux
    port map (
            O => \N__27886\,
            I => \N__27870\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__27883\,
            I => \N__27865\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__27878\,
            I => \N__27862\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__27875\,
            I => \N__27859\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27874\,
            I => \N__27854\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27854\
        );

    \I__5793\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27851\
        );

    \I__5792\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27846\
        );

    \I__5791\ : InMux
    port map (
            O => \N__27868\,
            I => \N__27846\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__27865\,
            I => \N__27843\
        );

    \I__5789\ : Span4Mux_v
    port map (
            O => \N__27862\,
            I => \N__27838\
        );

    \I__5788\ : Span4Mux_h
    port map (
            O => \N__27859\,
            I => \N__27838\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__27854\,
            I => \N__27833\
        );

    \I__5786\ : LocalMux
    port map (
            O => \N__27851\,
            I => \N__27833\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__27846\,
            I => \N__27830\
        );

    \I__5784\ : Odrv4
    port map (
            O => \N__27843\,
            I => \N_247\
        );

    \I__5783\ : Odrv4
    port map (
            O => \N__27838\,
            I => \N_247\
        );

    \I__5782\ : Odrv12
    port map (
            O => \N__27833\,
            I => \N_247\
        );

    \I__5781\ : Odrv12
    port map (
            O => \N__27830\,
            I => \N_247\
        );

    \I__5780\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27818\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__27818\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_0\
        );

    \I__5778\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27811\
        );

    \I__5777\ : CascadeMux
    port map (
            O => \N__27814\,
            I => \N__27808\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__27811\,
            I => \N__27803\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27800\
        );

    \I__5774\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27792\
        );

    \I__5773\ : InMux
    port map (
            O => \N__27806\,
            I => \N__27792\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__27803\,
            I => \N__27787\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__27800\,
            I => \N__27787\
        );

    \I__5770\ : CascadeMux
    port map (
            O => \N__27799\,
            I => \N__27784\
        );

    \I__5769\ : CascadeMux
    port map (
            O => \N__27798\,
            I => \N__27781\
        );

    \I__5768\ : InMux
    port map (
            O => \N__27797\,
            I => \N__27778\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__27792\,
            I => \N__27775\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__27787\,
            I => \N__27772\
        );

    \I__5765\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27767\
        );

    \I__5764\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27767\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__27778\,
            I => \RSMRSTn_rep1\
        );

    \I__5762\ : Odrv4
    port map (
            O => \N__27775\,
            I => \RSMRSTn_rep1\
        );

    \I__5761\ : Odrv4
    port map (
            O => \N__27772\,
            I => \RSMRSTn_rep1\
        );

    \I__5760\ : LocalMux
    port map (
            O => \N__27767\,
            I => \RSMRSTn_rep1\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__27758\,
            I => \POWERLED.N_506_cascade_\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__27755\,
            I => \N__27752\
        );

    \I__5757\ : InMux
    port map (
            O => \N__27752\,
            I => \N__27749\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__27749\,
            I => \N__27746\
        );

    \I__5755\ : Span4Mux_h
    port map (
            O => \N__27746\,
            I => \N__27743\
        );

    \I__5754\ : Odrv4
    port map (
            O => \N__27743\,
            I => \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_10\
        );

    \I__5753\ : InMux
    port map (
            O => \N__27740\,
            I => \N__27737\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__27737\,
            I => \N__27734\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__27734\,
            I => \N__27731\
        );

    \I__5750\ : Odrv4
    port map (
            O => \N__27731\,
            I => \POWERLED.g0_i_0_1\
        );

    \I__5749\ : CascadeMux
    port map (
            O => \N__27728\,
            I => \POWERLED.un1_dutycycle_53_25_0_tz_1_1_cascade_\
        );

    \I__5748\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27721\
        );

    \I__5747\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27718\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__27721\,
            I => \N__27713\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27718\,
            I => \N__27713\
        );

    \I__5744\ : Span4Mux_h
    port map (
            O => \N__27713\,
            I => \N__27710\
        );

    \I__5743\ : Odrv4
    port map (
            O => \N__27710\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_4\
        );

    \I__5742\ : CascadeMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__5741\ : InMux
    port map (
            O => \N__27704\,
            I => \N__27700\
        );

    \I__5740\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27697\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__27700\,
            I => \N__27694\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__27697\,
            I => \N__27689\
        );

    \I__5737\ : Span4Mux_s2_h
    port map (
            O => \N__27694\,
            I => \N__27689\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__27689\,
            I => \N__27686\
        );

    \I__5735\ : Odrv4
    port map (
            O => \N__27686\,
            I => \POWERLED.func_state_RNI_0Z0Z_1\
        );

    \I__5734\ : InMux
    port map (
            O => \N__27683\,
            I => \N__27678\
        );

    \I__5733\ : InMux
    port map (
            O => \N__27682\,
            I => \N__27673\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__27681\,
            I => \N__27670\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__27678\,
            I => \N__27667\
        );

    \I__5730\ : InMux
    port map (
            O => \N__27677\,
            I => \N__27662\
        );

    \I__5729\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27662\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__27673\,
            I => \N__27657\
        );

    \I__5727\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27652\
        );

    \I__5726\ : Span4Mux_v
    port map (
            O => \N__27667\,
            I => \N__27647\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__27662\,
            I => \N__27647\
        );

    \I__5724\ : InMux
    port map (
            O => \N__27661\,
            I => \N__27642\
        );

    \I__5723\ : InMux
    port map (
            O => \N__27660\,
            I => \N__27642\
        );

    \I__5722\ : Span4Mux_s1_h
    port map (
            O => \N__27657\,
            I => \N__27639\
        );

    \I__5721\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27634\
        );

    \I__5720\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27634\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__27652\,
            I => \N__27629\
        );

    \I__5718\ : Span4Mux_h
    port map (
            O => \N__27647\,
            I => \N__27629\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27626\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__27639\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__27634\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5714\ : Odrv4
    port map (
            O => \N__27629\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5713\ : Odrv12
    port map (
            O => \N__27626\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__27617\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_1_cascade_\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__27614\,
            I => \POWERLED.func_state_RNI_8Z0Z_1_cascade_\
        );

    \I__5710\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27608\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__27608\,
            I => \N__27605\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__27605\,
            I => \POWERLED.func_state_RNIMQ0F_0Z0Z_1\
        );

    \I__5707\ : InMux
    port map (
            O => \N__27602\,
            I => \N__27599\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__27599\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__27596\,
            I => \POWERLED.func_state_RNIMQ0F_0Z0Z_1_cascade_\
        );

    \I__5704\ : InMux
    port map (
            O => \N__27593\,
            I => \N__27590\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__27590\,
            I => \POWERLED.dutycycle_RNI2MQDZ0Z_7\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__27587\,
            I => \N__27584\
        );

    \I__5701\ : InMux
    port map (
            O => \N__27584\,
            I => \N__27581\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__27581\,
            I => \N__27578\
        );

    \I__5699\ : Odrv12
    port map (
            O => \N__27578\,
            I => \POWERLED.dutycycle_RNIEBSB1Z0Z_7\
        );

    \I__5698\ : InMux
    port map (
            O => \N__27575\,
            I => \N__27572\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__27572\,
            I => \N__27569\
        );

    \I__5696\ : Span12Mux_s3_h
    port map (
            O => \N__27569\,
            I => \N__27566\
        );

    \I__5695\ : Odrv12
    port map (
            O => \N__27566\,
            I => \POWERLED.N_545\
        );

    \I__5694\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27560\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__27560\,
            I => \N__27557\
        );

    \I__5692\ : Span4Mux_s2_h
    port map (
            O => \N__27557\,
            I => \N__27554\
        );

    \I__5691\ : Odrv4
    port map (
            O => \N__27554\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\
        );

    \I__5690\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27545\
        );

    \I__5689\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27545\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__27545\,
            I => \N__27542\
        );

    \I__5687\ : Span4Mux_h
    port map (
            O => \N__27542\,
            I => \N__27539\
        );

    \I__5686\ : Span4Mux_v
    port map (
            O => \N__27539\,
            I => \N__27536\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__27536\,
            I => \POWERLED.N_71\
        );

    \I__5684\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27527\
        );

    \I__5683\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27527\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__27527\,
            I => \N__27524\
        );

    \I__5681\ : Span4Mux_s2_h
    port map (
            O => \N__27524\,
            I => \N__27521\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__27521\,
            I => \POWERLED.un1_clk_100khz_36_and_i_0_a2_d\
        );

    \I__5679\ : InMux
    port map (
            O => \N__27518\,
            I => \N__27515\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__27515\,
            I => \N__27512\
        );

    \I__5677\ : Odrv12
    port map (
            O => \N__27512\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__5676\ : InMux
    port map (
            O => \N__27509\,
            I => \N__27506\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__27506\,
            I => \POWERLED.dutycycle_e_1_4\
        );

    \I__5674\ : CascadeMux
    port map (
            O => \N__27503\,
            I => \POWERLED.dutycycle_e_1_4_cascade_\
        );

    \I__5673\ : InMux
    port map (
            O => \N__27500\,
            I => \N__27494\
        );

    \I__5672\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27494\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__27494\,
            I => \POWERLED.func_state_RNIJ17U4Z0Z_1\
        );

    \I__5670\ : InMux
    port map (
            O => \N__27491\,
            I => \N__27487\
        );

    \I__5669\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27484\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__27487\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__27484\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__5666\ : InMux
    port map (
            O => \N__27479\,
            I => \N__27476\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__27476\,
            I => \N__27473\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__27473\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__5663\ : InMux
    port map (
            O => \N__27470\,
            I => \N__27467\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27467\,
            I => \POWERLED.dutycycle_e_1_7\
        );

    \I__5661\ : InMux
    port map (
            O => \N__27464\,
            I => \N__27460\
        );

    \I__5660\ : InMux
    port map (
            O => \N__27463\,
            I => \N__27457\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__27460\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__27457\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__27452\,
            I => \POWERLED.dutycycle_e_1_7_cascade_\
        );

    \I__5656\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27443\
        );

    \I__5655\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27443\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__27443\,
            I => \POWERLED.func_state_RNI9S7D5Z0Z_1\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__27440\,
            I => \POWERLED.dutycycleZ1Z_6_cascade_\
        );

    \I__5652\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27433\
        );

    \I__5651\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27430\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__27433\,
            I => \N__27425\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27425\
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__27425\,
            I => \POWERLED.N_133\
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__27422\,
            I => \N__27417\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__27421\,
            I => \N__27412\
        );

    \I__5645\ : InMux
    port map (
            O => \N__27420\,
            I => \N__27409\
        );

    \I__5644\ : InMux
    port map (
            O => \N__27417\,
            I => \N__27406\
        );

    \I__5643\ : InMux
    port map (
            O => \N__27416\,
            I => \N__27403\
        );

    \I__5642\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27400\
        );

    \I__5641\ : InMux
    port map (
            O => \N__27412\,
            I => \N__27397\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__27409\,
            I => \N__27393\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__27406\,
            I => \N__27390\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__27403\,
            I => \N__27386\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__27400\,
            I => \N__27381\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__27397\,
            I => \N__27381\
        );

    \I__5635\ : InMux
    port map (
            O => \N__27396\,
            I => \N__27378\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__27393\,
            I => \N__27373\
        );

    \I__5633\ : Span4Mux_v
    port map (
            O => \N__27390\,
            I => \N__27373\
        );

    \I__5632\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27370\
        );

    \I__5631\ : Span4Mux_s2_h
    port map (
            O => \N__27386\,
            I => \N__27365\
        );

    \I__5630\ : Span4Mux_h
    port map (
            O => \N__27381\,
            I => \N__27365\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__27378\,
            I => \N__27362\
        );

    \I__5628\ : Odrv4
    port map (
            O => \N__27373\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__27370\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__27365\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5625\ : Odrv4
    port map (
            O => \N__27362\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__27353\,
            I => \N__27349\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27352\,
            I => \N__27342\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27342\
        );

    \I__5621\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27333\
        );

    \I__5620\ : InMux
    port map (
            O => \N__27347\,
            I => \N__27333\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__27342\,
            I => \N__27329\
        );

    \I__5618\ : InMux
    port map (
            O => \N__27341\,
            I => \N__27326\
        );

    \I__5617\ : InMux
    port map (
            O => \N__27340\,
            I => \N__27321\
        );

    \I__5616\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27321\
        );

    \I__5615\ : InMux
    port map (
            O => \N__27338\,
            I => \N__27318\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__27333\,
            I => \N__27313\
        );

    \I__5613\ : InMux
    port map (
            O => \N__27332\,
            I => \N__27310\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__27329\,
            I => \N__27307\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__27326\,
            I => \N__27300\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__27321\,
            I => \N__27300\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__27318\,
            I => \N__27300\
        );

    \I__5608\ : InMux
    port map (
            O => \N__27317\,
            I => \N__27297\
        );

    \I__5607\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27294\
        );

    \I__5606\ : Span4Mux_s3_h
    port map (
            O => \N__27313\,
            I => \N__27289\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__27310\,
            I => \N__27289\
        );

    \I__5604\ : Span4Mux_v
    port map (
            O => \N__27307\,
            I => \N__27284\
        );

    \I__5603\ : Span4Mux_v
    port map (
            O => \N__27300\,
            I => \N__27284\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__27297\,
            I => \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__27294\,
            I => \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__27289\,
            I => \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0\
        );

    \I__5599\ : Odrv4
    port map (
            O => \N__27284\,
            I => \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0\
        );

    \I__5598\ : InMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__27272\,
            I => \POWERLED.N_490\
        );

    \I__5596\ : InMux
    port map (
            O => \N__27269\,
            I => \N__27266\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__27266\,
            I => \N__27263\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__27263\,
            I => \N__27260\
        );

    \I__5593\ : Odrv4
    port map (
            O => \N__27260\,
            I => \POWERLED.g1_0_2\
        );

    \I__5592\ : CascadeMux
    port map (
            O => \N__27257\,
            I => \POWERLED.func_state_RNI2MQDZ0Z_0_cascade_\
        );

    \I__5591\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27251\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__27251\,
            I => \N__27248\
        );

    \I__5589\ : Span4Mux_v
    port map (
            O => \N__27248\,
            I => \N__27245\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__27245\,
            I => \POWERLED.dutycycle_eena_13_1_0\
        );

    \I__5587\ : InMux
    port map (
            O => \N__27242\,
            I => \N__27239\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__27239\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6\
        );

    \I__5585\ : CascadeMux
    port map (
            O => \N__27236\,
            I => \N__27232\
        );

    \I__5584\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__5583\ : InMux
    port map (
            O => \N__27232\,
            I => \N__27226\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27223\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__27226\,
            I => \N__27220\
        );

    \I__5580\ : Span4Mux_s1_h
    port map (
            O => \N__27223\,
            I => \N__27215\
        );

    \I__5579\ : Span4Mux_v
    port map (
            O => \N__27220\,
            I => \N__27215\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__5577\ : Span4Mux_v
    port map (
            O => \N__27212\,
            I => \N__27209\
        );

    \I__5576\ : Odrv4
    port map (
            O => \N__27209\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__27206\,
            I => \POWERLED.count_offZ0Z_3_cascade_\
        );

    \I__5574\ : CascadeMux
    port map (
            O => \N__27203\,
            I => \N__27199\
        );

    \I__5573\ : InMux
    port map (
            O => \N__27202\,
            I => \N__27196\
        );

    \I__5572\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27193\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__27196\,
            I => \N__27190\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__27193\,
            I => \N__27187\
        );

    \I__5569\ : Span12Mux_s5_h
    port map (
            O => \N__27190\,
            I => \N__27184\
        );

    \I__5568\ : Span12Mux_v
    port map (
            O => \N__27187\,
            I => \N__27181\
        );

    \I__5567\ : Odrv12
    port map (
            O => \N__27184\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__5566\ : Odrv12
    port map (
            O => \N__27181\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__5565\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27173\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__27173\,
            I => \N__27170\
        );

    \I__5563\ : Span4Mux_v
    port map (
            O => \N__27170\,
            I => \N__27167\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__27167\,
            I => \POWERLED.un34_clk_100khz_11\
        );

    \I__5561\ : CascadeMux
    port map (
            O => \N__27164\,
            I => \POWERLED.un34_clk_100khz_8_cascade_\
        );

    \I__5560\ : CascadeMux
    port map (
            O => \N__27161\,
            I => \POWERLED.count_off_RNI_0Z0Z_10_cascade_\
        );

    \I__5559\ : CascadeMux
    port map (
            O => \N__27158\,
            I => \POWERLED.count_off_RNI8AQHZ0Z_10_cascade_\
        );

    \I__5558\ : InMux
    port map (
            O => \N__27155\,
            I => \N__27152\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__27152\,
            I => \POWERLED.func_state_1_m2_ns_1_1\
        );

    \I__5556\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27146\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27143\
        );

    \I__5554\ : Span4Mux_v
    port map (
            O => \N__27143\,
            I => \N__27140\
        );

    \I__5553\ : Span4Mux_v
    port map (
            O => \N__27140\,
            I => \N__27137\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__27137\,
            I => \POWERLED.N_494\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__27134\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_\
        );

    \I__5550\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27128\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__27128\,
            I => \N__27125\
        );

    \I__5548\ : Span4Mux_s2_h
    port map (
            O => \N__27125\,
            I => \N__27122\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__27122\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__27119\,
            I => \POWERLED.dutycycle_1_0_iv_i_i_m2_1_6_cascade_\
        );

    \I__5545\ : InMux
    port map (
            O => \N__27116\,
            I => \N__27113\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__27113\,
            I => \N__27110\
        );

    \I__5543\ : Span4Mux_v
    port map (
            O => \N__27110\,
            I => \N__27107\
        );

    \I__5542\ : Span4Mux_h
    port map (
            O => \N__27107\,
            I => \N__27104\
        );

    \I__5541\ : Odrv4
    port map (
            O => \N__27104\,
            I => \POWERLED.N_453\
        );

    \I__5540\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27098\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27095\
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__27095\,
            I => \POWERLED.N_426_i\
        );

    \I__5537\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27089\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__27089\,
            I => \POWERLED.N_562\
        );

    \I__5535\ : CascadeMux
    port map (
            O => \N__27086\,
            I => \N__27083\
        );

    \I__5534\ : InMux
    port map (
            O => \N__27083\,
            I => \N__27079\
        );

    \I__5533\ : InMux
    port map (
            O => \N__27082\,
            I => \N__27076\
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__27079\,
            I => \N__27071\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__27076\,
            I => \N__27071\
        );

    \I__5530\ : Odrv12
    port map (
            O => \N__27071\,
            I => \POWERLED.func_state_enZ0\
        );

    \I__5529\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27065\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__27065\,
            I => \POWERLED.func_state_1_m2_1\
        );

    \I__5527\ : InMux
    port map (
            O => \N__27062\,
            I => \N__27056\
        );

    \I__5526\ : InMux
    port map (
            O => \N__27061\,
            I => \N__27056\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__27056\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__5524\ : InMux
    port map (
            O => \N__27053\,
            I => \N__27050\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__27050\,
            I => \POWERLED.count_off_0_4\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__27047\,
            I => \N__27044\
        );

    \I__5521\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27038\
        );

    \I__5520\ : InMux
    port map (
            O => \N__27043\,
            I => \N__27038\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__27038\,
            I => \N__27035\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__27035\,
            I => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\
        );

    \I__5517\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27029\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__27029\,
            I => \POWERLED.count_off_0_3\
        );

    \I__5515\ : InMux
    port map (
            O => \N__27026\,
            I => \N__27020\
        );

    \I__5514\ : InMux
    port map (
            O => \N__27025\,
            I => \N__27020\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__27020\,
            I => \N__27017\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__27017\,
            I => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\
        );

    \I__5511\ : InMux
    port map (
            O => \N__27014\,
            I => \N__27011\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__27011\,
            I => \N__27008\
        );

    \I__5509\ : Odrv4
    port map (
            O => \N__27008\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__5508\ : CascadeMux
    port map (
            O => \N__27005\,
            I => \N__27002\
        );

    \I__5507\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26998\
        );

    \I__5506\ : InMux
    port map (
            O => \N__27001\,
            I => \N__26995\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__26998\,
            I => \N__26992\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__26995\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__5503\ : Odrv4
    port map (
            O => \N__26992\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__5502\ : InMux
    port map (
            O => \N__26987\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__26984\,
            I => \N__26981\
        );

    \I__5500\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26977\
        );

    \I__5499\ : InMux
    port map (
            O => \N__26980\,
            I => \N__26974\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__26977\,
            I => \N__26971\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__26974\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__5496\ : Odrv4
    port map (
            O => \N__26971\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__5495\ : InMux
    port map (
            O => \N__26966\,
            I => \N__26960\
        );

    \I__5494\ : InMux
    port map (
            O => \N__26965\,
            I => \N__26960\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__26960\,
            I => \N__26957\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__26957\,
            I => \POWERLED.count_off_1_12\
        );

    \I__5491\ : InMux
    port map (
            O => \N__26954\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__5490\ : InMux
    port map (
            O => \N__26951\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__5489\ : InMux
    port map (
            O => \N__26948\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__5488\ : InMux
    port map (
            O => \N__26945\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__5487\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26939\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__26939\,
            I => \N__26936\
        );

    \I__5485\ : Span4Mux_v
    port map (
            O => \N__26936\,
            I => \N__26933\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__26933\,
            I => \POWERLED.N_627\
        );

    \I__5483\ : CascadeMux
    port map (
            O => \N__26930\,
            I => \N__26927\
        );

    \I__5482\ : InMux
    port map (
            O => \N__26927\,
            I => \N__26924\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__26924\,
            I => \N__26921\
        );

    \I__5480\ : Odrv12
    port map (
            O => \N__26921\,
            I => \POWERLED.N_688\
        );

    \I__5479\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26914\
        );

    \I__5478\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26911\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__26914\,
            I => \N__26908\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__26911\,
            I => \N__26904\
        );

    \I__5475\ : Span4Mux_h
    port map (
            O => \N__26908\,
            I => \N__26901\
        );

    \I__5474\ : CascadeMux
    port map (
            O => \N__26907\,
            I => \N__26898\
        );

    \I__5473\ : Span4Mux_s3_h
    port map (
            O => \N__26904\,
            I => \N__26893\
        );

    \I__5472\ : Span4Mux_v
    port map (
            O => \N__26901\,
            I => \N__26893\
        );

    \I__5471\ : InMux
    port map (
            O => \N__26898\,
            I => \N__26890\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__26893\,
            I => \POWERLED.N_74\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__26890\,
            I => \POWERLED.N_74\
        );

    \I__5468\ : CascadeMux
    port map (
            O => \N__26885\,
            I => \POWERLED.N_6_1_cascade_\
        );

    \I__5467\ : CascadeMux
    port map (
            O => \N__26882\,
            I => \POWERLED.func_state_1_m2_1_cascade_\
        );

    \I__5466\ : CascadeMux
    port map (
            O => \N__26879\,
            I => \POWERLED.func_state_cascade_\
        );

    \I__5465\ : InMux
    port map (
            O => \N__26876\,
            I => \POWERLED.un3_count_off_1_cry_1\
        );

    \I__5464\ : InMux
    port map (
            O => \N__26873\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__5463\ : InMux
    port map (
            O => \N__26870\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__5462\ : InMux
    port map (
            O => \N__26867\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__5461\ : InMux
    port map (
            O => \N__26864\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__5460\ : InMux
    port map (
            O => \N__26861\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__5459\ : InMux
    port map (
            O => \N__26858\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__5458\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26852\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__26852\,
            I => \N__26849\
        );

    \I__5456\ : Odrv4
    port map (
            O => \N__26849\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__5455\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26840\
        );

    \I__5454\ : InMux
    port map (
            O => \N__26845\,
            I => \N__26840\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__26840\,
            I => \N__26837\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__26837\,
            I => \POWERLED.count_off_1_9\
        );

    \I__5451\ : InMux
    port map (
            O => \N__26834\,
            I => \bfn_11_4_0_\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__26831\,
            I => \N__26828\
        );

    \I__5449\ : InMux
    port map (
            O => \N__26828\,
            I => \N__26824\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26821\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__26824\,
            I => \N__26818\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__26821\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__5445\ : Odrv4
    port map (
            O => \N__26818\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__5444\ : InMux
    port map (
            O => \N__26813\,
            I => \N__26807\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26812\,
            I => \N__26807\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__26807\,
            I => \N__26804\
        );

    \I__5441\ : Odrv4
    port map (
            O => \N__26804\,
            I => \POWERLED.count_off_1_10\
        );

    \I__5440\ : InMux
    port map (
            O => \N__26801\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__5439\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26794\
        );

    \I__5438\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26791\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__26794\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__26791\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__5435\ : InMux
    port map (
            O => \N__26786\,
            I => \N__26783\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__26783\,
            I => \POWERLED.count_off_0_9\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__26780\,
            I => \POWERLED.count_offZ0Z_9_cascade_\
        );

    \I__5432\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26774\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__26774\,
            I => \POWERLED.count_off_0_10\
        );

    \I__5430\ : InMux
    port map (
            O => \N__26771\,
            I => \N__26768\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__26768\,
            I => \POWERLED.count_off_0_12\
        );

    \I__5428\ : InMux
    port map (
            O => \N__26765\,
            I => \N__26758\
        );

    \I__5427\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26758\
        );

    \I__5426\ : InMux
    port map (
            O => \N__26763\,
            I => \N__26755\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__26758\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__26755\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__5423\ : InMux
    port map (
            O => \N__26750\,
            I => \N__26746\
        );

    \I__5422\ : InMux
    port map (
            O => \N__26749\,
            I => \N__26743\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__26746\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__26743\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__26738\,
            I => \POWERLED.count_clkZ0Z_7_cascade_\
        );

    \I__5418\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26732\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__26732\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3\
        );

    \I__5416\ : InMux
    port map (
            O => \N__26729\,
            I => \N__26723\
        );

    \I__5415\ : InMux
    port map (
            O => \N__26728\,
            I => \N__26723\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__26723\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__5413\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26717\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__26717\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__5411\ : InMux
    port map (
            O => \N__26714\,
            I => \N__26711\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__26711\,
            I => \N__26707\
        );

    \I__5409\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26704\
        );

    \I__5408\ : Span4Mux_h
    port map (
            O => \N__26707\,
            I => \N__26699\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__26704\,
            I => \N__26699\
        );

    \I__5406\ : Odrv4
    port map (
            O => \N__26699\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__5405\ : InMux
    port map (
            O => \N__26696\,
            I => \N__26693\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__26693\,
            I => \N__26688\
        );

    \I__5403\ : InMux
    port map (
            O => \N__26692\,
            I => \N__26685\
        );

    \I__5402\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26682\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__26688\,
            I => \N__26679\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__26685\,
            I => \POWERLED.count_clk_1_10\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__26682\,
            I => \POWERLED.count_clk_1_10\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__26679\,
            I => \POWERLED.count_clk_1_10\
        );

    \I__5397\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26669\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26665\
        );

    \I__5395\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26662\
        );

    \I__5394\ : Span4Mux_s2_v
    port map (
            O => \N__26665\,
            I => \N__26659\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26656\
        );

    \I__5392\ : Odrv4
    port map (
            O => \N__26659\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__26656\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__5390\ : CascadeMux
    port map (
            O => \N__26651\,
            I => \N__26647\
        );

    \I__5389\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26644\
        );

    \I__5388\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26641\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__26644\,
            I => \N__26638\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__26641\,
            I => \N__26635\
        );

    \I__5385\ : Odrv4
    port map (
            O => \N__26638\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__26635\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__5383\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26627\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__26627\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_0\
        );

    \I__5381\ : CascadeMux
    port map (
            O => \N__26624\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_2_cascade_\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26621\,
            I => \N__26618\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__26618\,
            I => \N__26614\
        );

    \I__5378\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26611\
        );

    \I__5377\ : Odrv4
    port map (
            O => \N__26614\,
            I => \POWERLED.count_clk_RNINSEUCZ0Z_10\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__26611\,
            I => \POWERLED.count_clk_RNINSEUCZ0Z_10\
        );

    \I__5375\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26603\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__26603\,
            I => \POWERLED.un2_count_clk_17_0_o2_1_1\
        );

    \I__5373\ : InMux
    port map (
            O => \N__26600\,
            I => \N__26594\
        );

    \I__5372\ : InMux
    port map (
            O => \N__26599\,
            I => \N__26594\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__26594\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__5370\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26582\
        );

    \I__5369\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26582\
        );

    \I__5368\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26582\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__26582\,
            I => \POWERLED.count_clk_1_12\
        );

    \I__5366\ : InMux
    port map (
            O => \N__26579\,
            I => \N__26576\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__26576\,
            I => \POWERLED.un1_count_clk_2_axb_12\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26566\
        );

    \I__5363\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26566\
        );

    \I__5362\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26563\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__26566\,
            I => \POWERLED.count_clk_1_14\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__26563\,
            I => \POWERLED.count_clk_1_14\
        );

    \I__5359\ : InMux
    port map (
            O => \N__26558\,
            I => \N__26552\
        );

    \I__5358\ : InMux
    port map (
            O => \N__26557\,
            I => \N__26552\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__26552\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__5356\ : InMux
    port map (
            O => \N__26549\,
            I => \N__26543\
        );

    \I__5355\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26543\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__26543\,
            I => \N__26539\
        );

    \I__5353\ : InMux
    port map (
            O => \N__26542\,
            I => \N__26536\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__26539\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26536\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__5350\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26524\
        );

    \I__5349\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26524\
        );

    \I__5348\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26521\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__26524\,
            I => \N__26518\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__26521\,
            I => \N__26515\
        );

    \I__5345\ : Span4Mux_s3_h
    port map (
            O => \N__26518\,
            I => \N__26510\
        );

    \I__5344\ : Span4Mux_s2_v
    port map (
            O => \N__26515\,
            I => \N__26510\
        );

    \I__5343\ : Odrv4
    port map (
            O => \N__26510\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__5342\ : InMux
    port map (
            O => \N__26507\,
            I => \N__26502\
        );

    \I__5341\ : InMux
    port map (
            O => \N__26506\,
            I => \N__26499\
        );

    \I__5340\ : InMux
    port map (
            O => \N__26505\,
            I => \N__26496\
        );

    \I__5339\ : LocalMux
    port map (
            O => \N__26502\,
            I => \N__26493\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__26499\,
            I => \N__26488\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__26496\,
            I => \N__26488\
        );

    \I__5336\ : Span4Mux_s2_v
    port map (
            O => \N__26493\,
            I => \N__26485\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__26488\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__26485\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__5333\ : CascadeMux
    port map (
            O => \N__26480\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_\
        );

    \I__5332\ : InMux
    port map (
            O => \N__26477\,
            I => \N__26472\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26476\,
            I => \N__26467\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26475\,
            I => \N__26467\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__26472\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__26467\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__5327\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26459\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__26459\,
            I => \POWERLED.N_625\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__26456\,
            I => \POWERLED.N_625_cascade_\
        );

    \I__5324\ : CascadeMux
    port map (
            O => \N__26453\,
            I => \POWERLED.count_clkZ0Z_9_cascade_\
        );

    \I__5323\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26444\
        );

    \I__5322\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26444\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__26444\,
            I => \POWERLED.count_clk_RNINSEUC_0Z0Z_10\
        );

    \I__5320\ : InMux
    port map (
            O => \N__26441\,
            I => \N__26435\
        );

    \I__5319\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26435\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__26435\,
            I => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\
        );

    \I__5317\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26429\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__26429\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__5315\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__26420\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__5312\ : InMux
    port map (
            O => \N__26417\,
            I => \N__26411\
        );

    \I__5311\ : InMux
    port map (
            O => \N__26416\,
            I => \N__26411\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__26411\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__5309\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26401\
        );

    \I__5308\ : InMux
    port map (
            O => \N__26407\,
            I => \N__26401\
        );

    \I__5307\ : InMux
    port map (
            O => \N__26406\,
            I => \N__26398\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__26401\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__26398\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__5304\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26387\
        );

    \I__5303\ : InMux
    port map (
            O => \N__26392\,
            I => \N__26387\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__26387\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__26384\,
            I => \N__26380\
        );

    \I__5300\ : InMux
    port map (
            O => \N__26383\,
            I => \N__26375\
        );

    \I__5299\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26375\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__5297\ : Odrv12
    port map (
            O => \N__26372\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26369\,
            I => \N__26366\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__26366\,
            I => \POWERLED.dutycycle_RNIHDMC5Z0Z_9\
        );

    \I__5294\ : CascadeMux
    port map (
            O => \N__26363\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__5293\ : CascadeMux
    port map (
            O => \N__26360\,
            I => \POWERLED.N_17_cascade_\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26354\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__26354\,
            I => \N__26351\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__26351\,
            I => \POWERLED.N_8_2\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26345\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__26345\,
            I => \POWERLED.G_7_i_0\
        );

    \I__5287\ : InMux
    port map (
            O => \N__26342\,
            I => \N__26339\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__26339\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \POWERLED.count_clkZ0Z_3_cascade_\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__26333\,
            I => \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_\
        );

    \I__5283\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26321\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26321\
        );

    \I__5281\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26321\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__26321\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__26318\,
            I => \POWERLED.dutycycleZ0Z_2_cascade_\
        );

    \I__5278\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__26312\,
            I => \POWERLED.g0_9_1\
        );

    \I__5276\ : InMux
    port map (
            O => \N__26309\,
            I => \N__26306\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__26306\,
            I => \POWERLED.g0_9_1_1_0\
        );

    \I__5274\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26299\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__26302\,
            I => \N__26296\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__26299\,
            I => \N__26293\
        );

    \I__5271\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26290\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__26293\,
            I => \POWERLED.dutycycle_RNIHDMC5Z0Z_10\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__26290\,
            I => \POWERLED.dutycycle_RNIHDMC5Z0Z_10\
        );

    \I__5268\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26279\
        );

    \I__5267\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26279\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__26276\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__26273\,
            I => \N__26270\
        );

    \I__5263\ : InMux
    port map (
            O => \N__26270\,
            I => \N__26264\
        );

    \I__5262\ : InMux
    port map (
            O => \N__26269\,
            I => \N__26264\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__26264\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__5260\ : InMux
    port map (
            O => \N__26261\,
            I => \N__26258\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__5258\ : Span4Mux_v
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__5257\ : Span4Mux_v
    port map (
            O => \N__26252\,
            I => \N__26249\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__26249\,
            I => \POWERLED.dutycycle_RNI6SKJ1Z0Z_9\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__26246\,
            I => \POWERLED.dutycycle_RNIHDMC5Z0Z_9_cascade_\
        );

    \I__5254\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26239\
        );

    \I__5253\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26234\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__26239\,
            I => \N__26229\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \N__26224\
        );

    \I__5250\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26221\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__26234\,
            I => \N__26218\
        );

    \I__5248\ : InMux
    port map (
            O => \N__26233\,
            I => \N__26213\
        );

    \I__5247\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26213\
        );

    \I__5246\ : Span4Mux_v
    port map (
            O => \N__26229\,
            I => \N__26210\
        );

    \I__5245\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26207\
        );

    \I__5244\ : InMux
    port map (
            O => \N__26227\,
            I => \N__26204\
        );

    \I__5243\ : InMux
    port map (
            O => \N__26224\,
            I => \N__26201\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__26221\,
            I => \N__26196\
        );

    \I__5241\ : Span4Mux_h
    port map (
            O => \N__26218\,
            I => \N__26196\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26193\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__26210\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__26207\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__26204\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__26201\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5235\ : Odrv4
    port map (
            O => \N__26196\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5234\ : Odrv12
    port map (
            O => \N__26193\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5233\ : InMux
    port map (
            O => \N__26180\,
            I => \N__26177\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__26177\,
            I => \POWERLED.un1_dutycycle_53_7_0\
        );

    \I__5231\ : CascadeMux
    port map (
            O => \N__26174\,
            I => \POWERLED.un1_dutycycle_53_41_0_cascade_\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__5229\ : InMux
    port map (
            O => \N__26168\,
            I => \N__26165\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__26165\,
            I => \N__26162\
        );

    \I__5227\ : Span4Mux_h
    port map (
            O => \N__26162\,
            I => \N__26159\
        );

    \I__5226\ : Odrv4
    port map (
            O => \N__26159\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_13\
        );

    \I__5225\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26153\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__26153\,
            I => \POWERLED.un1_dutycycle_53_59_a0_0\
        );

    \I__5223\ : CascadeMux
    port map (
            O => \N__26150\,
            I => \N__26147\
        );

    \I__5222\ : InMux
    port map (
            O => \N__26147\,
            I => \N__26141\
        );

    \I__5221\ : InMux
    port map (
            O => \N__26146\,
            I => \N__26141\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__26141\,
            I => \POWERLED.dutycycleZ1Z_11\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__26138\,
            I => \N__26134\
        );

    \I__5218\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26129\
        );

    \I__5217\ : InMux
    port map (
            O => \N__26134\,
            I => \N__26129\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__26129\,
            I => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\
        );

    \I__5215\ : CascadeMux
    port map (
            O => \N__26126\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__5214\ : CascadeMux
    port map (
            O => \N__26123\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_\
        );

    \I__5213\ : InMux
    port map (
            O => \N__26120\,
            I => \N__26116\
        );

    \I__5212\ : InMux
    port map (
            O => \N__26119\,
            I => \N__26113\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__26116\,
            I => \POWERLED.un1_dutycycle_53_56_a1_2\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__26113\,
            I => \POWERLED.un1_dutycycle_53_56_a1_2\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__5208\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26099\
        );

    \I__5206\ : Span4Mux_h
    port map (
            O => \N__26099\,
            I => \N__26096\
        );

    \I__5205\ : Odrv4
    port map (
            O => \N__26096\,
            I => \POWERLED.un1_dutycycle_53_8_2\
        );

    \I__5204\ : InMux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__26090\,
            I => \POWERLED.un1_dutycycle_53_8_0\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__26087\,
            I => \N__26084\
        );

    \I__5201\ : InMux
    port map (
            O => \N__26084\,
            I => \N__26081\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__26081\,
            I => \N__26078\
        );

    \I__5199\ : Odrv4
    port map (
            O => \N__26078\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__5198\ : CascadeMux
    port map (
            O => \N__26075\,
            I => \POWERLED.G_7_i_a5_1_1_cascade_\
        );

    \I__5197\ : InMux
    port map (
            O => \N__26072\,
            I => \N__26069\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__26069\,
            I => \POWERLED.N_11_1\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__26066\,
            I => \POWERLED.N_16_1_cascade_\
        );

    \I__5194\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__26060\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_9\
        );

    \I__5192\ : InMux
    port map (
            O => \N__26057\,
            I => \POWERLED.un1_dutycycle_94_cry_9\
        );

    \I__5191\ : InMux
    port map (
            O => \N__26054\,
            I => \POWERLED.un1_dutycycle_94_cry_10\
        );

    \I__5190\ : CascadeMux
    port map (
            O => \N__26051\,
            I => \N__26047\
        );

    \I__5189\ : InMux
    port map (
            O => \N__26050\,
            I => \N__26042\
        );

    \I__5188\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26042\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__26042\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\
        );

    \I__5186\ : InMux
    port map (
            O => \N__26039\,
            I => \POWERLED.un1_dutycycle_94_cry_11\
        );

    \I__5185\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26030\
        );

    \I__5184\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26030\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__26030\,
            I => \N__26027\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__26027\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\
        );

    \I__5181\ : InMux
    port map (
            O => \N__26024\,
            I => \POWERLED.un1_dutycycle_94_cry_12_cZ0\
        );

    \I__5180\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26012\
        );

    \I__5179\ : InMux
    port map (
            O => \N__26020\,
            I => \N__26012\
        );

    \I__5178\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26012\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__26012\,
            I => \N__26002\
        );

    \I__5176\ : InMux
    port map (
            O => \N__26011\,
            I => \N__25993\
        );

    \I__5175\ : InMux
    port map (
            O => \N__26010\,
            I => \N__25993\
        );

    \I__5174\ : InMux
    port map (
            O => \N__26009\,
            I => \N__25993\
        );

    \I__5173\ : InMux
    port map (
            O => \N__26008\,
            I => \N__25993\
        );

    \I__5172\ : CascadeMux
    port map (
            O => \N__26007\,
            I => \N__25990\
        );

    \I__5171\ : CascadeMux
    port map (
            O => \N__26006\,
            I => \N__25984\
        );

    \I__5170\ : CascadeMux
    port map (
            O => \N__26005\,
            I => \N__25980\
        );

    \I__5169\ : Span4Mux_s3_h
    port map (
            O => \N__26002\,
            I => \N__25977\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__25993\,
            I => \N__25974\
        );

    \I__5167\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25967\
        );

    \I__5166\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25967\
        );

    \I__5165\ : InMux
    port map (
            O => \N__25988\,
            I => \N__25967\
        );

    \I__5164\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25958\
        );

    \I__5163\ : InMux
    port map (
            O => \N__25984\,
            I => \N__25958\
        );

    \I__5162\ : InMux
    port map (
            O => \N__25983\,
            I => \N__25958\
        );

    \I__5161\ : InMux
    port map (
            O => \N__25980\,
            I => \N__25958\
        );

    \I__5160\ : Odrv4
    port map (
            O => \N__25977\,
            I => \POWERLED.N_435_i\
        );

    \I__5159\ : Odrv12
    port map (
            O => \N__25974\,
            I => \POWERLED.N_435_i\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__25967\,
            I => \POWERLED.N_435_i\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__25958\,
            I => \POWERLED.N_435_i\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25949\,
            I => \N__25943\
        );

    \I__5155\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25943\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__25940\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\
        );

    \I__5152\ : InMux
    port map (
            O => \N__25937\,
            I => \POWERLED.un1_dutycycle_94_cry_13\
        );

    \I__5151\ : InMux
    port map (
            O => \N__25934\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__5150\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25925\
        );

    \I__5149\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25925\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__25925\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\
        );

    \I__5147\ : CascadeMux
    port map (
            O => \N__25922\,
            I => \N__25919\
        );

    \I__5146\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25913\
        );

    \I__5145\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25913\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25910\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__25910\,
            I => \POWERLED.un1_dutycycle_53_2_1\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25901\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__25901\,
            I => \N__25896\
        );

    \I__5139\ : InMux
    port map (
            O => \N__25900\,
            I => \N__25891\
        );

    \I__5138\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25891\
        );

    \I__5137\ : Span4Mux_v
    port map (
            O => \N__25896\,
            I => \N__25888\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__25891\,
            I => \N__25885\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__25888\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_11\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__25885\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_11\
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__25880\,
            I => \N__25877\
        );

    \I__5132\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25864\
        );

    \I__5131\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25861\
        );

    \I__5130\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25856\
        );

    \I__5129\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25856\
        );

    \I__5128\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25853\
        );

    \I__5127\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25849\
        );

    \I__5126\ : InMux
    port map (
            O => \N__25871\,
            I => \N__25845\
        );

    \I__5125\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25842\
        );

    \I__5124\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25837\
        );

    \I__5123\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25837\
        );

    \I__5122\ : CascadeMux
    port map (
            O => \N__25867\,
            I => \N__25832\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__25864\,
            I => \N__25823\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__25861\,
            I => \N__25823\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__25856\,
            I => \N__25823\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__25853\,
            I => \N__25823\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25852\,
            I => \N__25819\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__25849\,
            I => \N__25816\
        );

    \I__5115\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25813\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__25845\,
            I => \N__25806\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__25842\,
            I => \N__25806\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__25837\,
            I => \N__25806\
        );

    \I__5111\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25799\
        );

    \I__5110\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25799\
        );

    \I__5109\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25799\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__25823\,
            I => \N__25796\
        );

    \I__5107\ : InMux
    port map (
            O => \N__25822\,
            I => \N__25793\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__25819\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__25816\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__25813\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__25806\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__25799\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__25796\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__25793\,
            I => \dutycycle_RNII6848_0_1\
        );

    \I__5099\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25775\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__25775\,
            I => \N__25772\
        );

    \I__5097\ : Span4Mux_h
    port map (
            O => \N__25772\,
            I => \N__25769\
        );

    \I__5096\ : Odrv4
    port map (
            O => \N__25769\,
            I => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\
        );

    \I__5095\ : InMux
    port map (
            O => \N__25766\,
            I => \POWERLED.un1_dutycycle_94_cry_0_cZ0\
        );

    \I__5094\ : InMux
    port map (
            O => \N__25763\,
            I => \POWERLED.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__5093\ : InMux
    port map (
            O => \N__25760\,
            I => \POWERLED.un1_dutycycle_94_cry_2_cZ0\
        );

    \I__5092\ : InMux
    port map (
            O => \N__25757\,
            I => \POWERLED.un1_dutycycle_94_cry_3_cZ0\
        );

    \I__5091\ : InMux
    port map (
            O => \N__25754\,
            I => \N__25751\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__25751\,
            I => \N__25748\
        );

    \I__5089\ : Span12Mux_s8_v
    port map (
            O => \N__25748\,
            I => \N__25745\
        );

    \I__5088\ : Odrv12
    port map (
            O => \N__25745\,
            I => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\
        );

    \I__5087\ : InMux
    port map (
            O => \N__25742\,
            I => \POWERLED.un1_dutycycle_94_cry_4_cZ0\
        );

    \I__5086\ : InMux
    port map (
            O => \N__25739\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__5085\ : InMux
    port map (
            O => \N__25736\,
            I => \POWERLED.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__5084\ : CascadeMux
    port map (
            O => \N__25733\,
            I => \N__25729\
        );

    \I__5083\ : InMux
    port map (
            O => \N__25732\,
            I => \N__25724\
        );

    \I__5082\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25724\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__25724\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\
        );

    \I__5080\ : InMux
    port map (
            O => \N__25721\,
            I => \bfn_9_10_0_\
        );

    \I__5079\ : InMux
    port map (
            O => \N__25718\,
            I => \POWERLED.un1_dutycycle_94_cry_8\
        );

    \I__5078\ : CascadeMux
    port map (
            O => \N__25715\,
            I => \POWERLED.g1_0_1_cascade_\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25712\,
            I => \N__25704\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25701\
        );

    \I__5075\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25696\
        );

    \I__5074\ : InMux
    port map (
            O => \N__25709\,
            I => \N__25696\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25708\,
            I => \N__25691\
        );

    \I__5072\ : InMux
    port map (
            O => \N__25707\,
            I => \N__25691\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__25704\,
            I => \N_43\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__25701\,
            I => \N_43\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__25696\,
            I => \N_43\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__25691\,
            I => \N_43\
        );

    \I__5067\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25679\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__25679\,
            I => \POWERLED.g2_1\
        );

    \I__5065\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25673\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25669\
        );

    \I__5063\ : CascadeMux
    port map (
            O => \N__25672\,
            I => \N__25666\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__25669\,
            I => \N__25659\
        );

    \I__5061\ : InMux
    port map (
            O => \N__25666\,
            I => \N__25656\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25665\,
            I => \N__25653\
        );

    \I__5059\ : InMux
    port map (
            O => \N__25664\,
            I => \N__25648\
        );

    \I__5058\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25648\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25645\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__25659\,
            I => \N__25642\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__25656\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__25653\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__25648\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__25645\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__25642\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__5050\ : InMux
    port map (
            O => \N__25631\,
            I => \N__25628\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__25628\,
            I => \N__25625\
        );

    \I__5048\ : Span4Mux_h
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__25622\,
            I => \N__25618\
        );

    \I__5046\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25615\
        );

    \I__5045\ : Odrv4
    port map (
            O => \N__25618\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__25615\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__5043\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25607\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__25607\,
            I => \N__25603\
        );

    \I__5041\ : InMux
    port map (
            O => \N__25606\,
            I => \N__25600\
        );

    \I__5040\ : Span4Mux_s2_h
    port map (
            O => \N__25603\,
            I => \N__25595\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__25600\,
            I => \N__25595\
        );

    \I__5038\ : Span4Mux_v
    port map (
            O => \N__25595\,
            I => \N__25592\
        );

    \I__5037\ : Span4Mux_h
    port map (
            O => \N__25592\,
            I => \N__25589\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__25589\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__5035\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25577\
        );

    \I__5034\ : CEMux
    port map (
            O => \N__25585\,
            I => \N__25577\
        );

    \I__5033\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25574\
        );

    \I__5032\ : CEMux
    port map (
            O => \N__25583\,
            I => \N__25567\
        );

    \I__5031\ : CEMux
    port map (
            O => \N__25582\,
            I => \N__25563\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__25577\,
            I => \N__25557\
        );

    \I__5029\ : InMux
    port map (
            O => \N__25574\,
            I => \N__25552\
        );

    \I__5028\ : CEMux
    port map (
            O => \N__25573\,
            I => \N__25552\
        );

    \I__5027\ : CascadeMux
    port map (
            O => \N__25572\,
            I => \N__25545\
        );

    \I__5026\ : InMux
    port map (
            O => \N__25571\,
            I => \N__25529\
        );

    \I__5025\ : CEMux
    port map (
            O => \N__25570\,
            I => \N__25529\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__25567\,
            I => \N__25526\
        );

    \I__5023\ : CEMux
    port map (
            O => \N__25566\,
            I => \N__25523\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__25563\,
            I => \N__25520\
        );

    \I__5021\ : CEMux
    port map (
            O => \N__25562\,
            I => \N__25517\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25512\
        );

    \I__5019\ : CEMux
    port map (
            O => \N__25560\,
            I => \N__25512\
        );

    \I__5018\ : Span4Mux_h
    port map (
            O => \N__25557\,
            I => \N__25507\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__25552\,
            I => \N__25507\
        );

    \I__5016\ : InMux
    port map (
            O => \N__25551\,
            I => \N__25498\
        );

    \I__5015\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25498\
        );

    \I__5014\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25498\
        );

    \I__5013\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25498\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25491\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25491\
        );

    \I__5010\ : InMux
    port map (
            O => \N__25543\,
            I => \N__25491\
        );

    \I__5009\ : InMux
    port map (
            O => \N__25542\,
            I => \N__25484\
        );

    \I__5008\ : InMux
    port map (
            O => \N__25541\,
            I => \N__25484\
        );

    \I__5007\ : InMux
    port map (
            O => \N__25540\,
            I => \N__25484\
        );

    \I__5006\ : InMux
    port map (
            O => \N__25539\,
            I => \N__25479\
        );

    \I__5005\ : InMux
    port map (
            O => \N__25538\,
            I => \N__25479\
        );

    \I__5004\ : InMux
    port map (
            O => \N__25537\,
            I => \N__25470\
        );

    \I__5003\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25470\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25535\,
            I => \N__25470\
        );

    \I__5001\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25470\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__25529\,
            I => \N__25464\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__25526\,
            I => \N__25461\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__25523\,
            I => \N__25452\
        );

    \I__4997\ : Span4Mux_v
    port map (
            O => \N__25520\,
            I => \N__25452\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25452\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__25512\,
            I => \N__25452\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__25507\,
            I => \N__25447\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25447\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__25491\,
            I => \N__25438\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__25484\,
            I => \N__25438\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__25479\,
            I => \N__25438\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__25470\,
            I => \N__25438\
        );

    \I__4988\ : InMux
    port map (
            O => \N__25469\,
            I => \N__25431\
        );

    \I__4987\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25431\
        );

    \I__4986\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25431\
        );

    \I__4985\ : Span12Mux_s4_h
    port map (
            O => \N__25464\,
            I => \N__25428\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__25461\,
            I => \N__25417\
        );

    \I__4983\ : Span4Mux_v
    port map (
            O => \N__25452\,
            I => \N__25417\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__25447\,
            I => \N__25417\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__25438\,
            I => \N__25417\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25417\
        );

    \I__4979\ : Odrv12
    port map (
            O => \N__25428\,
            I => \PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__25417\,
            I => \PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0\
        );

    \I__4977\ : CascadeMux
    port map (
            O => \N__25412\,
            I => \N__25396\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__25411\,
            I => \N__25393\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__25410\,
            I => \N__25387\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__25409\,
            I => \N__25381\
        );

    \I__4973\ : SRMux
    port map (
            O => \N__25408\,
            I => \N__25377\
        );

    \I__4972\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25374\
        );

    \I__4971\ : InMux
    port map (
            O => \N__25406\,
            I => \N__25368\
        );

    \I__4970\ : SRMux
    port map (
            O => \N__25405\,
            I => \N__25368\
        );

    \I__4969\ : InMux
    port map (
            O => \N__25404\,
            I => \N__25360\
        );

    \I__4968\ : SRMux
    port map (
            O => \N__25403\,
            I => \N__25360\
        );

    \I__4967\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25351\
        );

    \I__4966\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25351\
        );

    \I__4965\ : SRMux
    port map (
            O => \N__25400\,
            I => \N__25351\
        );

    \I__4964\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25351\
        );

    \I__4963\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25344\
        );

    \I__4962\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25344\
        );

    \I__4961\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25344\
        );

    \I__4960\ : SRMux
    port map (
            O => \N__25391\,
            I => \N__25335\
        );

    \I__4959\ : InMux
    port map (
            O => \N__25390\,
            I => \N__25335\
        );

    \I__4958\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25335\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25386\,
            I => \N__25335\
        );

    \I__4956\ : InMux
    port map (
            O => \N__25385\,
            I => \N__25326\
        );

    \I__4955\ : InMux
    port map (
            O => \N__25384\,
            I => \N__25326\
        );

    \I__4954\ : InMux
    port map (
            O => \N__25381\,
            I => \N__25326\
        );

    \I__4953\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25326\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__25377\,
            I => \N__25323\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__25374\,
            I => \N__25320\
        );

    \I__4950\ : SRMux
    port map (
            O => \N__25373\,
            I => \N__25316\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__25368\,
            I => \N__25313\
        );

    \I__4948\ : InMux
    port map (
            O => \N__25367\,
            I => \N__25307\
        );

    \I__4947\ : SRMux
    port map (
            O => \N__25366\,
            I => \N__25304\
        );

    \I__4946\ : SRMux
    port map (
            O => \N__25365\,
            I => \N__25301\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__25360\,
            I => \N__25284\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25284\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__25344\,
            I => \N__25284\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__25335\,
            I => \N__25284\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__25326\,
            I => \N__25284\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__25323\,
            I => \N__25281\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__25320\,
            I => \N__25278\
        );

    \I__4938\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25275\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__25316\,
            I => \N__25270\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__25313\,
            I => \N__25270\
        );

    \I__4935\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25267\
        );

    \I__4934\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25262\
        );

    \I__4933\ : InMux
    port map (
            O => \N__25310\,
            I => \N__25262\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__25307\,
            I => \N__25255\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__25304\,
            I => \N__25255\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25255\
        );

    \I__4929\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25252\
        );

    \I__4928\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25247\
        );

    \I__4927\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25247\
        );

    \I__4926\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25240\
        );

    \I__4925\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25240\
        );

    \I__4924\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25240\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__25284\,
            I => \N__25231\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__25281\,
            I => \N__25231\
        );

    \I__4921\ : Span4Mux_h
    port map (
            O => \N__25278\,
            I => \N__25231\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__25275\,
            I => \N__25231\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__25270\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__25267\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__25262\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__25255\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__25252\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__25247\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__25240\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4912\ : Odrv4
    port map (
            O => \N__25231\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__4911\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25211\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__25211\,
            I => \N__25208\
        );

    \I__4909\ : Span4Mux_v
    port map (
            O => \N__25208\,
            I => \N__25204\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__25207\,
            I => \N__25201\
        );

    \I__4907\ : Sp12to4
    port map (
            O => \N__25204\,
            I => \N__25198\
        );

    \I__4906\ : InMux
    port map (
            O => \N__25201\,
            I => \N__25195\
        );

    \I__4905\ : Odrv12
    port map (
            O => \N__25198\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__25195\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__4903\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25187\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__25187\,
            I => \N__25184\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__25184\,
            I => \N__25181\
        );

    \I__4900\ : Span4Mux_h
    port map (
            O => \N__25181\,
            I => \N__25178\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__25178\,
            I => \POWERLED.mult1_un124_sum_axb_7_l_fx\
        );

    \I__4898\ : InMux
    port map (
            O => \N__25175\,
            I => \N__25169\
        );

    \I__4897\ : InMux
    port map (
            O => \N__25174\,
            I => \N__25169\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25166\
        );

    \I__4895\ : Span4Mux_v
    port map (
            O => \N__25166\,
            I => \N__25161\
        );

    \I__4894\ : InMux
    port map (
            O => \N__25165\,
            I => \N__25158\
        );

    \I__4893\ : CascadeMux
    port map (
            O => \N__25164\,
            I => \N__25155\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__25161\,
            I => \N__25147\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__25158\,
            I => \N__25147\
        );

    \I__4890\ : InMux
    port map (
            O => \N__25155\,
            I => \N__25140\
        );

    \I__4889\ : InMux
    port map (
            O => \N__25154\,
            I => \N__25140\
        );

    \I__4888\ : InMux
    port map (
            O => \N__25153\,
            I => \N__25140\
        );

    \I__4887\ : InMux
    port map (
            O => \N__25152\,
            I => \N__25137\
        );

    \I__4886\ : Odrv4
    port map (
            O => \N__25147\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__25140\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__25137\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__4883\ : InMux
    port map (
            O => \N__25130\,
            I => \N__25127\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__4881\ : Span12Mux_s8_v
    port map (
            O => \N__25124\,
            I => \N__25121\
        );

    \I__4880\ : Odrv12
    port map (
            O => \N__25121\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__4879\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25115\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__25115\,
            I => \N__25111\
        );

    \I__4877\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25108\
        );

    \I__4876\ : Span12Mux_v
    port map (
            O => \N__25111\,
            I => \N__25101\
        );

    \I__4875\ : LocalMux
    port map (
            O => \N__25108\,
            I => \N__25101\
        );

    \I__4874\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25098\
        );

    \I__4873\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25095\
        );

    \I__4872\ : Odrv12
    port map (
            O => \N__25101\,
            I => \N_428\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__25098\,
            I => \N_428\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N_428\
        );

    \I__4869\ : IoInMux
    port map (
            O => \N__25088\,
            I => \N__25085\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__25085\,
            I => \N__25081\
        );

    \I__4867\ : IoInMux
    port map (
            O => \N__25084\,
            I => \N__25078\
        );

    \I__4866\ : IoSpan4Mux
    port map (
            O => \N__25081\,
            I => \N__25075\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__25078\,
            I => \N__25072\
        );

    \I__4864\ : IoSpan4Mux
    port map (
            O => \N__25075\,
            I => \N__25069\
        );

    \I__4863\ : Span4Mux_s2_h
    port map (
            O => \N__25072\,
            I => \N__25066\
        );

    \I__4862\ : Sp12to4
    port map (
            O => \N__25069\,
            I => \N__25063\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__25066\,
            I => \N__25060\
        );

    \I__4860\ : Odrv12
    port map (
            O => \N__25063\,
            I => pch_pwrok
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__25060\,
            I => pch_pwrok
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__25055\,
            I => \POWERLED.func_state_RNI12ASZ0Z_1_cascade_\
        );

    \I__4857\ : InMux
    port map (
            O => \N__25052\,
            I => \N__25049\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__25049\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3\
        );

    \I__4855\ : InMux
    port map (
            O => \N__25046\,
            I => \N__25043\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__25043\,
            I => \POWERLED.dutycycle_eena_13\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__25040\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3_cascade_\
        );

    \I__4852\ : InMux
    port map (
            O => \N__25037\,
            I => \N__25031\
        );

    \I__4851\ : InMux
    port map (
            O => \N__25036\,
            I => \N__25031\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__25031\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__4849\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25025\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__25025\,
            I => \POWERLED.dutycycle_RNI_13Z0Z_0\
        );

    \I__4847\ : CascadeMux
    port map (
            O => \N__25022\,
            I => \POWERLED.N_2363_0_cascade_\
        );

    \I__4846\ : InMux
    port map (
            O => \N__25019\,
            I => \N__25016\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__25016\,
            I => \POWERLED.N_12_3_0\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__25013\,
            I => \G_11_i_a10_2_1_cascade_\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__25010\,
            I => \N__25007\
        );

    \I__4842\ : InMux
    port map (
            O => \N__25007\,
            I => \N__25004\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__25004\,
            I => \N__25001\
        );

    \I__4840\ : Span4Mux_h
    port map (
            O => \N__25001\,
            I => \N__24997\
        );

    \I__4839\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24994\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__24997\,
            I => \POWERLED.g2_3\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__24994\,
            I => \POWERLED.g2_3\
        );

    \I__4836\ : InMux
    port map (
            O => \N__24989\,
            I => \N__24986\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__24986\,
            I => \N_28\
        );

    \I__4834\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__24980\,
            I => \N_7\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__24977\,
            I => \N__24973\
        );

    \I__4831\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24968\
        );

    \I__4830\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24968\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__24968\,
            I => \N__24965\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__24965\,
            I => \N_50\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__24962\,
            I => \N_7_cascade_\
        );

    \I__4826\ : InMux
    port map (
            O => \N__24959\,
            I => \N__24955\
        );

    \I__4825\ : InMux
    port map (
            O => \N__24958\,
            I => \N__24952\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__24955\,
            I => \N__24949\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__24952\,
            I => \POWERLED.N_2363_0\
        );

    \I__4822\ : Odrv4
    port map (
            O => \N__24949\,
            I => \POWERLED.N_2363_0\
        );

    \I__4821\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24941\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24941\,
            I => \N__24937\
        );

    \I__4819\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24934\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__24937\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_0\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__24934\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_0\
        );

    \I__4816\ : InMux
    port map (
            O => \N__24929\,
            I => \N__24925\
        );

    \I__4815\ : InMux
    port map (
            O => \N__24928\,
            I => \N__24918\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__24925\,
            I => \N__24915\
        );

    \I__4813\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24912\
        );

    \I__4812\ : InMux
    port map (
            O => \N__24923\,
            I => \N__24907\
        );

    \I__4811\ : InMux
    port map (
            O => \N__24922\,
            I => \N__24907\
        );

    \I__4810\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24904\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__24918\,
            I => \N__24901\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__24915\,
            I => \N__24898\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__24912\,
            I => \N__24891\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__24907\,
            I => \N__24891\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__24904\,
            I => \N__24891\
        );

    \I__4804\ : Span4Mux_s3_h
    port map (
            O => \N__24901\,
            I => \N__24884\
        );

    \I__4803\ : Span4Mux_s3_h
    port map (
            O => \N__24898\,
            I => \N__24884\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__24891\,
            I => \N__24884\
        );

    \I__4801\ : Odrv4
    port map (
            O => \N__24884\,
            I => \POWERLED.N_613\
        );

    \I__4800\ : CascadeMux
    port map (
            O => \N__24881\,
            I => \POWERLED.un1_clk_100khz_51_and_i_3_1_cascade_\
        );

    \I__4799\ : InMux
    port map (
            O => \N__24878\,
            I => \N__24874\
        );

    \I__4798\ : InMux
    port map (
            O => \N__24877\,
            I => \N__24871\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__24874\,
            I => \N__24866\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__24871\,
            I => \N__24866\
        );

    \I__4795\ : Odrv4
    port map (
            O => \N__24866\,
            I => \POWERLED.N_252_N\
        );

    \I__4794\ : CascadeMux
    port map (
            O => \N__24863\,
            I => \POWERLED.dutycycle_eena_13_1_cascade_\
        );

    \I__4793\ : CascadeMux
    port map (
            O => \N__24860\,
            I => \POWERLED.dutycycle_eena_13_cascade_\
        );

    \I__4792\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24854\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__24854\,
            I => \N__24851\
        );

    \I__4790\ : Span4Mux_h
    port map (
            O => \N__24851\,
            I => \N__24848\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__24848\,
            I => \POWERLED.N_452\
        );

    \I__4788\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24839\
        );

    \I__4787\ : InMux
    port map (
            O => \N__24844\,
            I => \N__24839\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__24839\,
            I => \N__24836\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__24836\,
            I => \POWERLED.dutycycle_set_1\
        );

    \I__4784\ : InMux
    port map (
            O => \N__24833\,
            I => \N__24830\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__24830\,
            I => \POWERLED.func_state_RNI12ASZ0Z_1\
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__24827\,
            I => \POWERLED.dutycycle_e_N_3L4_0_1_cascade_\
        );

    \I__4781\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24821\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__24821\,
            I => \POWERLED.g0_8Z0Z_0\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__24818\,
            I => \POWERLED.N_435_cascade_\
        );

    \I__4778\ : InMux
    port map (
            O => \N__24815\,
            I => \N__24812\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__4776\ : Odrv4
    port map (
            O => \N__24809\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_0\
        );

    \I__4775\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__24803\,
            I => \POWERLED.func_state_1_m2s2_i_0_0\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__24800\,
            I => \POWERLED.N_423_cascade_\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24794\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__24794\,
            I => \POWERLED.N_542\
        );

    \I__4770\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24788\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__24788\,
            I => \N__24785\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__24785\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__4767\ : InMux
    port map (
            O => \N__24782\,
            I => \N__24779\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__24779\,
            I => \POWERLED.g2\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__24776\,
            I => \N__24773\
        );

    \I__4764\ : InMux
    port map (
            O => \N__24773\,
            I => \N__24770\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__24770\,
            I => \N__24767\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__4761\ : Span4Mux_s2_h
    port map (
            O => \N__24764\,
            I => \N__24760\
        );

    \I__4760\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24757\
        );

    \I__4759\ : Odrv4
    port map (
            O => \N__24760\,
            I => \POWERLED.g0_0_5\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__24757\,
            I => \POWERLED.g0_0_5\
        );

    \I__4757\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24748\
        );

    \I__4756\ : InMux
    port map (
            O => \N__24751\,
            I => \N__24745\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__24748\,
            I => \POWERLED.g2_0\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__24745\,
            I => \POWERLED.g2_0\
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__24740\,
            I => \POWERLED.g2_cascade_\
        );

    \I__4752\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24731\
        );

    \I__4751\ : InMux
    port map (
            O => \N__24736\,
            I => \N__24731\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24728\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__24728\,
            I => \N__24725\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__24725\,
            I => \POWERLED.N_13_0_0_0\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__24722\,
            I => \POWERLED.func_stateZ0Z_0_cascade_\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24714\
        );

    \I__4745\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24709\
        );

    \I__4744\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24709\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__24714\,
            I => \N__24706\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__24709\,
            I => \N__24701\
        );

    \I__4741\ : Span4Mux_s3_v
    port map (
            O => \N__24706\,
            I => \N__24701\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__24701\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_0\
        );

    \I__4739\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24684\
        );

    \I__4738\ : IoInMux
    port map (
            O => \N__24697\,
            I => \N__24680\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__24696\,
            I => \N__24677\
        );

    \I__4736\ : InMux
    port map (
            O => \N__24695\,
            I => \N__24670\
        );

    \I__4735\ : InMux
    port map (
            O => \N__24694\,
            I => \N__24670\
        );

    \I__4734\ : InMux
    port map (
            O => \N__24693\,
            I => \N__24656\
        );

    \I__4733\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24656\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__24691\,
            I => \N__24650\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__24690\,
            I => \N__24645\
        );

    \I__4730\ : InMux
    port map (
            O => \N__24689\,
            I => \N__24632\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24632\
        );

    \I__4728\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24632\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24627\
        );

    \I__4726\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24624\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__24680\,
            I => \N__24621\
        );

    \I__4724\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24617\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__24676\,
            I => \N__24612\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24675\,
            I => \N__24608\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__24670\,
            I => \N__24605\
        );

    \I__4720\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24602\
        );

    \I__4719\ : InMux
    port map (
            O => \N__24668\,
            I => \N__24599\
        );

    \I__4718\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24596\
        );

    \I__4717\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24591\
        );

    \I__4716\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24591\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24664\,
            I => \N__24588\
        );

    \I__4714\ : InMux
    port map (
            O => \N__24663\,
            I => \N__24581\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24662\,
            I => \N__24581\
        );

    \I__4712\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24581\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__24656\,
            I => \N__24578\
        );

    \I__4710\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24565\
        );

    \I__4709\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24565\
        );

    \I__4708\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24565\
        );

    \I__4707\ : InMux
    port map (
            O => \N__24650\,
            I => \N__24565\
        );

    \I__4706\ : InMux
    port map (
            O => \N__24649\,
            I => \N__24565\
        );

    \I__4705\ : InMux
    port map (
            O => \N__24648\,
            I => \N__24565\
        );

    \I__4704\ : InMux
    port map (
            O => \N__24645\,
            I => \N__24556\
        );

    \I__4703\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24556\
        );

    \I__4702\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24556\
        );

    \I__4701\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24556\
        );

    \I__4700\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24548\
        );

    \I__4699\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24548\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24548\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24632\,
            I => \N__24545\
        );

    \I__4696\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24542\
        );

    \I__4695\ : InMux
    port map (
            O => \N__24630\,
            I => \N__24539\
        );

    \I__4694\ : Span4Mux_v
    port map (
            O => \N__24627\,
            I => \N__24534\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__24624\,
            I => \N__24534\
        );

    \I__4692\ : IoSpan4Mux
    port map (
            O => \N__24621\,
            I => \N__24531\
        );

    \I__4691\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24528\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__24617\,
            I => \N__24525\
        );

    \I__4689\ : InMux
    port map (
            O => \N__24616\,
            I => \N__24516\
        );

    \I__4688\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24516\
        );

    \I__4687\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24516\
        );

    \I__4686\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24516\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__24608\,
            I => \N__24513\
        );

    \I__4684\ : Span4Mux_s0_v
    port map (
            O => \N__24605\,
            I => \N__24510\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__24602\,
            I => \N__24507\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__24599\,
            I => \N__24502\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__24596\,
            I => \N__24499\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__24591\,
            I => \N__24486\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24486\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__24581\,
            I => \N__24486\
        );

    \I__4677\ : Span4Mux_h
    port map (
            O => \N__24578\,
            I => \N__24486\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__24565\,
            I => \N__24486\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__24556\,
            I => \N__24486\
        );

    \I__4674\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24483\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__24548\,
            I => \N__24476\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__24545\,
            I => \N__24476\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24476\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__24539\,
            I => \N__24471\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__24534\,
            I => \N__24471\
        );

    \I__4668\ : Span4Mux_s2_h
    port map (
            O => \N__24531\,
            I => \N__24466\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__24528\,
            I => \N__24466\
        );

    \I__4666\ : Span4Mux_s2_h
    port map (
            O => \N__24525\,
            I => \N__24461\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__24516\,
            I => \N__24461\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__24513\,
            I => \N__24454\
        );

    \I__4663\ : Span4Mux_v
    port map (
            O => \N__24510\,
            I => \N__24454\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__24507\,
            I => \N__24454\
        );

    \I__4661\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24449\
        );

    \I__4660\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24449\
        );

    \I__4659\ : Span12Mux_s8_v
    port map (
            O => \N__24502\,
            I => \N__24446\
        );

    \I__4658\ : Span4Mux_h
    port map (
            O => \N__24499\,
            I => \N__24439\
        );

    \I__4657\ : Span4Mux_v
    port map (
            O => \N__24486\,
            I => \N__24439\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__24483\,
            I => \N__24439\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__24476\,
            I => \N__24434\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__24471\,
            I => \N__24434\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__24466\,
            I => \N__24427\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__24461\,
            I => \N__24427\
        );

    \I__4651\ : Span4Mux_v
    port map (
            O => \N__24454\,
            I => \N__24427\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__24449\,
            I => suswarn_n
        );

    \I__4649\ : Odrv12
    port map (
            O => \N__24446\,
            I => suswarn_n
        );

    \I__4648\ : Odrv4
    port map (
            O => \N__24439\,
            I => suswarn_n
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__24434\,
            I => suswarn_n
        );

    \I__4646\ : Odrv4
    port map (
            O => \N__24427\,
            I => suswarn_n
        );

    \I__4645\ : CascadeMux
    port map (
            O => \N__24416\,
            I => \POWERLED.N_8_0_cascade_\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24410\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__24410\,
            I => \N__24407\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__24407\,
            I => \N__24404\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__24404\,
            I => \POWERLED.N_16_2\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__24401\,
            I => \POWERLED.N_423_0_cascade_\
        );

    \I__4639\ : CascadeMux
    port map (
            O => \N__24398\,
            I => \POWERLED.g1_cascade_\
        );

    \I__4638\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24392\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24392\,
            I => \POWERLED.g0_0_0\
        );

    \I__4636\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24386\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__24386\,
            I => \POWERLED.N_8_0_0\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__24383\,
            I => \POWERLED.g0_0_2_cascade_\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__24380\,
            I => \POWERLED.N_541_cascade_\
        );

    \I__4632\ : InMux
    port map (
            O => \N__24377\,
            I => \N__24373\
        );

    \I__4631\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24370\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__24373\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__24370\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__24365\,
            I => \N__24361\
        );

    \I__4627\ : InMux
    port map (
            O => \N__24364\,
            I => \N__24358\
        );

    \I__4626\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24355\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__24358\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__24355\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__4623\ : InMux
    port map (
            O => \N__24350\,
            I => \N__24346\
        );

    \I__4622\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24343\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__24346\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__24343\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24338\,
            I => \N__24335\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__4617\ : Span4Mux_h
    port map (
            O => \N__24332\,
            I => \N__24329\
        );

    \I__4616\ : Odrv4
    port map (
            O => \N__24329\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11\
        );

    \I__4615\ : CascadeMux
    port map (
            O => \N__24326\,
            I => \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\
        );

    \I__4614\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \N__24319\
        );

    \I__4613\ : InMux
    port map (
            O => \N__24322\,
            I => \N__24316\
        );

    \I__4612\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24313\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__24316\,
            I => \RSMRST_PWRGD.N_264_i\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__24313\,
            I => \RSMRST_PWRGD.N_264_i\
        );

    \I__4609\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24291\
        );

    \I__4608\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24291\
        );

    \I__4607\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24291\
        );

    \I__4606\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24291\
        );

    \I__4605\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24291\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__24303\,
            I => \N__24288\
        );

    \I__4603\ : CascadeMux
    port map (
            O => \N__24302\,
            I => \N__24285\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24280\
        );

    \I__4601\ : InMux
    port map (
            O => \N__24288\,
            I => \N__24271\
        );

    \I__4600\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24271\
        );

    \I__4599\ : InMux
    port map (
            O => \N__24284\,
            I => \N__24271\
        );

    \I__4598\ : InMux
    port map (
            O => \N__24283\,
            I => \N__24271\
        );

    \I__4597\ : Span4Mux_s0_v
    port map (
            O => \N__24280\,
            I => \N__24268\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__24271\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__24268\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__4594\ : InMux
    port map (
            O => \N__24263\,
            I => \N__24251\
        );

    \I__4593\ : InMux
    port map (
            O => \N__24262\,
            I => \N__24251\
        );

    \I__4592\ : InMux
    port map (
            O => \N__24261\,
            I => \N__24251\
        );

    \I__4591\ : InMux
    port map (
            O => \N__24260\,
            I => \N__24251\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__24251\,
            I => \N__24248\
        );

    \I__4589\ : Span4Mux_h
    port map (
            O => \N__24248\,
            I => \N__24239\
        );

    \I__4588\ : InMux
    port map (
            O => \N__24247\,
            I => \N__24226\
        );

    \I__4587\ : InMux
    port map (
            O => \N__24246\,
            I => \N__24226\
        );

    \I__4586\ : InMux
    port map (
            O => \N__24245\,
            I => \N__24226\
        );

    \I__4585\ : InMux
    port map (
            O => \N__24244\,
            I => \N__24226\
        );

    \I__4584\ : InMux
    port map (
            O => \N__24243\,
            I => \N__24226\
        );

    \I__4583\ : InMux
    port map (
            O => \N__24242\,
            I => \N__24226\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__24239\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__24226\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__4580\ : InMux
    port map (
            O => \N__24221\,
            I => \N__24214\
        );

    \I__4579\ : InMux
    port map (
            O => \N__24220\,
            I => \N__24214\
        );

    \I__4578\ : InMux
    port map (
            O => \N__24219\,
            I => \N__24211\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__24214\,
            I => \N__24208\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__24211\,
            I => \N__24205\
        );

    \I__4575\ : Span4Mux_s1_v
    port map (
            O => \N__24208\,
            I => \N__24202\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__24205\,
            I => \RSMRST_PWRGD.N_662\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__24202\,
            I => \RSMRST_PWRGD.N_662\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__24197\,
            I => \RSMRST_PWRGD.N_555_cascade_\
        );

    \I__4571\ : SRMux
    port map (
            O => \N__24194\,
            I => \N__24190\
        );

    \I__4570\ : SRMux
    port map (
            O => \N__24193\,
            I => \N__24187\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24183\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__24187\,
            I => \N__24180\
        );

    \I__4567\ : SRMux
    port map (
            O => \N__24186\,
            I => \N__24177\
        );

    \I__4566\ : Span4Mux_v
    port map (
            O => \N__24183\,
            I => \N__24170\
        );

    \I__4565\ : Span4Mux_h
    port map (
            O => \N__24180\,
            I => \N__24170\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__24177\,
            I => \N__24170\
        );

    \I__4563\ : Odrv4
    port map (
            O => \N__24170\,
            I => \RSMRST_PWRGD.G_14\
        );

    \I__4562\ : CascadeMux
    port map (
            O => \N__24167\,
            I => \N__24149\
        );

    \I__4561\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24121\
        );

    \I__4560\ : InMux
    port map (
            O => \N__24165\,
            I => \N__24121\
        );

    \I__4559\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24121\
        );

    \I__4558\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24121\
        );

    \I__4557\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24114\
        );

    \I__4556\ : InMux
    port map (
            O => \N__24161\,
            I => \N__24114\
        );

    \I__4555\ : InMux
    port map (
            O => \N__24160\,
            I => \N__24114\
        );

    \I__4554\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24105\
        );

    \I__4553\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24105\
        );

    \I__4552\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24105\
        );

    \I__4551\ : InMux
    port map (
            O => \N__24156\,
            I => \N__24105\
        );

    \I__4550\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24096\
        );

    \I__4549\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24096\
        );

    \I__4548\ : InMux
    port map (
            O => \N__24153\,
            I => \N__24096\
        );

    \I__4547\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24096\
        );

    \I__4546\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24093\
        );

    \I__4545\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24084\
        );

    \I__4544\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24084\
        );

    \I__4543\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24084\
        );

    \I__4542\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24084\
        );

    \I__4541\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24077\
        );

    \I__4540\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24077\
        );

    \I__4539\ : InMux
    port map (
            O => \N__24142\,
            I => \N__24077\
        );

    \I__4538\ : InMux
    port map (
            O => \N__24141\,
            I => \N__24068\
        );

    \I__4537\ : InMux
    port map (
            O => \N__24140\,
            I => \N__24068\
        );

    \I__4536\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24068\
        );

    \I__4535\ : InMux
    port map (
            O => \N__24138\,
            I => \N__24068\
        );

    \I__4534\ : InMux
    port map (
            O => \N__24137\,
            I => \N__24059\
        );

    \I__4533\ : InMux
    port map (
            O => \N__24136\,
            I => \N__24059\
        );

    \I__4532\ : InMux
    port map (
            O => \N__24135\,
            I => \N__24059\
        );

    \I__4531\ : InMux
    port map (
            O => \N__24134\,
            I => \N__24059\
        );

    \I__4530\ : InMux
    port map (
            O => \N__24133\,
            I => \N__24054\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24054\
        );

    \I__4528\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24049\
        );

    \I__4527\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24049\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__24121\,
            I => \N__24044\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__24114\,
            I => \N__24041\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24032\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__24096\,
            I => \N__24029\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__24093\,
            I => \N__24025\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__24022\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__24077\,
            I => \N__24019\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__24068\,
            I => \N__24016\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24013\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24010\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__24049\,
            I => \N__24007\
        );

    \I__4515\ : CEMux
    port map (
            O => \N__24048\,
            I => \N__23966\
        );

    \I__4514\ : CEMux
    port map (
            O => \N__24047\,
            I => \N__23966\
        );

    \I__4513\ : Glb2LocalMux
    port map (
            O => \N__24044\,
            I => \N__23966\
        );

    \I__4512\ : Glb2LocalMux
    port map (
            O => \N__24041\,
            I => \N__23966\
        );

    \I__4511\ : CEMux
    port map (
            O => \N__24040\,
            I => \N__23966\
        );

    \I__4510\ : CEMux
    port map (
            O => \N__24039\,
            I => \N__23966\
        );

    \I__4509\ : CEMux
    port map (
            O => \N__24038\,
            I => \N__23966\
        );

    \I__4508\ : CEMux
    port map (
            O => \N__24037\,
            I => \N__23966\
        );

    \I__4507\ : CEMux
    port map (
            O => \N__24036\,
            I => \N__23966\
        );

    \I__4506\ : CEMux
    port map (
            O => \N__24035\,
            I => \N__23966\
        );

    \I__4505\ : Glb2LocalMux
    port map (
            O => \N__24032\,
            I => \N__23966\
        );

    \I__4504\ : Glb2LocalMux
    port map (
            O => \N__24029\,
            I => \N__23966\
        );

    \I__4503\ : CEMux
    port map (
            O => \N__24028\,
            I => \N__23966\
        );

    \I__4502\ : Glb2LocalMux
    port map (
            O => \N__24025\,
            I => \N__23966\
        );

    \I__4501\ : Glb2LocalMux
    port map (
            O => \N__24022\,
            I => \N__23966\
        );

    \I__4500\ : Glb2LocalMux
    port map (
            O => \N__24019\,
            I => \N__23966\
        );

    \I__4499\ : Glb2LocalMux
    port map (
            O => \N__24016\,
            I => \N__23966\
        );

    \I__4498\ : Glb2LocalMux
    port map (
            O => \N__24013\,
            I => \N__23966\
        );

    \I__4497\ : Glb2LocalMux
    port map (
            O => \N__24010\,
            I => \N__23966\
        );

    \I__4496\ : Glb2LocalMux
    port map (
            O => \N__24007\,
            I => \N__23966\
        );

    \I__4495\ : GlobalMux
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__4494\ : gio2CtrlBuf
    port map (
            O => \N__23963\,
            I => \N_92_g\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__23960\,
            I => \RSMRST_PWRGD.G_14_cascade_\
        );

    \I__4492\ : CEMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__4490\ : Span4Mux_h
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__4489\ : Odrv4
    port map (
            O => \N__23948\,
            I => \RSMRST_PWRGD.N_92_1\
        );

    \I__4488\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23939\
        );

    \I__4487\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23939\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__23939\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__4485\ : InMux
    port map (
            O => \N__23936\,
            I => \POWERLED.un1_count_clk_2_cry_7_cZ0\
        );

    \I__4484\ : InMux
    port map (
            O => \N__23933\,
            I => \bfn_8_16_0_\
        );

    \I__4483\ : InMux
    port map (
            O => \N__23930\,
            I => \N__23927\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__4481\ : Span4Mux_s2_v
    port map (
            O => \N__23924\,
            I => \N__23921\
        );

    \I__4480\ : Odrv4
    port map (
            O => \N__23921\,
            I => \POWERLED.un1_count_clk_2_axb_10\
        );

    \I__4479\ : InMux
    port map (
            O => \N__23918\,
            I => \POWERLED.un1_count_clk_2_cry_9_cZ0\
        );

    \I__4478\ : InMux
    port map (
            O => \N__23915\,
            I => \POWERLED.un1_count_clk_2_cry_10\
        );

    \I__4477\ : InMux
    port map (
            O => \N__23912\,
            I => \POWERLED.un1_count_clk_2_cry_11\
        );

    \I__4476\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23903\
        );

    \I__4475\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23903\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__23903\,
            I => \N__23900\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__23900\,
            I => \POWERLED.count_clk_1_13\
        );

    \I__4472\ : InMux
    port map (
            O => \N__23897\,
            I => \POWERLED.un1_count_clk_2_cry_12_cZ0\
        );

    \I__4471\ : InMux
    port map (
            O => \N__23894\,
            I => \POWERLED.un1_count_clk_2_cry_13\
        );

    \I__4470\ : InMux
    port map (
            O => \N__23891\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23882\
        );

    \I__4468\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23882\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__4466\ : Odrv4
    port map (
            O => \N__23879\,
            I => \POWERLED.count_clk_1_15\
        );

    \I__4465\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23873\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__23873\,
            I => \POWERLED.un1_count_clk_2_axb_14\
        );

    \I__4463\ : InMux
    port map (
            O => \N__23870\,
            I => \N__23867\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__23867\,
            I => \N__23864\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__23864\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__4460\ : InMux
    port map (
            O => \N__23861\,
            I => \N__23855\
        );

    \I__4459\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23855\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__23855\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__4457\ : InMux
    port map (
            O => \N__23852\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__4456\ : InMux
    port map (
            O => \N__23849\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__4455\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__23843\,
            I => \N__23839\
        );

    \I__4453\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23836\
        );

    \I__4452\ : Span4Mux_h
    port map (
            O => \N__23839\,
            I => \N__23833\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__23836\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__4450\ : Odrv4
    port map (
            O => \N__23833\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__4449\ : InMux
    port map (
            O => \N__23828\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__4448\ : InMux
    port map (
            O => \N__23825\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__4447\ : InMux
    port map (
            O => \N__23822\,
            I => \N__23818\
        );

    \I__4446\ : InMux
    port map (
            O => \N__23821\,
            I => \N__23815\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__23818\,
            I => \N__23812\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__23815\,
            I => \N__23809\
        );

    \I__4443\ : Span12Mux_s7_h
    port map (
            O => \N__23812\,
            I => \N__23806\
        );

    \I__4442\ : Span4Mux_h
    port map (
            O => \N__23809\,
            I => \N__23803\
        );

    \I__4441\ : Odrv12
    port map (
            O => \N__23806\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__23803\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__4439\ : InMux
    port map (
            O => \N__23798\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__4438\ : InMux
    port map (
            O => \N__23795\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__4437\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23784\
        );

    \I__4436\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23784\
        );

    \I__4435\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23779\
        );

    \I__4434\ : InMux
    port map (
            O => \N__23789\,
            I => \N__23779\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23776\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__23779\,
            I => \N__23773\
        );

    \I__4431\ : Odrv4
    port map (
            O => \N__23776\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_6\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__23773\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_6\
        );

    \I__4429\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23765\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__23765\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_8\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23762\,
            I => \N__23756\
        );

    \I__4426\ : InMux
    port map (
            O => \N__23761\,
            I => \N__23756\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__23756\,
            I => \POWERLED.dutycycleZ1Z_14\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__23753\,
            I => \POWERLED.dutycycleZ0Z_10_cascade_\
        );

    \I__4423\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23746\
        );

    \I__4422\ : InMux
    port map (
            O => \N__23749\,
            I => \N__23743\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__23746\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_13\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__23743\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_13\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__23738\,
            I => \N__23735\
        );

    \I__4418\ : InMux
    port map (
            O => \N__23735\,
            I => \N__23732\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__23732\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_15\
        );

    \I__4416\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23726\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__23726\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__4414\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23720\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__4412\ : Span12Mux_s3_v
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__4411\ : Odrv12
    port map (
            O => \N__23714\,
            I => \POWERLED.N_492\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__23711\,
            I => \POWERLED.count_clk_en_cascade_\
        );

    \I__4409\ : InMux
    port map (
            O => \N__23708\,
            I => \N__23705\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__23705\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__4407\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23699\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__23699\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__4405\ : CascadeMux
    port map (
            O => \N__23696\,
            I => \POWERLED.dutycycle_RNI_15Z0Z_3_cascade_\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__23693\,
            I => \N__23690\
        );

    \I__4403\ : InMux
    port map (
            O => \N__23690\,
            I => \N__23687\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__23687\,
            I => \POWERLED.dutycycle_RNIZ0Z_15\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__23684\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_\
        );

    \I__4400\ : CascadeMux
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__4399\ : InMux
    port map (
            O => \N__23678\,
            I => \N__23675\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__23675\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_10\
        );

    \I__4397\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23669\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__23669\,
            I => \POWERLED.N_4_0\
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \N__23663\
        );

    \I__4394\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23660\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__23660\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_13\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__23657\,
            I => \POWERLED.un1_dutycycle_53_12_1_0_cascade_\
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__23654\,
            I => \N__23651\
        );

    \I__4390\ : InMux
    port map (
            O => \N__23651\,
            I => \N__23645\
        );

    \I__4389\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23645\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__23645\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__4387\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23636\
        );

    \I__4386\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23636\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__23633\,
            I => \POWERLED.dutycycle_RNIT70K5Z0Z_8\
        );

    \I__4383\ : CascadeMux
    port map (
            O => \N__23630\,
            I => \POWERLED.dutycycleZ0Z_3_cascade_\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_8_cascade_\
        );

    \I__4381\ : CascadeMux
    port map (
            O => \N__23624\,
            I => \POWERLED.N_6_3_cascade_\
        );

    \I__4380\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23618\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__23618\,
            I => \POWERLED.g0_9_1_0\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__23615\,
            I => \POWERLED.N_9_1_cascade_\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__23612\,
            I => \POWERLED.un1_m2_e_1_cascade_\
        );

    \I__4376\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23606\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__23606\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_8\
        );

    \I__4374\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23597\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23597\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__23597\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__4371\ : CascadeMux
    port map (
            O => \N__23594\,
            I => \POWERLED.dutycycleZ0Z_7_cascade_\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__23591\,
            I => \POWERLED.un1_dutycycle_53_56_a1_2_cascade_\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__23588\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_8_cascade_\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23582\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__23582\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_8\
        );

    \I__4366\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23576\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__23576\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_8\
        );

    \I__4364\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23567\
        );

    \I__4363\ : InMux
    port map (
            O => \N__23572\,
            I => \N__23567\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__23567\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__23564\,
            I => \N__23561\
        );

    \I__4360\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23555\
        );

    \I__4359\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23555\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__23555\,
            I => \N_16_0\
        );

    \I__4357\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23549\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23546\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__23546\,
            I => \POWERLED.g0_0_1\
        );

    \I__4354\ : CascadeMux
    port map (
            O => \N__23543\,
            I => \POWERLED.N_598_cascade_\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__23540\,
            I => \POWERLED.N_450_cascade_\
        );

    \I__4352\ : InMux
    port map (
            O => \N__23537\,
            I => \N__23534\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__23534\,
            I => \POWERLED.dutycycle_RNI5FJ65Z0Z_13\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__23531\,
            I => \N__23528\
        );

    \I__4349\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23522\
        );

    \I__4348\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23522\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__23522\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__23519\,
            I => \POWERLED.dutycycle_RNI5FJ65Z0Z_13_cascade_\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__23516\,
            I => \POWERLED.dutycycleZ0Z_11_cascade_\
        );

    \I__4344\ : InMux
    port map (
            O => \N__23513\,
            I => \N__23509\
        );

    \I__4343\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23506\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__23509\,
            I => \POWERLED.N_2336_i\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__23506\,
            I => \POWERLED.N_2336_i\
        );

    \I__4340\ : InMux
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__23498\,
            I => \POWERLED.N_449\
        );

    \I__4338\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23492\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__23492\,
            I => \G_11_i_a10_0_1\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__23489\,
            I => \N_8_3_cascade_\
        );

    \I__4335\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23483\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__23483\,
            I => \POWERLED.N_10_1\
        );

    \I__4333\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23477\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__23477\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_1\
        );

    \I__4331\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23468\
        );

    \I__4330\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23468\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__23468\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__23465\,
            I => \N__23461\
        );

    \I__4327\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23456\
        );

    \I__4326\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23456\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__23456\,
            I => \POWERLED.g0_i_o4_2\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__23453\,
            I => \POWERLED.dutycycleZ1Z_5_cascade_\
        );

    \I__4323\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23441\
        );

    \I__4322\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23441\
        );

    \I__4321\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23441\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__23441\,
            I => \POWERLED.N_546\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__23438\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__23435\,
            I => \N__23432\
        );

    \I__4317\ : InMux
    port map (
            O => \N__23432\,
            I => \N__23429\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__23429\,
            I => \N__23426\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__23426\,
            I => \POWERLED.dutycycle_RNIZ0Z_5\
        );

    \I__4314\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23417\
        );

    \I__4313\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23414\
        );

    \I__4312\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23409\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23409\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__23417\,
            I => \N__23404\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23404\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__23409\,
            I => \POWERLED.N_612\
        );

    \I__4307\ : Odrv12
    port map (
            O => \N__23404\,
            I => \POWERLED.N_612\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__23399\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_0_cascade_\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_0_cascade_\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__23393\,
            I => \POWERLED.N_676_cascade_\
        );

    \I__4303\ : CascadeMux
    port map (
            O => \N__23390\,
            I => \G_11_i_a10_0_1_cascade_\
        );

    \I__4302\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23384\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__23384\,
            I => \G_11_i_2\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__23381\,
            I => \N_9_2_cascade_\
        );

    \I__4299\ : InMux
    port map (
            O => \N__23378\,
            I => \N__23375\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__23375\,
            I => \N_8_3\
        );

    \I__4297\ : CascadeMux
    port map (
            O => \N__23372\,
            I => \POWERLED.N_413_N_cascade_\
        );

    \I__4296\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23363\
        );

    \I__4295\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23363\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__23363\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__4293\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23356\
        );

    \I__4292\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23353\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__23356\,
            I => \N__23348\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23348\
        );

    \I__4289\ : Odrv4
    port map (
            O => \N__23348\,
            I => \POWERLED.N_413_N\
        );

    \I__4288\ : CascadeMux
    port map (
            O => \N__23345\,
            I => \POWERLED.N_430_cascade_\
        );

    \I__4287\ : CascadeMux
    port map (
            O => \N__23342\,
            I => \N__23339\
        );

    \I__4286\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23333\
        );

    \I__4285\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23333\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__23333\,
            I => \POWERLED.dutycycle_eena_1\
        );

    \I__4283\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23321\
        );

    \I__4282\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23321\
        );

    \I__4281\ : InMux
    port map (
            O => \N__23328\,
            I => \N__23321\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__23321\,
            I => \SUSWARN_N_fast\
        );

    \I__4279\ : CascadeMux
    port map (
            O => \N__23318\,
            I => \N__23315\
        );

    \I__4278\ : InMux
    port map (
            O => \N__23315\,
            I => \N__23312\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__23312\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m0\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__23309\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m1_ns_1_cascade_\
        );

    \I__4275\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23303\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__23303\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m1\
        );

    \I__4273\ : CascadeMux
    port map (
            O => \N__23300\,
            I => \N__23297\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23294\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__23294\,
            I => \COUNTER.tmp_0_fast_RNI0RLUZ0Z1\
        );

    \I__4270\ : InMux
    port map (
            O => \N__23291\,
            I => \bfn_8_3_0_\
        );

    \I__4269\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23284\
        );

    \I__4268\ : InMux
    port map (
            O => \N__23287\,
            I => \N__23281\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__23284\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__23281\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__23276\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__4264\ : InMux
    port map (
            O => \N__23273\,
            I => \N__23269\
        );

    \I__4263\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__23269\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__23266\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__4260\ : InMux
    port map (
            O => \N__23261\,
            I => \bfn_8_2_0_\
        );

    \I__4259\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23254\
        );

    \I__4258\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23251\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__23254\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__23251\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__4255\ : InMux
    port map (
            O => \N__23246\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__4254\ : InMux
    port map (
            O => \N__23243\,
            I => \N__23239\
        );

    \I__4253\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__23239\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__23236\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__4250\ : InMux
    port map (
            O => \N__23231\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__4249\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23224\
        );

    \I__4248\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23221\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__23224\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__23221\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__4245\ : InMux
    port map (
            O => \N__23216\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__4244\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23209\
        );

    \I__4243\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23206\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__23209\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__23206\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__4240\ : InMux
    port map (
            O => \N__23201\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__4239\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23194\
        );

    \I__4238\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23191\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__23194\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__23191\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__4235\ : InMux
    port map (
            O => \N__23186\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__4234\ : InMux
    port map (
            O => \N__23183\,
            I => \N__23179\
        );

    \I__4233\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__23179\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__23176\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__4230\ : InMux
    port map (
            O => \N__23171\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__4229\ : CascadeMux
    port map (
            O => \N__23168\,
            I => \N__23164\
        );

    \I__4228\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23160\
        );

    \I__4227\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23155\
        );

    \I__4226\ : InMux
    port map (
            O => \N__23163\,
            I => \N__23155\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23152\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23149\
        );

    \I__4223\ : Span4Mux_h
    port map (
            O => \N__23152\,
            I => \N__23142\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__23149\,
            I => \N__23142\
        );

    \I__4221\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23139\
        );

    \I__4220\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23136\
        );

    \I__4219\ : IoSpan4Mux
    port map (
            O => \N__23142\,
            I => \N__23131\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__23139\,
            I => \N__23126\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__23136\,
            I => \N__23126\
        );

    \I__4216\ : IoInMux
    port map (
            O => \N__23135\,
            I => \N__23123\
        );

    \I__4215\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23120\
        );

    \I__4214\ : Span4Mux_s3_v
    port map (
            O => \N__23131\,
            I => \N__23115\
        );

    \I__4213\ : Span4Mux_s3_v
    port map (
            O => \N__23126\,
            I => \N__23115\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__23123\,
            I => \N__23112\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__23120\,
            I => \N__23109\
        );

    \I__4210\ : Span4Mux_v
    port map (
            O => \N__23115\,
            I => \N__23106\
        );

    \I__4209\ : Span12Mux_s4_h
    port map (
            O => \N__23112\,
            I => \N__23103\
        );

    \I__4208\ : Span4Mux_h
    port map (
            O => \N__23109\,
            I => \N__23100\
        );

    \I__4207\ : Odrv4
    port map (
            O => \N__23106\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4206\ : Odrv12
    port map (
            O => \N__23103\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__23100\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__23093\,
            I => \N__23089\
        );

    \I__4203\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23086\
        );

    \I__4202\ : InMux
    port map (
            O => \N__23089\,
            I => \N__23083\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__23086\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__23083\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__23078\,
            I => \N__23074\
        );

    \I__4198\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23071\
        );

    \I__4197\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23068\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__23071\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__23068\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__4194\ : InMux
    port map (
            O => \N__23063\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23056\
        );

    \I__4192\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23053\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__23056\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__23053\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__4189\ : InMux
    port map (
            O => \N__23048\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__4188\ : InMux
    port map (
            O => \N__23045\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__4187\ : InMux
    port map (
            O => \N__23042\,
            I => \N__23038\
        );

    \I__4186\ : InMux
    port map (
            O => \N__23041\,
            I => \N__23035\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__23038\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__23035\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__4183\ : InMux
    port map (
            O => \N__23030\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__4182\ : InMux
    port map (
            O => \N__23027\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__4181\ : InMux
    port map (
            O => \N__23024\,
            I => \N__23020\
        );

    \I__4180\ : InMux
    port map (
            O => \N__23023\,
            I => \N__23017\
        );

    \I__4179\ : LocalMux
    port map (
            O => \N__23020\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__23017\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__4177\ : InMux
    port map (
            O => \N__23012\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__4176\ : InMux
    port map (
            O => \N__23009\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__23006\,
            I => \N__23003\
        );

    \I__4174\ : InMux
    port map (
            O => \N__23003\,
            I => \N__22999\
        );

    \I__4173\ : InMux
    port map (
            O => \N__23002\,
            I => \N__22996\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__22999\,
            I => \N__22993\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__22996\,
            I => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__22993\,
            I => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\
        );

    \I__4169\ : InMux
    port map (
            O => \N__22988\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__22985\,
            I => \N__22982\
        );

    \I__4167\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22979\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__22979\,
            I => \POWERLED.mult1_un47_sum_axb_4\
        );

    \I__4165\ : CascadeMux
    port map (
            O => \N__22976\,
            I => \N__22973\
        );

    \I__4164\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22970\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__22970\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__4162\ : InMux
    port map (
            O => \N__22967\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__4161\ : CascadeMux
    port map (
            O => \N__22964\,
            I => \N__22961\
        );

    \I__4160\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22958\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__22958\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__22955\,
            I => \N__22952\
        );

    \I__4157\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22949\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__22949\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__4155\ : InMux
    port map (
            O => \N__22946\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__4154\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22940\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22937\
        );

    \I__4152\ : Odrv4
    port map (
            O => \N__22937\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_5\
        );

    \I__4151\ : InMux
    port map (
            O => \N__22934\,
            I => \N__22927\
        );

    \I__4150\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22927\
        );

    \I__4149\ : InMux
    port map (
            O => \N__22932\,
            I => \N__22924\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__22927\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__22924\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__4146\ : InMux
    port map (
            O => \N__22919\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__4144\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22910\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__22910\,
            I => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__4142\ : InMux
    port map (
            O => \N__22907\,
            I => \POWERLED.mult1_un47_sum_cry_6\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__22904\,
            I => \N__22901\
        );

    \I__4140\ : InMux
    port map (
            O => \N__22901\,
            I => \N__22893\
        );

    \I__4139\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22893\
        );

    \I__4138\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22890\
        );

    \I__4137\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22887\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__22893\,
            I => \N__22882\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__22890\,
            I => \N__22882\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__22887\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__22882\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__22877\,
            I => \N__22874\
        );

    \I__4131\ : InMux
    port map (
            O => \N__22874\,
            I => \N__22864\
        );

    \I__4130\ : InMux
    port map (
            O => \N__22873\,
            I => \N__22864\
        );

    \I__4129\ : InMux
    port map (
            O => \N__22872\,
            I => \N__22864\
        );

    \I__4128\ : InMux
    port map (
            O => \N__22871\,
            I => \N__22861\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__22864\,
            I => \N__22856\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__22861\,
            I => \N__22856\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__22856\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__4123\ : InMux
    port map (
            O => \N__22850\,
            I => \N__22847\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__22847\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__4121\ : InMux
    port map (
            O => \N__22844\,
            I => \N__22839\
        );

    \I__4120\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22836\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22833\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__22839\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__22836\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__22833\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__22826\,
            I => \N__22823\
        );

    \I__4114\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22820\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__22820\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__22817\,
            I => \N__22814\
        );

    \I__4111\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22811\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__22811\,
            I => \N__22808\
        );

    \I__4109\ : Span4Mux_s3_v
    port map (
            O => \N__22808\,
            I => \N__22805\
        );

    \I__4108\ : Odrv4
    port map (
            O => \N__22805\,
            I => \POWERLED.un1_dutycycle_53_i_28\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__22802\,
            I => \N__22798\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22794\
        );

    \I__4105\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22787\
        );

    \I__4104\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22787\
        );

    \I__4103\ : InMux
    port map (
            O => \N__22794\,
            I => \N__22787\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__22787\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__22784\,
            I => \N__22781\
        );

    \I__4100\ : InMux
    port map (
            O => \N__22781\,
            I => \N__22778\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__22778\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_14\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22772\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__22772\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__4096\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22763\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22763\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__22763\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__22760\,
            I => \N__22755\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__22759\,
            I => \N__22752\
        );

    \I__4091\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22745\
        );

    \I__4090\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22745\
        );

    \I__4089\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22745\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__22745\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__4087\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__22739\,
            I => \N__22735\
        );

    \I__4085\ : InMux
    port map (
            O => \N__22738\,
            I => \N__22732\
        );

    \I__4084\ : Span4Mux_v
    port map (
            O => \N__22735\,
            I => \N__22729\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__22732\,
            I => \N__22726\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__22729\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__22726\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__4080\ : InMux
    port map (
            O => \N__22721\,
            I => \POWERLED.un1_dutycycle_53_cry_9\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22715\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__22715\,
            I => \N__22711\
        );

    \I__4077\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22708\
        );

    \I__4076\ : Odrv4
    port map (
            O => \N__22711\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__22708\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__4074\ : InMux
    port map (
            O => \N__22703\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__4073\ : InMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__22697\,
            I => \N__22693\
        );

    \I__4071\ : InMux
    port map (
            O => \N__22696\,
            I => \N__22690\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__22693\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__22690\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__4068\ : InMux
    port map (
            O => \N__22685\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__4066\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__4065\ : LocalMux
    port map (
            O => \N__22676\,
            I => \N__22673\
        );

    \I__4064\ : Odrv4
    port map (
            O => \N__22673\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__4062\ : InMux
    port map (
            O => \N__22667\,
            I => \N__22663\
        );

    \I__4061\ : InMux
    port map (
            O => \N__22666\,
            I => \N__22660\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__22663\,
            I => \N__22657\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__22660\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__22657\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__4057\ : InMux
    port map (
            O => \N__22652\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__4056\ : InMux
    port map (
            O => \N__22649\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__4055\ : InMux
    port map (
            O => \N__22646\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__4054\ : InMux
    port map (
            O => \N__22643\,
            I => \bfn_7_13_0_\
        );

    \I__4053\ : InMux
    port map (
            O => \N__22640\,
            I => \POWERLED.CO2\
        );

    \I__4052\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22634\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__22634\,
            I => \N__22631\
        );

    \I__4050\ : Span4Mux_v
    port map (
            O => \N__22631\,
            I => \N__22628\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__22628\,
            I => \POWERLED.dutycycle_RNIZ0Z_2\
        );

    \I__4048\ : InMux
    port map (
            O => \N__22625\,
            I => \N__22622\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__22622\,
            I => \N__22618\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22621\,
            I => \N__22615\
        );

    \I__4045\ : Span12Mux_s10_v
    port map (
            O => \N__22618\,
            I => \N__22612\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__22615\,
            I => \N__22609\
        );

    \I__4043\ : Odrv12
    port map (
            O => \N__22612\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__22609\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__4041\ : InMux
    port map (
            O => \N__22604\,
            I => \POWERLED.un1_dutycycle_53_cry_1\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__4037\ : Span4Mux_v
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__22589\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_2\
        );

    \I__4035\ : InMux
    port map (
            O => \N__22586\,
            I => \N__22582\
        );

    \I__4034\ : InMux
    port map (
            O => \N__22585\,
            I => \N__22579\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__22582\,
            I => \N__22574\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__22579\,
            I => \N__22574\
        );

    \I__4031\ : Span12Mux_s6_h
    port map (
            O => \N__22574\,
            I => \N__22571\
        );

    \I__4030\ : Odrv12
    port map (
            O => \N__22571\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__4029\ : InMux
    port map (
            O => \N__22568\,
            I => \POWERLED.un1_dutycycle_53_cry_2\
        );

    \I__4028\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__4026\ : Span4Mux_v
    port map (
            O => \N__22559\,
            I => \N__22556\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__22556\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_3\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__22553\,
            I => \N__22549\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__22552\,
            I => \N__22546\
        );

    \I__4022\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22543\
        );

    \I__4021\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22540\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__22543\,
            I => \N__22537\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__22540\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_3\
        );

    \I__4018\ : Odrv4
    port map (
            O => \N__22537\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_3\
        );

    \I__4017\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22528\
        );

    \I__4016\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22525\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22522\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__22525\,
            I => \N__22519\
        );

    \I__4013\ : Span4Mux_h
    port map (
            O => \N__22522\,
            I => \N__22514\
        );

    \I__4012\ : Span4Mux_v
    port map (
            O => \N__22519\,
            I => \N__22514\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__22514\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22511\,
            I => \POWERLED.un1_dutycycle_53_cry_3\
        );

    \I__4009\ : InMux
    port map (
            O => \N__22508\,
            I => \N__22504\
        );

    \I__4008\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22501\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__22504\,
            I => \N__22498\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__22501\,
            I => \N__22495\
        );

    \I__4005\ : Odrv12
    port map (
            O => \N__22498\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__4004\ : Odrv4
    port map (
            O => \N__22495\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__4003\ : InMux
    port map (
            O => \N__22490\,
            I => \POWERLED.un1_dutycycle_53_cry_4\
        );

    \I__4002\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22483\
        );

    \I__4001\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22480\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22475\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__22480\,
            I => \N__22475\
        );

    \I__3998\ : Span4Mux_v
    port map (
            O => \N__22475\,
            I => \N__22472\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__22472\,
            I => \N__22469\
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__22469\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__3995\ : InMux
    port map (
            O => \N__22466\,
            I => \POWERLED.un1_dutycycle_53_cry_5\
        );

    \I__3994\ : InMux
    port map (
            O => \N__22463\,
            I => \N__22459\
        );

    \I__3993\ : InMux
    port map (
            O => \N__22462\,
            I => \N__22456\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22451\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22451\
        );

    \I__3990\ : Span4Mux_v
    port map (
            O => \N__22451\,
            I => \N__22448\
        );

    \I__3989\ : Span4Mux_h
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__3988\ : Odrv4
    port map (
            O => \N__22445\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__3987\ : InMux
    port map (
            O => \N__22442\,
            I => \POWERLED.un1_dutycycle_53_cry_6\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__22439\,
            I => \N__22436\
        );

    \I__3985\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22433\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__22433\,
            I => \N__22430\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__22430\,
            I => \POWERLED.dutycycle_RNIZ0Z_11\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22424\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__22424\,
            I => \N__22420\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22417\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__22420\,
            I => \N__22412\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22412\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__22412\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__3976\ : InMux
    port map (
            O => \N__22409\,
            I => \bfn_7_12_0_\
        );

    \I__3975\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__22400\,
            I => \POWERLED.dutycycle_RNIZ0Z_12\
        );

    \I__3972\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22393\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22390\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__22393\,
            I => \N__22385\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__22390\,
            I => \N__22385\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__22385\,
            I => \N__22382\
        );

    \I__3967\ : Odrv4
    port map (
            O => \N__22382\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__3966\ : InMux
    port map (
            O => \N__22379\,
            I => \POWERLED.un1_dutycycle_53_cry_8\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__22376\,
            I => \POWERLED.N_9_i_1_cascade_\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__22373\,
            I => \POWERLED.dutycycle_RNIZ0Z_8_cascade_\
        );

    \I__3963\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__22364\,
            I => \N__22361\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__22361\,
            I => \POWERLED.un1_clk_100khz_32_and_i_0_a2_0_0_0\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__22358\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_6_cascade_\
        );

    \I__3958\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22352\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__22352\,
            I => \POWERLED.un2_count_clk_17_0_0_a2_0_3\
        );

    \I__3956\ : InMux
    port map (
            O => \N__22349\,
            I => \N__22346\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__22346\,
            I => \N__22342\
        );

    \I__3954\ : InMux
    port map (
            O => \N__22345\,
            I => \N__22339\
        );

    \I__3953\ : Span4Mux_v
    port map (
            O => \N__22342\,
            I => \N__22336\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__22339\,
            I => \N__22333\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__22336\,
            I => \POWERLED.un1_dutycycle_53_axb_0\
        );

    \I__3950\ : Odrv12
    port map (
            O => \N__22333\,
            I => \POWERLED.un1_dutycycle_53_axb_0\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__22328\,
            I => \N__22325\
        );

    \I__3948\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22322\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__22322\,
            I => \N__22319\
        );

    \I__3946\ : Odrv4
    port map (
            O => \N__22319\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_0\
        );

    \I__3945\ : InMux
    port map (
            O => \N__22316\,
            I => \N__22313\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22310\
        );

    \I__3943\ : Span4Mux_v
    port map (
            O => \N__22310\,
            I => \N__22306\
        );

    \I__3942\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22303\
        );

    \I__3941\ : Span4Mux_h
    port map (
            O => \N__22306\,
            I => \N__22300\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__22303\,
            I => \N__22297\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__22300\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__22297\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3937\ : InMux
    port map (
            O => \N__22292\,
            I => \POWERLED.un1_dutycycle_53_cry_0\
        );

    \I__3936\ : InMux
    port map (
            O => \N__22289\,
            I => \N__22283\
        );

    \I__3935\ : InMux
    port map (
            O => \N__22288\,
            I => \N__22283\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__22283\,
            I => \N__22280\
        );

    \I__3933\ : Odrv12
    port map (
            O => \N__22280\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_0\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__22277\,
            I => \POWERLED.un2_count_clk_17_0_0_a2_0_4_cascade_\
        );

    \I__3931\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22270\
        );

    \I__3930\ : InMux
    port map (
            O => \N__22273\,
            I => \N__22267\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__22270\,
            I => \POWERLED.N_604\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__22267\,
            I => \POWERLED.N_604\
        );

    \I__3927\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22259\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__22259\,
            I => \POWERLED.func_state_RNI1O2V5Z0Z_1\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__22256\,
            I => \N__22253\
        );

    \I__3924\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__3922\ : Span4Mux_h
    port map (
            O => \N__22247\,
            I => \N__22244\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__22244\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__3920\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22237\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__22240\,
            I => \N__22233\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22229\
        );

    \I__3917\ : InMux
    port map (
            O => \N__22236\,
            I => \N__22226\
        );

    \I__3916\ : InMux
    port map (
            O => \N__22233\,
            I => \N__22221\
        );

    \I__3915\ : InMux
    port map (
            O => \N__22232\,
            I => \N__22221\
        );

    \I__3914\ : Span4Mux_v
    port map (
            O => \N__22229\,
            I => \N__22218\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__22226\,
            I => \N__22213\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__22221\,
            I => \N__22213\
        );

    \I__3911\ : Span4Mux_v
    port map (
            O => \N__22218\,
            I => \N__22209\
        );

    \I__3910\ : Span4Mux_v
    port map (
            O => \N__22213\,
            I => \N__22206\
        );

    \I__3909\ : InMux
    port map (
            O => \N__22212\,
            I => \N__22203\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__22209\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__22206\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__22203\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__22196\,
            I => \N__22193\
        );

    \I__3904\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__22190\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__3902\ : InMux
    port map (
            O => \N__22187\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__22184\,
            I => \N__22180\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22172\
        );

    \I__3899\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22172\
        );

    \I__3898\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22172\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__22172\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__3895\ : InMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__3893\ : Span4Mux_v
    port map (
            O => \N__22160\,
            I => \N__22157\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__22157\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__3891\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22151\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__22151\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__3889\ : InMux
    port map (
            O => \N__22148\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__3888\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22142\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__22142\,
            I => \N__22139\
        );

    \I__3886\ : Odrv12
    port map (
            O => \N__22139\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__3885\ : InMux
    port map (
            O => \N__22136\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__3884\ : InMux
    port map (
            O => \N__22133\,
            I => \N__22130\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22126\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__22129\,
            I => \N__22123\
        );

    \I__3881\ : Span4Mux_v
    port map (
            O => \N__22126\,
            I => \N__22117\
        );

    \I__3880\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22110\
        );

    \I__3879\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22110\
        );

    \I__3878\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22110\
        );

    \I__3877\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22107\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__22117\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__22110\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__22107\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__3872\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__22094\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__3870\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__22088\,
            I => \N__22085\
        );

    \I__3868\ : Odrv12
    port map (
            O => \N__22085\,
            I => \POWERLED.un1_dutycycle_53_axb_4_1\
        );

    \I__3867\ : InMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__22079\,
            I => \N__22076\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__22076\,
            I => \POWERLED.g0_7_a2_2\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__3863\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__3861\ : Span4Mux_s3_v
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__3860\ : Odrv4
    port map (
            O => \N__22061\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__3859\ : CascadeMux
    port map (
            O => \N__22058\,
            I => \POWERLED.N_672_cascade_\
        );

    \I__3858\ : InMux
    port map (
            O => \N__22055\,
            I => \N__22049\
        );

    \I__3857\ : InMux
    port map (
            O => \N__22054\,
            I => \N__22049\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__22049\,
            I => \dutycycle_RNI_1_5\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__22043\,
            I => \POWERLED_un1_dutycycle_172_m1\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__22040\,
            I => \dutycycle_RNI_3_1_cascade_\
        );

    \I__3852\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22034\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__22034\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__3850\ : InMux
    port map (
            O => \N__22031\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__3849\ : InMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__3847\ : Odrv12
    port map (
            O => \N__22022\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__3845\ : InMux
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__22013\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__3843\ : InMux
    port map (
            O => \N__22010\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__22007\,
            I => \N__22004\
        );

    \I__3841\ : InMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__3839\ : Span4Mux_v
    port map (
            O => \N__21998\,
            I => \N__21995\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__21995\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__3837\ : InMux
    port map (
            O => \N__21992\,
            I => \N__21989\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__21989\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__3835\ : InMux
    port map (
            O => \N__21986\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__3834\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21980\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21977\
        );

    \I__3832\ : Odrv12
    port map (
            O => \N__21977\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__21974\,
            I => \POWERLED.dutycycle_cascade_\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__3829\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__21965\,
            I => \POWERLED.dutycycle_1_0_0\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__21962\,
            I => \POWERLED.dutycycle_1_0_0_cascade_\
        );

    \I__3826\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21953\
        );

    \I__3825\ : InMux
    port map (
            O => \N__21958\,
            I => \N__21953\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__21953\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__21950\,
            I => \POWERLED.dutycycle_1_0_1_cascade_\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__21947\,
            I => \dutycycle_RNII6848_0_1_cascade_\
        );

    \I__3821\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__21941\,
            I => \POWERLED.dutycycle_eena_0\
        );

    \I__3819\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__21935\,
            I => \POWERLED.dutycycle_1_0_1\
        );

    \I__3817\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \POWERLED.dutycycle_eena_0_cascade_\
        );

    \I__3816\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21923\
        );

    \I__3815\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21923\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__21923\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__3813\ : CascadeMux
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__3812\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__3810\ : Span12Mux_s6_h
    port map (
            O => \N__21911\,
            I => \N__21908\
        );

    \I__3809\ : Odrv12
    port map (
            O => \N__21908\,
            I => \POWERLED.N_15\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__21905\,
            I => \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_\
        );

    \I__3807\ : InMux
    port map (
            O => \N__21902\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__3805\ : InMux
    port map (
            O => \N__21896\,
            I => \N__21887\
        );

    \I__3804\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21887\
        );

    \I__3803\ : InMux
    port map (
            O => \N__21894\,
            I => \N__21887\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__3801\ : Span12Mux_s7_v
    port map (
            O => \N__21884\,
            I => \N__21879\
        );

    \I__3800\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21876\
        );

    \I__3799\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21873\
        );

    \I__3798\ : Odrv12
    port map (
            O => \N__21879\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__21876\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__21873\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__21866\,
            I => \N__21862\
        );

    \I__3794\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21854\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21862\,
            I => \N__21854\
        );

    \I__3792\ : InMux
    port map (
            O => \N__21861\,
            I => \N__21854\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__21854\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__3790\ : InMux
    port map (
            O => \N__21851\,
            I => \N__21845\
        );

    \I__3789\ : InMux
    port map (
            O => \N__21850\,
            I => \N__21845\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__21845\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__21842\,
            I => \POWERLED.dutycycleZ0Z_0_cascade_\
        );

    \I__3786\ : CascadeMux
    port map (
            O => \N__21839\,
            I => \POWERLED.un1_dutycycle_53_axb_3_1_cascade_\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__21836\,
            I => \POWERLED.un1_dutycycle_53_axb_3_cascade_\
        );

    \I__3784\ : InMux
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__21830\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10\
        );

    \I__3782\ : CascadeMux
    port map (
            O => \N__21827\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12_cascade_\
        );

    \I__3781\ : InMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__21821\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9\
        );

    \I__3779\ : InMux
    port map (
            O => \N__21818\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__3778\ : InMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__3776\ : Span4Mux_s3_v
    port map (
            O => \N__21809\,
            I => \N__21806\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__21803\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__3773\ : InMux
    port map (
            O => \N__21800\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__3771\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__3769\ : Span4Mux_s3_v
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__3768\ : Span4Mux_v
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__21782\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21779\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__3765\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21773\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__3763\ : Span4Mux_s3_v
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__21767\,
            I => \N__21764\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__21764\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__3760\ : InMux
    port map (
            O => \N__21761\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__21758\,
            I => \N__21755\
        );

    \I__3758\ : InMux
    port map (
            O => \N__21755\,
            I => \N__21752\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__21752\,
            I => \N__21749\
        );

    \I__3756\ : Span4Mux_s3_v
    port map (
            O => \N__21749\,
            I => \N__21746\
        );

    \I__3755\ : Span4Mux_v
    port map (
            O => \N__21746\,
            I => \N__21743\
        );

    \I__3754\ : Odrv4
    port map (
            O => \N__21743\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__3753\ : InMux
    port map (
            O => \N__21740\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__3752\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21734\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__21734\,
            I => \N__21731\
        );

    \I__3750\ : Span4Mux_h
    port map (
            O => \N__21731\,
            I => \N__21728\
        );

    \I__3749\ : Span4Mux_v
    port map (
            O => \N__21728\,
            I => \N__21725\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__21725\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__21722\,
            I => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1_cascade_\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__21719\,
            I => \N__21699\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__21718\,
            I => \N__21695\
        );

    \I__3744\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21682\
        );

    \I__3743\ : InMux
    port map (
            O => \N__21716\,
            I => \N__21682\
        );

    \I__3742\ : InMux
    port map (
            O => \N__21715\,
            I => \N__21682\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21682\
        );

    \I__3740\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21682\
        );

    \I__3739\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21673\
        );

    \I__3738\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21673\
        );

    \I__3737\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21673\
        );

    \I__3736\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21673\
        );

    \I__3735\ : InMux
    port map (
            O => \N__21708\,
            I => \N__21670\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21707\,
            I => \N__21661\
        );

    \I__3733\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21661\
        );

    \I__3732\ : InMux
    port map (
            O => \N__21705\,
            I => \N__21661\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21661\
        );

    \I__3730\ : InMux
    port map (
            O => \N__21703\,
            I => \N__21652\
        );

    \I__3729\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21652\
        );

    \I__3728\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21652\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21652\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21649\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__21694\,
            I => \N__21640\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__21693\,
            I => \N__21637\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21629\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21624\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__21670\,
            I => \N__21624\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21621\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__21652\,
            I => \N__21616\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__21649\,
            I => \N__21616\
        );

    \I__3717\ : InMux
    port map (
            O => \N__21648\,
            I => \N__21613\
        );

    \I__3716\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21610\
        );

    \I__3715\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21607\
        );

    \I__3714\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21604\
        );

    \I__3713\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21593\
        );

    \I__3712\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21593\
        );

    \I__3711\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21593\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21593\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21593\
        );

    \I__3708\ : InMux
    port map (
            O => \N__21635\,
            I => \N__21584\
        );

    \I__3707\ : InMux
    port map (
            O => \N__21634\,
            I => \N__21584\
        );

    \I__3706\ : InMux
    port map (
            O => \N__21633\,
            I => \N__21584\
        );

    \I__3705\ : InMux
    port map (
            O => \N__21632\,
            I => \N__21584\
        );

    \I__3704\ : Span4Mux_s1_v
    port map (
            O => \N__21629\,
            I => \N__21577\
        );

    \I__3703\ : Span4Mux_v
    port map (
            O => \N__21624\,
            I => \N__21577\
        );

    \I__3702\ : Span4Mux_v
    port map (
            O => \N__21621\,
            I => \N__21577\
        );

    \I__3701\ : Span4Mux_h
    port map (
            O => \N__21616\,
            I => \N__21574\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__21613\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__21610\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__21607\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__21604\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__21593\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__21584\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__21577\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__21574\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__21557\,
            I => \VPP_VDDQ.N_664_cascade_\
        );

    \I__3691\ : CascadeMux
    port map (
            O => \N__21554\,
            I => \VPP_VDDQ.m4_0_0_cascade_\
        );

    \I__3690\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21533\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21524\
        );

    \I__3688\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21524\
        );

    \I__3687\ : InMux
    port map (
            O => \N__21548\,
            I => \N__21524\
        );

    \I__3686\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21524\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__21546\,
            I => \N__21519\
        );

    \I__3684\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21513\
        );

    \I__3683\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21504\
        );

    \I__3682\ : InMux
    port map (
            O => \N__21543\,
            I => \N__21504\
        );

    \I__3681\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21504\
        );

    \I__3680\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21504\
        );

    \I__3679\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21497\
        );

    \I__3678\ : InMux
    port map (
            O => \N__21539\,
            I => \N__21497\
        );

    \I__3677\ : InMux
    port map (
            O => \N__21538\,
            I => \N__21497\
        );

    \I__3676\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21492\
        );

    \I__3675\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21492\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21475\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__21524\,
            I => \N__21475\
        );

    \I__3672\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21466\
        );

    \I__3671\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21466\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21466\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21518\,
            I => \N__21466\
        );

    \I__3668\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21461\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21516\,
            I => \N__21461\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__21513\,
            I => \N__21456\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__21504\,
            I => \N__21456\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__21497\,
            I => \N__21451\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__21492\,
            I => \N__21451\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21491\,
            I => \N__21440\
        );

    \I__3661\ : InMux
    port map (
            O => \N__21490\,
            I => \N__21440\
        );

    \I__3660\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21440\
        );

    \I__3659\ : InMux
    port map (
            O => \N__21488\,
            I => \N__21440\
        );

    \I__3658\ : InMux
    port map (
            O => \N__21487\,
            I => \N__21440\
        );

    \I__3657\ : InMux
    port map (
            O => \N__21486\,
            I => \N__21429\
        );

    \I__3656\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21429\
        );

    \I__3655\ : InMux
    port map (
            O => \N__21484\,
            I => \N__21429\
        );

    \I__3654\ : InMux
    port map (
            O => \N__21483\,
            I => \N__21429\
        );

    \I__3653\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21429\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21422\
        );

    \I__3651\ : InMux
    port map (
            O => \N__21480\,
            I => \N__21419\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21414\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__21466\,
            I => \N__21414\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__21461\,
            I => \N__21409\
        );

    \I__3647\ : Span4Mux_h
    port map (
            O => \N__21456\,
            I => \N__21409\
        );

    \I__3646\ : Span4Mux_v
    port map (
            O => \N__21451\,
            I => \N__21402\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__21440\,
            I => \N__21402\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__21429\,
            I => \N__21402\
        );

    \I__3643\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21397\
        );

    \I__3642\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21397\
        );

    \I__3641\ : InMux
    port map (
            O => \N__21426\,
            I => \N__21394\
        );

    \I__3640\ : InMux
    port map (
            O => \N__21425\,
            I => \N__21391\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__21422\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__21419\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3637\ : Odrv4
    port map (
            O => \N__21414\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__21409\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__21402\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__21397\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__21394\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__21391\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__3631\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21364\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21364\
        );

    \I__3629\ : InMux
    port map (
            O => \N__21372\,
            I => \N__21364\
        );

    \I__3628\ : InMux
    port map (
            O => \N__21371\,
            I => \N__21361\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__21364\,
            I => \N__21358\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21355\
        );

    \I__3625\ : Odrv4
    port map (
            O => \N__21358\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__21355\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__21350\,
            I => \N__21345\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__21349\,
            I => \N__21341\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__21348\,
            I => \N__21338\
        );

    \I__3620\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21329\
        );

    \I__3619\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21329\
        );

    \I__3618\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21329\
        );

    \I__3617\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21322\
        );

    \I__3616\ : InMux
    port map (
            O => \N__21337\,
            I => \N__21322\
        );

    \I__3615\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21322\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21317\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__21322\,
            I => \N__21317\
        );

    \I__3612\ : Span4Mux_s1_v
    port map (
            O => \N__21317\,
            I => \N__21314\
        );

    \I__3611\ : Span4Mux_v
    port map (
            O => \N__21314\,
            I => \N__21310\
        );

    \I__3610\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21307\
        );

    \I__3609\ : Span4Mux_h
    port map (
            O => \N__21310\,
            I => \N__21301\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__21307\,
            I => \N__21301\
        );

    \I__3607\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21298\
        );

    \I__3606\ : Span4Mux_v
    port map (
            O => \N__21301\,
            I => \N__21295\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21292\
        );

    \I__3604\ : Span4Mux_v
    port map (
            O => \N__21295\,
            I => \N__21289\
        );

    \I__3603\ : Span12Mux_v
    port map (
            O => \N__21292\,
            I => \N__21286\
        );

    \I__3602\ : Sp12to4
    port map (
            O => \N__21289\,
            I => \N__21283\
        );

    \I__3601\ : Odrv12
    port map (
            O => \N__21286\,
            I => vddq_ok
        );

    \I__3600\ : Odrv12
    port map (
            O => \N__21283\,
            I => vddq_ok
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__21278\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__3598\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21269\
        );

    \I__3597\ : InMux
    port map (
            O => \N__21274\,
            I => \N__21269\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__21269\,
            I => \VPP_VDDQ.N_664\
        );

    \I__3595\ : InMux
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__21263\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__3593\ : InMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__21257\,
            I => \VPP_VDDQ.N_53\
        );

    \I__3591\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__21251\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__21248\,
            I => \N__21242\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__21247\,
            I => \N__21239\
        );

    \I__3587\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21234\
        );

    \I__3586\ : InMux
    port map (
            O => \N__21245\,
            I => \N__21231\
        );

    \I__3585\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21228\
        );

    \I__3584\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21225\
        );

    \I__3583\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21222\
        );

    \I__3582\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21219\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__21234\,
            I => \N__21216\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21203\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__21228\,
            I => \N__21200\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__21225\,
            I => \N__21196\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21193\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__21219\,
            I => \N__21190\
        );

    \I__3575\ : Glb2LocalMux
    port map (
            O => \N__21216\,
            I => \N__21155\
        );

    \I__3574\ : CEMux
    port map (
            O => \N__21215\,
            I => \N__21155\
        );

    \I__3573\ : CEMux
    port map (
            O => \N__21214\,
            I => \N__21155\
        );

    \I__3572\ : CEMux
    port map (
            O => \N__21213\,
            I => \N__21155\
        );

    \I__3571\ : CEMux
    port map (
            O => \N__21212\,
            I => \N__21155\
        );

    \I__3570\ : CEMux
    port map (
            O => \N__21211\,
            I => \N__21155\
        );

    \I__3569\ : CEMux
    port map (
            O => \N__21210\,
            I => \N__21155\
        );

    \I__3568\ : CEMux
    port map (
            O => \N__21209\,
            I => \N__21155\
        );

    \I__3567\ : CEMux
    port map (
            O => \N__21208\,
            I => \N__21155\
        );

    \I__3566\ : CEMux
    port map (
            O => \N__21207\,
            I => \N__21155\
        );

    \I__3565\ : CEMux
    port map (
            O => \N__21206\,
            I => \N__21155\
        );

    \I__3564\ : Glb2LocalMux
    port map (
            O => \N__21203\,
            I => \N__21155\
        );

    \I__3563\ : Glb2LocalMux
    port map (
            O => \N__21200\,
            I => \N__21155\
        );

    \I__3562\ : CEMux
    port map (
            O => \N__21199\,
            I => \N__21155\
        );

    \I__3561\ : Glb2LocalMux
    port map (
            O => \N__21196\,
            I => \N__21155\
        );

    \I__3560\ : Glb2LocalMux
    port map (
            O => \N__21193\,
            I => \N__21155\
        );

    \I__3559\ : Glb2LocalMux
    port map (
            O => \N__21190\,
            I => \N__21155\
        );

    \I__3558\ : GlobalMux
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__3557\ : gio2CtrlBuf
    port map (
            O => \N__21152\,
            I => \N_557_g\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__21149\,
            I => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__21146\,
            I => \N__21143\
        );

    \I__3554\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__3552\ : Odrv4
    port map (
            O => \N__21137\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__3551\ : InMux
    port map (
            O => \N__21134\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__21131\,
            I => \N__21128\
        );

    \I__3549\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__21125\,
            I => \N__21122\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__21122\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__3546\ : InMux
    port map (
            O => \N__21119\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__3545\ : InMux
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__21110\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__3542\ : InMux
    port map (
            O => \N__21107\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__3541\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__21098\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__3538\ : InMux
    port map (
            O => \N__21095\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__3537\ : InMux
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__21089\,
            I => \N__21086\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__21086\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__3534\ : InMux
    port map (
            O => \N__21083\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__3533\ : InMux
    port map (
            O => \N__21080\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__21077\,
            I => \N__21074\
        );

    \I__3531\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21071\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__21071\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__21068\,
            I => \VPP_VDDQ.N_53_cascade_\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__21065\,
            I => \N__21044\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__21064\,
            I => \N__21041\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__21063\,
            I => \N__21038\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__21062\,
            I => \N__21035\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__21061\,
            I => \N__21032\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__21060\,
            I => \N__21029\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__21059\,
            I => \N__21025\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__21058\,
            I => \N__21022\
        );

    \I__3520\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21019\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__21056\,
            I => \N__21016\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__21055\,
            I => \N__21012\
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__21054\,
            I => \N__21009\
        );

    \I__3516\ : CascadeMux
    port map (
            O => \N__21053\,
            I => \N__21005\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__21052\,
            I => \N__21001\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__21051\,
            I => \N__20994\
        );

    \I__3513\ : CascadeMux
    port map (
            O => \N__21050\,
            I => \N__20991\
        );

    \I__3512\ : CascadeMux
    port map (
            O => \N__21049\,
            I => \N__20988\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__21048\,
            I => \N__20983\
        );

    \I__3510\ : InMux
    port map (
            O => \N__21047\,
            I => \N__20970\
        );

    \I__3509\ : InMux
    port map (
            O => \N__21044\,
            I => \N__20970\
        );

    \I__3508\ : InMux
    port map (
            O => \N__21041\,
            I => \N__20970\
        );

    \I__3507\ : InMux
    port map (
            O => \N__21038\,
            I => \N__20970\
        );

    \I__3506\ : InMux
    port map (
            O => \N__21035\,
            I => \N__20970\
        );

    \I__3505\ : InMux
    port map (
            O => \N__21032\,
            I => \N__20961\
        );

    \I__3504\ : InMux
    port map (
            O => \N__21029\,
            I => \N__20961\
        );

    \I__3503\ : InMux
    port map (
            O => \N__21028\,
            I => \N__20961\
        );

    \I__3502\ : InMux
    port map (
            O => \N__21025\,
            I => \N__20961\
        );

    \I__3501\ : InMux
    port map (
            O => \N__21022\,
            I => \N__20958\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__21019\,
            I => \N__20954\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21016\,
            I => \N__20947\
        );

    \I__3498\ : InMux
    port map (
            O => \N__21015\,
            I => \N__20947\
        );

    \I__3497\ : InMux
    port map (
            O => \N__21012\,
            I => \N__20947\
        );

    \I__3496\ : InMux
    port map (
            O => \N__21009\,
            I => \N__20936\
        );

    \I__3495\ : InMux
    port map (
            O => \N__21008\,
            I => \N__20936\
        );

    \I__3494\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20936\
        );

    \I__3493\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20936\
        );

    \I__3492\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20936\
        );

    \I__3491\ : InMux
    port map (
            O => \N__21000\,
            I => \N__20927\
        );

    \I__3490\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20927\
        );

    \I__3489\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20927\
        );

    \I__3488\ : InMux
    port map (
            O => \N__20997\,
            I => \N__20927\
        );

    \I__3487\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20924\
        );

    \I__3486\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20915\
        );

    \I__3485\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20915\
        );

    \I__3484\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20915\
        );

    \I__3483\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20915\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20912\
        );

    \I__3481\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20909\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__20981\,
            I => \N__20906\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__20970\,
            I => \N__20899\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__20961\,
            I => \N__20899\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__20958\,
            I => \N__20899\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__20957\,
            I => \N__20896\
        );

    \I__3475\ : Span4Mux_h
    port map (
            O => \N__20954\,
            I => \N__20890\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__20947\,
            I => \N__20890\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20885\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__20927\,
            I => \N__20885\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__20924\,
            I => \N__20876\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__20915\,
            I => \N__20876\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__20912\,
            I => \N__20876\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20876\
        );

    \I__3467\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20873\
        );

    \I__3466\ : Span4Mux_v
    port map (
            O => \N__20899\,
            I => \N__20870\
        );

    \I__3465\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20865\
        );

    \I__3464\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20865\
        );

    \I__3463\ : Span4Mux_v
    port map (
            O => \N__20890\,
            I => \N__20858\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__20885\,
            I => \N__20858\
        );

    \I__3461\ : Span4Mux_v
    port map (
            O => \N__20876\,
            I => \N__20858\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__20873\,
            I => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1\
        );

    \I__3459\ : Odrv4
    port map (
            O => \N__20870\,
            I => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__20865\,
            I => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__20858\,
            I => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1\
        );

    \I__3456\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__20846\,
            I => \POWERLED.un79_clk_100khzlto15_3\
        );

    \I__3454\ : InMux
    port map (
            O => \N__20843\,
            I => \N__20838\
        );

    \I__3453\ : InMux
    port map (
            O => \N__20842\,
            I => \N__20835\
        );

    \I__3452\ : InMux
    port map (
            O => \N__20841\,
            I => \N__20832\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__20838\,
            I => \N__20829\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20824\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__20832\,
            I => \N__20824\
        );

    \I__3448\ : Span4Mux_v
    port map (
            O => \N__20829\,
            I => \N__20820\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__20824\,
            I => \N__20817\
        );

    \I__3446\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20814\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__20820\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__20817\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__20814\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__3442\ : InMux
    port map (
            O => \N__20807\,
            I => \N__20803\
        );

    \I__3441\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20799\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__20803\,
            I => \N__20796\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \N__20793\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20790\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__20796\,
            I => \N__20787\
        );

    \I__3436\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20784\
        );

    \I__3435\ : Odrv12
    port map (
            O => \N__20790\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__20787\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__20784\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20777\,
            I => \N__20774\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__20774\,
            I => \N__20771\
        );

    \I__3430\ : Span4Mux_s3_v
    port map (
            O => \N__20771\,
            I => \N__20768\
        );

    \I__3429\ : Span4Mux_h
    port map (
            O => \N__20768\,
            I => \N__20765\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__20765\,
            I => \POWERLED.g1_i_o4_5\
        );

    \I__3427\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20759\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__20759\,
            I => \N__20756\
        );

    \I__3425\ : Span4Mux_v
    port map (
            O => \N__20756\,
            I => \N__20751\
        );

    \I__3424\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \N__20748\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__20754\,
            I => \N__20744\
        );

    \I__3422\ : Span4Mux_v
    port map (
            O => \N__20751\,
            I => \N__20741\
        );

    \I__3421\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20736\
        );

    \I__3420\ : InMux
    port map (
            O => \N__20747\,
            I => \N__20736\
        );

    \I__3419\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20733\
        );

    \I__3418\ : Odrv4
    port map (
            O => \N__20741\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__20736\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__20733\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20720\
        );

    \I__3414\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20720\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__20720\,
            I => \POWERLED.count_1_7\
        );

    \I__3412\ : InMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__20711\,
            I => \POWERLED.count_0_7\
        );

    \I__3409\ : InMux
    port map (
            O => \N__20708\,
            I => \N__20705\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__20705\,
            I => \N__20702\
        );

    \I__3407\ : Odrv12
    port map (
            O => \N__20702\,
            I => \POWERLED.N_6\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20696\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__20696\,
            I => \N__20693\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__20693\,
            I => \N__20690\
        );

    \I__3403\ : Odrv4
    port map (
            O => \N__20690\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__3402\ : InMux
    port map (
            O => \N__20687\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__3401\ : CascadeMux
    port map (
            O => \N__20684\,
            I => \N__20681\
        );

    \I__3400\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20677\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__20680\,
            I => \N__20673\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__20677\,
            I => \N__20669\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20664\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20664\
        );

    \I__3395\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20661\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__20669\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20664\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__20661\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__20654\,
            I => \POWERLED.mult1_un61_sum_s_8_cascade_\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__20651\,
            I => \N__20647\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__20650\,
            I => \N__20643\
        );

    \I__3388\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20636\
        );

    \I__3387\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20636\
        );

    \I__3386\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20636\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__20636\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__3384\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__20630\,
            I => \N__20626\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__20629\,
            I => \N__20623\
        );

    \I__3381\ : Span4Mux_v
    port map (
            O => \N__20626\,
            I => \N__20620\
        );

    \I__3380\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20617\
        );

    \I__3379\ : Odrv4
    port map (
            O => \N__20620\,
            I => \POWERLED.mult1_un82_sum_i_8\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__20617\,
            I => \POWERLED.mult1_un82_sum_i_8\
        );

    \I__3377\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20606\
        );

    \I__3375\ : Span4Mux_h
    port map (
            O => \N__20606\,
            I => \N__20603\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__20603\,
            I => \POWERLED.count_RNICOIT_0Z0Z_12\
        );

    \I__3373\ : InMux
    port map (
            O => \N__20600\,
            I => \N__20597\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__20597\,
            I => \POWERLED.count_0_13\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__3370\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20585\
        );

    \I__3369\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20585\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__20585\,
            I => \POWERLED.count_1_13\
        );

    \I__3367\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20579\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__20579\,
            I => \N__20575\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__20578\,
            I => \N__20572\
        );

    \I__3364\ : Span4Mux_v
    port map (
            O => \N__20575\,
            I => \N__20569\
        );

    \I__3363\ : InMux
    port map (
            O => \N__20572\,
            I => \N__20566\
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__20569\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__20566\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3360\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20554\
        );

    \I__3359\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20554\
        );

    \I__3358\ : InMux
    port map (
            O => \N__20559\,
            I => \N__20551\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__20554\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__20551\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__20546\,
            I => \POWERLED.countZ0Z_13_cascade_\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__20543\,
            I => \N__20539\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__20542\,
            I => \N__20536\
        );

    \I__3352\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20527\
        );

    \I__3351\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20527\
        );

    \I__3350\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20527\
        );

    \I__3349\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20524\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__20527\,
            I => \POWERLED.count_1_12\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__20524\,
            I => \POWERLED.count_1_12\
        );

    \I__3346\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20514\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__20518\,
            I => \N__20511\
        );

    \I__3344\ : InMux
    port map (
            O => \N__20517\,
            I => \N__20508\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20505\
        );

    \I__3342\ : InMux
    port map (
            O => \N__20511\,
            I => \N__20502\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20499\
        );

    \I__3340\ : Span4Mux_v
    port map (
            O => \N__20505\,
            I => \N__20494\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__20502\,
            I => \N__20494\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__20499\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__20494\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__3336\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20486\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20480\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__20485\,
            I => \N__20477\
        );

    \I__3333\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20474\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__20483\,
            I => \N__20471\
        );

    \I__3331\ : Span4Mux_v
    port map (
            O => \N__20480\,
            I => \N__20468\
        );

    \I__3330\ : InMux
    port map (
            O => \N__20477\,
            I => \N__20465\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__20474\,
            I => \N__20462\
        );

    \I__3328\ : InMux
    port map (
            O => \N__20471\,
            I => \N__20459\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__20468\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__20465\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__20462\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__20459\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3323\ : CascadeMux
    port map (
            O => \N__20450\,
            I => \POWERLED.un79_clk_100khzlto15_3_cascade_\
        );

    \I__3322\ : InMux
    port map (
            O => \N__20447\,
            I => \N__20444\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__20444\,
            I => \N__20441\
        );

    \I__3320\ : Odrv12
    port map (
            O => \N__20441\,
            I => \POWERLED.un79_clk_100khzlto15_6\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__20438\,
            I => \N__20435\
        );

    \I__3318\ : InMux
    port map (
            O => \N__20435\,
            I => \N__20432\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__20432\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__3316\ : InMux
    port map (
            O => \N__20429\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__3315\ : InMux
    port map (
            O => \N__20426\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__20423\,
            I => \N__20418\
        );

    \I__3313\ : InMux
    port map (
            O => \N__20422\,
            I => \N__20413\
        );

    \I__3312\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20410\
        );

    \I__3311\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20405\
        );

    \I__3310\ : InMux
    port map (
            O => \N__20417\,
            I => \N__20405\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20402\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__20413\,
            I => \N__20399\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__20410\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__20405\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__20402\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__20399\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__3303\ : InMux
    port map (
            O => \N__20390\,
            I => \N__20387\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__20387\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__20384\,
            I => \N__20381\
        );

    \I__3300\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20378\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__20378\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__3298\ : InMux
    port map (
            O => \N__20375\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__3297\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20369\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__20369\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20366\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__3293\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__20357\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__3291\ : InMux
    port map (
            O => \N__20354\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__3290\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__20348\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__3288\ : InMux
    port map (
            O => \N__20345\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__20342\,
            I => \N__20339\
        );

    \I__3286\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20336\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__20336\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__3284\ : InMux
    port map (
            O => \N__20333\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__20330\,
            I => \N__20326\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__20329\,
            I => \N__20322\
        );

    \I__3281\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20315\
        );

    \I__3280\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20315\
        );

    \I__3279\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20315\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__20315\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__3277\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20309\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__20309\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__3275\ : InMux
    port map (
            O => \N__20306\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__3274\ : InMux
    port map (
            O => \N__20303\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__3273\ : CascadeMux
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__3272\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20287\
        );

    \I__3271\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20287\
        );

    \I__3270\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20287\
        );

    \I__3269\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20284\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__20287\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__20284\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__20279\,
            I => \POWERLED.mult1_un75_sum_s_8_cascade_\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__3264\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__20267\,
            I => \POWERLED.mult1_un75_sum_i_8\
        );

    \I__3261\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20261\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__20261\,
            I => \N__20258\
        );

    \I__3259\ : Odrv12
    port map (
            O => \N__20258\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__20255\,
            I => \N__20252\
        );

    \I__3257\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20249\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__20249\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__3255\ : InMux
    port map (
            O => \N__20246\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__3253\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__20237\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__3251\ : InMux
    port map (
            O => \N__20234\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__3250\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20228\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__20228\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__3248\ : InMux
    port map (
            O => \N__20225\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__3247\ : InMux
    port map (
            O => \N__20222\,
            I => \N__20219\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__20219\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__3245\ : InMux
    port map (
            O => \N__20216\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__20213\,
            I => \N__20210\
        );

    \I__3243\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__3241\ : Odrv12
    port map (
            O => \N__20204\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__3240\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20198\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__20198\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__3238\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__20192\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__3236\ : InMux
    port map (
            O => \N__20189\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__20186\,
            I => \N__20183\
        );

    \I__3234\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20180\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__20180\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__3232\ : InMux
    port map (
            O => \N__20177\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__3231\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20171\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__20171\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__3229\ : InMux
    port map (
            O => \N__20168\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__20165\,
            I => \N__20162\
        );

    \I__3227\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20159\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__20159\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__3225\ : InMux
    port map (
            O => \N__20156\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__20153\,
            I => \N__20149\
        );

    \I__3223\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20141\
        );

    \I__3222\ : InMux
    port map (
            O => \N__20149\,
            I => \N__20141\
        );

    \I__3221\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20141\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__20141\,
            I => \G_2161\
        );

    \I__3219\ : InMux
    port map (
            O => \N__20138\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__20135\,
            I => \N__20132\
        );

    \I__3217\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20129\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__20129\,
            I => \N__20126\
        );

    \I__3215\ : Span4Mux_v
    port map (
            O => \N__20126\,
            I => \N__20123\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__20123\,
            I => \POWERLED.mult1_un166_sum_i_8\
        );

    \I__3213\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20117\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__20117\,
            I => \N__20114\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__20114\,
            I => \N__20111\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__20111\,
            I => \POWERLED.mult1_un145_sum_i_8\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__20108\,
            I => \N__20105\
        );

    \I__3208\ : InMux
    port map (
            O => \N__20105\,
            I => \N__20102\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__20102\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__20099\,
            I => \N__20096\
        );

    \I__3205\ : InMux
    port map (
            O => \N__20096\,
            I => \N__20093\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20090\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__20090\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__20087\,
            I => \N__20084\
        );

    \I__3201\ : InMux
    port map (
            O => \N__20084\,
            I => \N__20081\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__20081\,
            I => \N__20078\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__20078\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__20075\,
            I => \N__20072\
        );

    \I__3197\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20069\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__20069\,
            I => \N__20066\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__20066\,
            I => \N__20063\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__20063\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20060\,
            I => \bfn_6_6_0_\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__20057\,
            I => \N__20054\
        );

    \I__3191\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20051\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__20051\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__20048\,
            I => \N__20043\
        );

    \I__3188\ : CEMux
    port map (
            O => \N__20047\,
            I => \N__20036\
        );

    \I__3187\ : CEMux
    port map (
            O => \N__20046\,
            I => \N__20031\
        );

    \I__3186\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20018\
        );

    \I__3185\ : CEMux
    port map (
            O => \N__20042\,
            I => \N__20018\
        );

    \I__3184\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20013\
        );

    \I__3183\ : CEMux
    port map (
            O => \N__20040\,
            I => \N__20013\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__20039\,
            I => \N__20010\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__20036\,
            I => \N__20005\
        );

    \I__3180\ : CEMux
    port map (
            O => \N__20035\,
            I => \N__20002\
        );

    \I__3179\ : CEMux
    port map (
            O => \N__20034\,
            I => \N__19999\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__20031\,
            I => \N__19996\
        );

    \I__3177\ : InMux
    port map (
            O => \N__20030\,
            I => \N__19989\
        );

    \I__3176\ : InMux
    port map (
            O => \N__20029\,
            I => \N__19989\
        );

    \I__3175\ : InMux
    port map (
            O => \N__20028\,
            I => \N__19989\
        );

    \I__3174\ : InMux
    port map (
            O => \N__20027\,
            I => \N__19984\
        );

    \I__3173\ : InMux
    port map (
            O => \N__20026\,
            I => \N__19984\
        );

    \I__3172\ : InMux
    port map (
            O => \N__20025\,
            I => \N__19981\
        );

    \I__3171\ : InMux
    port map (
            O => \N__20024\,
            I => \N__19974\
        );

    \I__3170\ : CEMux
    port map (
            O => \N__20023\,
            I => \N__19974\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__19971\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__20013\,
            I => \N__19968\
        );

    \I__3167\ : InMux
    port map (
            O => \N__20010\,
            I => \N__19961\
        );

    \I__3166\ : InMux
    port map (
            O => \N__20009\,
            I => \N__19961\
        );

    \I__3165\ : InMux
    port map (
            O => \N__20008\,
            I => \N__19961\
        );

    \I__3164\ : Span4Mux_v
    port map (
            O => \N__20005\,
            I => \N__19954\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__20002\,
            I => \N__19954\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__19999\,
            I => \N__19949\
        );

    \I__3161\ : Span4Mux_s0_v
    port map (
            O => \N__19996\,
            I => \N__19940\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__19989\,
            I => \N__19940\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__19984\,
            I => \N__19940\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__19981\,
            I => \N__19940\
        );

    \I__3157\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19935\
        );

    \I__3156\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19935\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19931\
        );

    \I__3154\ : Span4Mux_s2_v
    port map (
            O => \N__19971\,
            I => \N__19924\
        );

    \I__3153\ : Span4Mux_s2_v
    port map (
            O => \N__19968\,
            I => \N__19924\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__19961\,
            I => \N__19924\
        );

    \I__3151\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19919\
        );

    \I__3150\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19919\
        );

    \I__3149\ : Span4Mux_h
    port map (
            O => \N__19954\,
            I => \N__19916\
        );

    \I__3148\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19913\
        );

    \I__3147\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19910\
        );

    \I__3146\ : Span4Mux_v
    port map (
            O => \N__19949\,
            I => \N__19903\
        );

    \I__3145\ : Span4Mux_v
    port map (
            O => \N__19940\,
            I => \N__19903\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__19935\,
            I => \N__19903\
        );

    \I__3143\ : InMux
    port map (
            O => \N__19934\,
            I => \N__19900\
        );

    \I__3142\ : Span4Mux_h
    port map (
            O => \N__19931\,
            I => \N__19893\
        );

    \I__3141\ : Span4Mux_v
    port map (
            O => \N__19924\,
            I => \N__19893\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19893\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__19916\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__19913\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__19910\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__19903\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__19900\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__19893\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__19880\,
            I => \VPP_VDDQ.count_2_1_11_cascade_\
        );

    \I__3132\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__19874\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__3130\ : InMux
    port map (
            O => \N__19871\,
            I => \N__19867\
        );

    \I__3129\ : InMux
    port map (
            O => \N__19870\,
            I => \N__19864\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__19867\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__19864\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__3126\ : SRMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__19856\,
            I => \N__19853\
        );

    \I__3124\ : Span4Mux_s2_v
    port map (
            O => \N__19853\,
            I => \N__19850\
        );

    \I__3123\ : Span4Mux_h
    port map (
            O => \N__19850\,
            I => \N__19847\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__19847\,
            I => \VPP_VDDQ.N_60_i\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__19844\,
            I => \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_\
        );

    \I__3120\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19835\
        );

    \I__3119\ : InMux
    port map (
            O => \N__19840\,
            I => \N__19835\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19831\
        );

    \I__3117\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19828\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__19831\,
            I => \VPP_VDDQ.N_60\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__19828\,
            I => \VPP_VDDQ.N_60\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__19823\,
            I => \VPP_VDDQ.N_60_cascade_\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__19820\,
            I => \N__19816\
        );

    \I__3112\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19811\
        );

    \I__3111\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19811\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__19811\,
            I => \N__19808\
        );

    \I__3109\ : Odrv4
    port map (
            O => \N__19808\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__19805\,
            I => \N__19802\
        );

    \I__3107\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__19799\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__19796\,
            I => \N__19793\
        );

    \I__3104\ : InMux
    port map (
            O => \N__19793\,
            I => \N__19790\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__19790\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__3102\ : CascadeMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__3101\ : InMux
    port map (
            O => \N__19784\,
            I => \N__19781\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__19781\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__19778\,
            I => \N__19775\
        );

    \I__3098\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__19772\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__3096\ : IoInMux
    port map (
            O => \N__19769\,
            I => \N__19766\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__19766\,
            I => \N__19763\
        );

    \I__3094\ : Span4Mux_s2_h
    port map (
            O => \N__19763\,
            I => \N__19759\
        );

    \I__3093\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19756\
        );

    \I__3092\ : Sp12to4
    port map (
            O => \N__19759\,
            I => \N__19753\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__19756\,
            I => \N__19750\
        );

    \I__3090\ : Span12Mux_s11_v
    port map (
            O => \N__19753\,
            I => \N__19747\
        );

    \I__3089\ : Span12Mux_s11_v
    port map (
            O => \N__19750\,
            I => \N__19744\
        );

    \I__3088\ : Odrv12
    port map (
            O => \N__19747\,
            I => v1p8a_ok
        );

    \I__3087\ : Odrv12
    port map (
            O => \N__19744\,
            I => v1p8a_ok
        );

    \I__3086\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19736\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__19736\,
            I => \N__19733\
        );

    \I__3084\ : Span4Mux_v
    port map (
            O => \N__19733\,
            I => \N__19730\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__19730\,
            I => \N__19727\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__19727\,
            I => v5a_ok
        );

    \I__3081\ : IoInMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19717\
        );

    \I__3079\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19714\
        );

    \I__3078\ : IoSpan4Mux
    port map (
            O => \N__19717\,
            I => \N__19711\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__19714\,
            I => \N__19707\
        );

    \I__3076\ : IoSpan4Mux
    port map (
            O => \N__19711\,
            I => \N__19704\
        );

    \I__3075\ : IoInMux
    port map (
            O => \N__19710\,
            I => \N__19701\
        );

    \I__3074\ : Span4Mux_s2_v
    port map (
            O => \N__19707\,
            I => \N__19698\
        );

    \I__3073\ : IoSpan4Mux
    port map (
            O => \N__19704\,
            I => \N__19693\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19693\
        );

    \I__3071\ : Sp12to4
    port map (
            O => \N__19698\,
            I => \N__19690\
        );

    \I__3070\ : IoSpan4Mux
    port map (
            O => \N__19693\,
            I => \N__19687\
        );

    \I__3069\ : Span12Mux_s11_h
    port map (
            O => \N__19690\,
            I => \N__19684\
        );

    \I__3068\ : IoSpan4Mux
    port map (
            O => \N__19687\,
            I => \N__19681\
        );

    \I__3067\ : Span12Mux_v
    port map (
            O => \N__19684\,
            I => \N__19678\
        );

    \I__3066\ : IoSpan4Mux
    port map (
            O => \N__19681\,
            I => \N__19675\
        );

    \I__3065\ : Odrv12
    port map (
            O => \N__19678\,
            I => v33a_ok
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__19675\,
            I => v33a_ok
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__19670\,
            I => \N__19666\
        );

    \I__3062\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19661\
        );

    \I__3061\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19661\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__19658\,
            I => \N__19655\
        );

    \I__3058\ : Sp12to4
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__3057\ : Span12Mux_s8_h
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__3056\ : Odrv12
    port map (
            O => \N__19649\,
            I => slp_susn
        );

    \I__3055\ : IoInMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__3053\ : Span4Mux_s3_h
    port map (
            O => \N__19640\,
            I => \N__19637\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__3051\ : Span4Mux_v
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__19631\,
            I => v33a_enn
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__19628\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__19625\,
            I => \VPP_VDDQ.count_2_1_1_cascade_\
        );

    \I__3047\ : InMux
    port map (
            O => \N__19622\,
            I => \N__19618\
        );

    \I__3046\ : InMux
    port map (
            O => \N__19621\,
            I => \N__19615\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__19618\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__19615\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__3043\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19607\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__19607\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__19604\,
            I => \N__19600\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__19603\,
            I => \N__19596\
        );

    \I__3039\ : InMux
    port map (
            O => \N__19600\,
            I => \N__19592\
        );

    \I__3038\ : InMux
    port map (
            O => \N__19599\,
            I => \N__19589\
        );

    \I__3037\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19584\
        );

    \I__3036\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19584\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__19592\,
            I => \N__19581\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__19589\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__19584\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__19581\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__3031\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19571\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__19571\,
            I => \VPP_VDDQ.un9_clk_100khz_1\
        );

    \I__3029\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19565\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__19565\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1\
        );

    \I__3027\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19556\
        );

    \I__3026\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19556\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__19556\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__3024\ : InMux
    port map (
            O => \N__19553\,
            I => \N__19547\
        );

    \I__3023\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19547\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19547\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__3021\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19538\
        );

    \I__3020\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19538\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__19538\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__19535\,
            I => \VPP_VDDQ_delayed_vddq_ok_cascade_\
        );

    \I__3017\ : IoInMux
    port map (
            O => \N__19532\,
            I => \N__19529\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__19529\,
            I => vccst_pwrgd
        );

    \I__3015\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__19523\,
            I => \N__19519\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19522\,
            I => \N__19516\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__19519\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__19516\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__3010\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__19508\,
            I => \VPP_VDDQ.un9_clk_100khz_9\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__19505\,
            I => \VPP_VDDQ.un9_clk_100khz_0_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19499\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__19496\,
            I => \VPP_VDDQ.un9_clk_100khz_13\
        );

    \I__3004\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19487\
        );

    \I__3003\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19487\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__19487\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__19484\,
            I => \VPP_VDDQ.N_1_i_cascade_\
        );

    \I__3000\ : InMux
    port map (
            O => \N__19481\,
            I => \N__19478\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__19478\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__19475\,
            I => \VPP_VDDQ.count_2_1_6_cascade_\
        );

    \I__2997\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19466\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19466\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__19466\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__2994\ : InMux
    port map (
            O => \N__19463\,
            I => \N__19460\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__19460\,
            I => \VPP_VDDQ.un1_count_2_1_axb_6\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__19457\,
            I => \N__19453\
        );

    \I__2991\ : InMux
    port map (
            O => \N__19456\,
            I => \N__19448\
        );

    \I__2990\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19448\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__19448\,
            I => \POWERLED.count_1_9\
        );

    \I__2988\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19442\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__19442\,
            I => \POWERLED.count_0_9\
        );

    \I__2986\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19436\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__19436\,
            I => \N__19431\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19428\
        );

    \I__2983\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19425\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__19431\,
            I => \POWERLED.count_1_10\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__19428\,
            I => \POWERLED.count_1_10\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__19425\,
            I => \POWERLED.count_1_10\
        );

    \I__2979\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__19415\,
            I => \POWERLED.count_0_10\
        );

    \I__2977\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19407\
        );

    \I__2976\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19404\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__19410\,
            I => \N__19401\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19398\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19395\
        );

    \I__2972\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19392\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__19398\,
            I => \N__19389\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__19395\,
            I => \N__19384\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__19392\,
            I => \N__19384\
        );

    \I__2968\ : Odrv4
    port map (
            O => \N__19389\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__19384\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2966\ : InMux
    port map (
            O => \N__19379\,
            I => \N__19374\
        );

    \I__2965\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19369\
        );

    \I__2964\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19369\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__19374\,
            I => \N__19366\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__2961\ : Odrv12
    port map (
            O => \N__19366\,
            I => \POWERLED.count_1_6\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__19363\,
            I => \POWERLED.count_1_6\
        );

    \I__2959\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19355\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__19355\,
            I => \POWERLED.count_0_6\
        );

    \I__2957\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19349\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__19349\,
            I => \N__19344\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19341\
        );

    \I__2954\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19338\
        );

    \I__2953\ : Span4Mux_s3_v
    port map (
            O => \N__19344\,
            I => \N__19335\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__19341\,
            I => \N__19330\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__19338\,
            I => \N__19330\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__19335\,
            I => \POWERLED.count_1_8\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__19330\,
            I => \POWERLED.count_1_8\
        );

    \I__2948\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__19319\,
            I => \POWERLED.count_0_8\
        );

    \I__2945\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19312\
        );

    \I__2944\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19309\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__19312\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__19309\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__2941\ : InMux
    port map (
            O => \N__19304\,
            I => \N__19301\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__19301\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__19298\,
            I => \VPP_VDDQ.count_2_1_3_cascade_\
        );

    \I__2938\ : InMux
    port map (
            O => \N__19295\,
            I => \N__19291\
        );

    \I__2937\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__19291\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__19288\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__2934\ : InMux
    port map (
            O => \N__19283\,
            I => \bfn_5_14_0_\
        );

    \I__2933\ : InMux
    port map (
            O => \N__19280\,
            I => \N__19277\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__19277\,
            I => \N__19273\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__19276\,
            I => \N__19269\
        );

    \I__2930\ : Span4Mux_v
    port map (
            O => \N__19273\,
            I => \N__19266\
        );

    \I__2929\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19263\
        );

    \I__2928\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19260\
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__19266\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__19263\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__19260\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__2924\ : InMux
    port map (
            O => \N__19253\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__2923\ : InMux
    port map (
            O => \N__19250\,
            I => \N__19246\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__19249\,
            I => \N__19242\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__19246\,
            I => \N__19239\
        );

    \I__2920\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19236\
        );

    \I__2919\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19233\
        );

    \I__2918\ : Odrv12
    port map (
            O => \N__19239\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__19236\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__19233\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__2915\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19222\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__19225\,
            I => \N__19219\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__19222\,
            I => \N__19215\
        );

    \I__2912\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19210\
        );

    \I__2911\ : InMux
    port map (
            O => \N__19218\,
            I => \N__19210\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__19215\,
            I => \POWERLED.count_1_11\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__19210\,
            I => \POWERLED.count_1_11\
        );

    \I__2908\ : InMux
    port map (
            O => \N__19205\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__2907\ : InMux
    port map (
            O => \N__19202\,
            I => \POWERLED.un1_count_cry_11\
        );

    \I__2906\ : InMux
    port map (
            O => \N__19199\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__19196\,
            I => \N__19193\
        );

    \I__2904\ : InMux
    port map (
            O => \N__19193\,
            I => \N__19187\
        );

    \I__2903\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19187\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__19187\,
            I => \POWERLED.count_1_14\
        );

    \I__2901\ : InMux
    port map (
            O => \N__19184\,
            I => \POWERLED.un1_count_cry_13\
        );

    \I__2900\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19176\
        );

    \I__2899\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19167\
        );

    \I__2898\ : InMux
    port map (
            O => \N__19179\,
            I => \N__19167\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__19176\,
            I => \N__19164\
        );

    \I__2896\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19151\
        );

    \I__2895\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19151\
        );

    \I__2894\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19151\
        );

    \I__2893\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19151\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__19167\,
            I => \N__19148\
        );

    \I__2891\ : Span4Mux_v
    port map (
            O => \N__19164\,
            I => \N__19138\
        );

    \I__2890\ : InMux
    port map (
            O => \N__19163\,
            I => \N__19131\
        );

    \I__2889\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19131\
        );

    \I__2888\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19131\
        );

    \I__2887\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19128\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19123\
        );

    \I__2885\ : Span4Mux_v
    port map (
            O => \N__19148\,
            I => \N__19123\
        );

    \I__2884\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19114\
        );

    \I__2883\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19114\
        );

    \I__2882\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19114\
        );

    \I__2881\ : InMux
    port map (
            O => \N__19144\,
            I => \N__19114\
        );

    \I__2880\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19107\
        );

    \I__2879\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19107\
        );

    \I__2878\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19107\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__19138\,
            I => \POWERLED.count_0_sqmuxa\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__19131\,
            I => \POWERLED.count_0_sqmuxa\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__19128\,
            I => \POWERLED.count_0_sqmuxa\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__19123\,
            I => \POWERLED.count_0_sqmuxa\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__19114\,
            I => \POWERLED.count_0_sqmuxa\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__19107\,
            I => \POWERLED.count_0_sqmuxa\
        );

    \I__2871\ : InMux
    port map (
            O => \N__19094\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__19091\,
            I => \N__19088\
        );

    \I__2869\ : InMux
    port map (
            O => \N__19088\,
            I => \N__19084\
        );

    \I__2868\ : InMux
    port map (
            O => \N__19087\,
            I => \N__19081\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__19081\,
            I => \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__19078\,
            I => \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__19073\,
            I => \N__19070\
        );

    \I__2863\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19067\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__19067\,
            I => \POWERLED.un1_count_axb_12\
        );

    \I__2861\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19054\
        );

    \I__2859\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19047\
        );

    \I__2858\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19047\
        );

    \I__2857\ : InMux
    port map (
            O => \N__19058\,
            I => \N__19047\
        );

    \I__2856\ : InMux
    port map (
            O => \N__19057\,
            I => \N__19044\
        );

    \I__2855\ : Odrv12
    port map (
            O => \N__19054\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__19047\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__19044\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__19037\,
            I => \N__19033\
        );

    \I__2851\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__2850\ : InMux
    port map (
            O => \N__19033\,
            I => \N__19027\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__19030\,
            I => \POWERLED.un1_count_axb_1\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__19027\,
            I => \POWERLED.un1_count_axb_1\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__2846\ : InMux
    port map (
            O => \N__19019\,
            I => \N__19016\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__19016\,
            I => \POWERLED.un1_count_axb_2\
        );

    \I__2844\ : InMux
    port map (
            O => \N__19013\,
            I => \N__19001\
        );

    \I__2843\ : InMux
    port map (
            O => \N__19012\,
            I => \N__19001\
        );

    \I__2842\ : InMux
    port map (
            O => \N__19011\,
            I => \N__19001\
        );

    \I__2841\ : InMux
    port map (
            O => \N__19010\,
            I => \N__19001\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__19001\,
            I => \POWERLED.count_1_2\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18998\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__2838\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18991\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__18994\,
            I => \N__18987\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__18991\,
            I => \N__18984\
        );

    \I__2835\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18981\
        );

    \I__2834\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18978\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__18984\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__18981\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__18978\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18971\,
            I => \N__18965\
        );

    \I__2829\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18965\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__18965\,
            I => \POWERLED.un1_count_cry_2_c_RNICZ0Z419\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18962\,
            I => \POWERLED.un1_count_cry_2\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__2825\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18953\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__18953\,
            I => \POWERLED.un1_count_axb_4\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__18950\,
            I => \N__18947\
        );

    \I__2822\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18935\
        );

    \I__2821\ : InMux
    port map (
            O => \N__18946\,
            I => \N__18935\
        );

    \I__2820\ : InMux
    port map (
            O => \N__18945\,
            I => \N__18935\
        );

    \I__2819\ : InMux
    port map (
            O => \N__18944\,
            I => \N__18935\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__18935\,
            I => \POWERLED.count_1_4\
        );

    \I__2817\ : InMux
    port map (
            O => \N__18932\,
            I => \POWERLED.un1_count_cry_3\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \N__18926\
        );

    \I__2815\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18923\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__18923\,
            I => \N__18920\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__18920\,
            I => \POWERLED.un1_count_axb_5\
        );

    \I__2812\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18912\
        );

    \I__2811\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18907\
        );

    \I__2810\ : InMux
    port map (
            O => \N__18915\,
            I => \N__18907\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18904\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__18907\,
            I => \N__18901\
        );

    \I__2807\ : Odrv12
    port map (
            O => \N__18904\,
            I => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__18901\,
            I => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\
        );

    \I__2805\ : InMux
    port map (
            O => \N__18896\,
            I => \POWERLED.un1_count_cry_4\
        );

    \I__2804\ : InMux
    port map (
            O => \N__18893\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__2803\ : InMux
    port map (
            O => \N__18890\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__2802\ : InMux
    port map (
            O => \N__18887\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__2800\ : InMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__18878\,
            I => \N__18875\
        );

    \I__2798\ : Odrv12
    port map (
            O => \N__18875\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__2797\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__18866\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18863\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__2793\ : InMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__18857\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18851\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__18851\,
            I => \N__18848\
        );

    \I__2789\ : Odrv4
    port map (
            O => \N__18848\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__2788\ : InMux
    port map (
            O => \N__18845\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__18842\,
            I => \N__18839\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18836\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__18836\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__2783\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18827\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__18827\,
            I => \N__18824\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__18824\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__2780\ : InMux
    port map (
            O => \N__18821\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__2779\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__18815\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__2776\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__18806\,
            I => \N__18803\
        );

    \I__2774\ : Odrv12
    port map (
            O => \N__18803\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__2773\ : InMux
    port map (
            O => \N__18800\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__2771\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__18791\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__2769\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__18785\,
            I => \N__18782\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__18782\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__2766\ : InMux
    port map (
            O => \N__18779\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18773\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__18773\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__2763\ : InMux
    port map (
            O => \N__18770\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__18767\,
            I => \N__18763\
        );

    \I__2761\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18755\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18755\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18755\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__18755\,
            I => \N__18750\
        );

    \I__2757\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18747\
        );

    \I__2756\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18744\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__18750\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__18747\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__18744\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__18737\,
            I => \N__18733\
        );

    \I__2751\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18727\
        );

    \I__2750\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18720\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18720\
        );

    \I__2748\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18720\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18717\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__18727\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18720\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__18717\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__18710\,
            I => \N__18706\
        );

    \I__2742\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18698\
        );

    \I__2741\ : InMux
    port map (
            O => \N__18706\,
            I => \N__18698\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18705\,
            I => \N__18698\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__18698\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__2738\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18690\
        );

    \I__2737\ : InMux
    port map (
            O => \N__18694\,
            I => \N__18687\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__18693\,
            I => \N__18684\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__18690\,
            I => \N__18679\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__18687\,
            I => \N__18676\
        );

    \I__2733\ : InMux
    port map (
            O => \N__18684\,
            I => \N__18671\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18683\,
            I => \N__18671\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18668\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__18679\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2729\ : Odrv12
    port map (
            O => \N__18676\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__18671\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__18668\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2726\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18656\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__18656\,
            I => \POWERLED.mult1_un124_sum_i_8\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__2723\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18647\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__18644\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18641\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__2719\ : InMux
    port map (
            O => \N__18638\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__2718\ : InMux
    port map (
            O => \N__18635\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__2717\ : InMux
    port map (
            O => \N__18632\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__2716\ : InMux
    port map (
            O => \N__18629\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__2715\ : InMux
    port map (
            O => \N__18626\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__18623\,
            I => \N__18619\
        );

    \I__2713\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18611\
        );

    \I__2712\ : InMux
    port map (
            O => \N__18619\,
            I => \N__18611\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18611\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__18611\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__18608\,
            I => \N__18604\
        );

    \I__2708\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18596\
        );

    \I__2707\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18596\
        );

    \I__2706\ : InMux
    port map (
            O => \N__18603\,
            I => \N__18596\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__18596\,
            I => \N__18592\
        );

    \I__2704\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18589\
        );

    \I__2703\ : Span4Mux_v
    port map (
            O => \N__18592\,
            I => \N__18584\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__18589\,
            I => \N__18584\
        );

    \I__2701\ : Sp12to4
    port map (
            O => \N__18584\,
            I => \N__18580\
        );

    \I__2700\ : InMux
    port map (
            O => \N__18583\,
            I => \N__18577\
        );

    \I__2699\ : Odrv12
    port map (
            O => \N__18580\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__18577\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__18572\,
            I => \N__18568\
        );

    \I__2696\ : InMux
    port map (
            O => \N__18571\,
            I => \N__18560\
        );

    \I__2695\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18560\
        );

    \I__2694\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18560\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__18560\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__2692\ : IoInMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__2690\ : Span4Mux_s1_h
    port map (
            O => \N__18551\,
            I => \N__18548\
        );

    \I__2689\ : Span4Mux_h
    port map (
            O => \N__18548\,
            I => \N__18545\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__18545\,
            I => vccst_en
        );

    \I__2687\ : IoInMux
    port map (
            O => \N__18542\,
            I => \N__18539\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__18539\,
            I => \N__18536\
        );

    \I__2685\ : Odrv12
    port map (
            O => \N__18536\,
            I => \G_12\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__2683\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__18527\,
            I => \POWERLED.mult1_un68_sum_i_8\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__18524\,
            I => \N__18521\
        );

    \I__2680\ : InMux
    port map (
            O => \N__18521\,
            I => \N__18518\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__18518\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__2677\ : InMux
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__18509\,
            I => \N__18506\
        );

    \I__2675\ : Span4Mux_h
    port map (
            O => \N__18506\,
            I => \N__18503\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__18503\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__2672\ : InMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__2670\ : Odrv4
    port map (
            O => \N__18491\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18484\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18481\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__18484\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__18481\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__2665\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18472\
        );

    \I__2664\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18469\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__18472\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__18469\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__18464\,
            I => \N__18460\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18457\
        );

    \I__2659\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18454\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__18457\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__18454\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__2656\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18445\
        );

    \I__2655\ : InMux
    port map (
            O => \N__18448\,
            I => \N__18442\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18445\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__18442\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__2652\ : InMux
    port map (
            O => \N__18437\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__18431\,
            I => \N__18428\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__18428\,
            I => \N__18425\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__18425\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18422\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__2646\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18416\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__18416\,
            I => \N__18413\
        );

    \I__2644\ : Span4Mux_v
    port map (
            O => \N__18413\,
            I => \N__18410\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__18410\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__2642\ : InMux
    port map (
            O => \N__18407\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__2641\ : CascadeMux
    port map (
            O => \N__18404\,
            I => \N__18401\
        );

    \I__2640\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__18398\,
            I => \N__18395\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__2637\ : Odrv4
    port map (
            O => \N__18392\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__2636\ : InMux
    port map (
            O => \N__18389\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__18386\,
            I => \N__18383\
        );

    \I__2634\ : InMux
    port map (
            O => \N__18383\,
            I => \N__18380\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__18374\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__2630\ : InMux
    port map (
            O => \N__18371\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__2629\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18362\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__18362\,
            I => \N__18359\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__18359\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18356\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__2624\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18350\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__18350\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__18347\,
            I => \N__18342\
        );

    \I__2621\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18339\
        );

    \I__2620\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18336\
        );

    \I__2619\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18333\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__18339\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__18336\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__18333\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2615\ : InMux
    port map (
            O => \N__18326\,
            I => \N__18322\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18325\,
            I => \N__18319\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__18322\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__18319\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__2611\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18310\
        );

    \I__2610\ : InMux
    port map (
            O => \N__18313\,
            I => \N__18307\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__18310\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__18307\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \N__18298\
        );

    \I__2606\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18295\
        );

    \I__2605\ : InMux
    port map (
            O => \N__18298\,
            I => \N__18292\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__18295\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__18292\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__2602\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18283\
        );

    \I__2601\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18280\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__18283\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__18280\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__2598\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18271\
        );

    \I__2597\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__18271\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__18268\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__2594\ : InMux
    port map (
            O => \N__18263\,
            I => \N__18259\
        );

    \I__2593\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18256\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__18259\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__18256\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__18251\,
            I => \N__18247\
        );

    \I__2589\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18244\
        );

    \I__2588\ : InMux
    port map (
            O => \N__18247\,
            I => \N__18241\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__18244\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__18241\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__2585\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18232\
        );

    \I__2584\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18229\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__18232\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__18229\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__2581\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18220\
        );

    \I__2580\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18217\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__18220\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__18217\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__2577\ : InMux
    port map (
            O => \N__18212\,
            I => \N__18208\
        );

    \I__2576\ : InMux
    port map (
            O => \N__18211\,
            I => \N__18205\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__18208\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__18205\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__18200\,
            I => \N__18196\
        );

    \I__2572\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18193\
        );

    \I__2571\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18190\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__18193\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__18190\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__2568\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18181\
        );

    \I__2567\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18178\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__18181\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__18178\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__18173\,
            I => \N__18169\
        );

    \I__2563\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18166\
        );

    \I__2562\ : InMux
    port map (
            O => \N__18169\,
            I => \N__18163\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__18166\,
            I => \N__18156\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__18163\,
            I => \N__18156\
        );

    \I__2559\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18151\
        );

    \I__2558\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18151\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__18156\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__18151\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__18146\,
            I => \N__18143\
        );

    \I__2554\ : InMux
    port map (
            O => \N__18143\,
            I => \N__18140\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__18140\,
            I => \N__18136\
        );

    \I__2552\ : InMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__18136\,
            I => \N__18130\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__18133\,
            I => \PCH_PWRGD.N_670\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__18130\,
            I => \PCH_PWRGD.N_670\
        );

    \I__2548\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18121\
        );

    \I__2547\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18118\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__18118\,
            I => \N__18112\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__18115\,
            I => \N__18109\
        );

    \I__2543\ : Odrv12
    port map (
            O => \N__18112\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__18109\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2541\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18100\
        );

    \I__2540\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18097\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__18100\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__18097\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18092\,
            I => \N__18088\
        );

    \I__2536\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18085\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__18088\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__18085\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__18080\,
            I => \N__18076\
        );

    \I__2532\ : InMux
    port map (
            O => \N__18079\,
            I => \N__18073\
        );

    \I__2531\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18070\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__18073\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__18070\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2528\ : InMux
    port map (
            O => \N__18065\,
            I => \N__18061\
        );

    \I__2527\ : InMux
    port map (
            O => \N__18064\,
            I => \N__18058\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__18061\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__18058\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__18053\,
            I => \VPP_VDDQ.count_2_1_0_cascade_\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__18050\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__2522\ : InMux
    port map (
            O => \N__18047\,
            I => \N__18044\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__18044\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__2520\ : InMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__18038\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__2518\ : InMux
    port map (
            O => \N__18035\,
            I => \N__18030\
        );

    \I__2517\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18027\
        );

    \I__2516\ : InMux
    port map (
            O => \N__18033\,
            I => \N__18024\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__18030\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__18027\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__18024\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2512\ : InMux
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__18014\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__2510\ : InMux
    port map (
            O => \N__18011\,
            I => \N__18008\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__18008\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__18005\,
            I => \N__18000\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__18004\,
            I => \N__17997\
        );

    \I__2506\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17994\
        );

    \I__2505\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17989\
        );

    \I__2504\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17989\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__17994\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__17989\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2501\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17981\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__17981\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__17978\,
            I => \N__17974\
        );

    \I__2498\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17970\
        );

    \I__2497\ : InMux
    port map (
            O => \N__17974\,
            I => \N__17965\
        );

    \I__2496\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17965\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__17970\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__17965\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2493\ : InMux
    port map (
            O => \N__17960\,
            I => \N__17956\
        );

    \I__2492\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17953\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__17956\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__17953\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__17948\,
            I => \N__17944\
        );

    \I__2488\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17940\
        );

    \I__2487\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17935\
        );

    \I__2486\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17935\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__17940\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__17935\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2483\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17925\
        );

    \I__2482\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17920\
        );

    \I__2481\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17920\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__17925\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__17920\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2478\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17912\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17908\
        );

    \I__2476\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17905\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__17908\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__17905\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__2473\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17896\
        );

    \I__2472\ : InMux
    port map (
            O => \N__17899\,
            I => \N__17893\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__17896\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__17893\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__2469\ : InMux
    port map (
            O => \N__17888\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__2468\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17881\
        );

    \I__2467\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17878\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__17881\,
            I => \N__17873\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17873\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__17873\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__2463\ : InMux
    port map (
            O => \N__17870\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__2462\ : InMux
    port map (
            O => \N__17867\,
            I => \N__17861\
        );

    \I__2461\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17861\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17858\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__17858\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__17855\,
            I => \N__17852\
        );

    \I__2457\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17848\
        );

    \I__2456\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17845\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__17848\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__17845\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__2453\ : InMux
    port map (
            O => \N__17840\,
            I => \N__17837\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__17837\,
            I => \VPP_VDDQ.count_2_1_13\
        );

    \I__2451\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17830\
        );

    \I__2450\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17827\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__17830\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__17827\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__2447\ : CascadeMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__2446\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__17816\,
            I => \VPP_VDDQ.un9_clk_100khz_10\
        );

    \I__2444\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17809\
        );

    \I__2443\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17806\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__17809\,
            I => \N__17801\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__17806\,
            I => \N__17801\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__17801\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__2439\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__17795\,
            I => \VPP_VDDQ.un9_clk_100khz_7\
        );

    \I__2437\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__17789\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__17786\,
            I => \VPP_VDDQ.count_2_1_7_cascade_\
        );

    \I__2434\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17780\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__17780\,
            I => \N__17777\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__17777\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__2431\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17768\
        );

    \I__2430\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17768\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__17768\,
            I => \N__17765\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__17765\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17756\
        );

    \I__2426\ : InMux
    port map (
            O => \N__17761\,
            I => \N__17756\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__17756\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__2424\ : InMux
    port map (
            O => \N__17753\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__2423\ : InMux
    port map (
            O => \N__17750\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__2422\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17743\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17740\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__17743\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__17740\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__17735\,
            I => \N__17731\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__17734\,
            I => \N__17728\
        );

    \I__2416\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17723\
        );

    \I__2415\ : InMux
    port map (
            O => \N__17728\,
            I => \N__17723\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__17723\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\
        );

    \I__2413\ : InMux
    port map (
            O => \N__17720\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__2412\ : InMux
    port map (
            O => \N__17717\,
            I => \N__17711\
        );

    \I__2411\ : InMux
    port map (
            O => \N__17716\,
            I => \N__17711\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17711\,
            I => \N__17708\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__17708\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\
        );

    \I__2408\ : InMux
    port map (
            O => \N__17705\,
            I => \bfn_5_3_0_\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__17702\,
            I => \N__17699\
        );

    \I__2406\ : InMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__17696\,
            I => \N__17692\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17689\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__17692\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__17689\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17684\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__2400\ : InMux
    port map (
            O => \N__17681\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__2399\ : InMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__17675\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__2397\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17666\
        );

    \I__2396\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17666\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__17666\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\
        );

    \I__2394\ : InMux
    port map (
            O => \N__17663\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__2393\ : InMux
    port map (
            O => \N__17660\,
            I => \N__17656\
        );

    \I__2392\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17653\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__17656\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__17653\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__2389\ : InMux
    port map (
            O => \N__17648\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__17645\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__17639\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__2385\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17633\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__17633\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17624\
        );

    \I__2382\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17624\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__17624\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\
        );

    \I__2380\ : InMux
    port map (
            O => \N__17621\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__2379\ : InMux
    port map (
            O => \N__17618\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__2378\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17609\
        );

    \I__2377\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17609\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__17609\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\
        );

    \I__2375\ : InMux
    port map (
            O => \N__17606\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__2374\ : InMux
    port map (
            O => \N__17603\,
            I => \N__17600\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__17600\,
            I => \N__17596\
        );

    \I__2372\ : InMux
    port map (
            O => \N__17599\,
            I => \N__17593\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__17596\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__17593\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__17588\,
            I => \N__17585\
        );

    \I__2368\ : InMux
    port map (
            O => \N__17585\,
            I => \N__17579\
        );

    \I__2367\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17579\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__17579\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\
        );

    \I__2365\ : InMux
    port map (
            O => \N__17576\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__2364\ : InMux
    port map (
            O => \N__17573\,
            I => \N__17570\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__17570\,
            I => \POWERLED.count_0_14\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__17567\,
            I => \POWERLED.countZ0Z_14_cascade_\
        );

    \I__2361\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__17561\,
            I => \N__17558\
        );

    \I__2359\ : Span4Mux_s3_h
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__17555\,
            I => \POWERLED.un79_clk_100khzlto15_5\
        );

    \I__2357\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17546\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__2354\ : Odrv4
    port map (
            O => \N__17543\,
            I => \POWERLED.g1_i_o4_4\
        );

    \I__2353\ : InMux
    port map (
            O => \N__17540\,
            I => \N__17537\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__17537\,
            I => \POWERLED.count_0_15\
        );

    \I__2351\ : InMux
    port map (
            O => \N__17534\,
            I => \N__17531\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__17531\,
            I => \VPP_VDDQ.count_2_0_2\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__17528\,
            I => \VPP_VDDQ.count_2_1_2_cascade_\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__17525\,
            I => \VPP_VDDQ.count_2Z0Z_2_cascade_\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__17522\,
            I => \POWERLED.count_1_0_cascade_\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__17519\,
            I => \POWERLED.countZ0Z_0_cascade_\
        );

    \I__2345\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17513\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__17513\,
            I => \POWERLED.count_1_1\
        );

    \I__2343\ : CascadeMux
    port map (
            O => \N__17510\,
            I => \POWERLED.count_1_1_cascade_\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__17507\,
            I => \POWERLED.un1_count_axb_1_cascade_\
        );

    \I__2341\ : InMux
    port map (
            O => \N__17504\,
            I => \N__17498\
        );

    \I__2340\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17498\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__17498\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2338\ : InMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__17492\,
            I => \POWERLED.count_0_0\
        );

    \I__2336\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17486\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__17486\,
            I => \POWERLED.count_0_11\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__17483\,
            I => \N__17479\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17482\,
            I => \N__17475\
        );

    \I__2332\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17470\
        );

    \I__2331\ : InMux
    port map (
            O => \N__17478\,
            I => \N__17470\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__17475\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__17470\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__17465\,
            I => \POWERLED.un79_clk_100khzlto4_0_cascade_\
        );

    \I__2327\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17458\
        );

    \I__2326\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17455\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__17458\,
            I => \N__17452\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__17455\,
            I => \N__17449\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__17452\,
            I => \POWERLED.un79_clk_100khzlt6\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__17449\,
            I => \POWERLED.un79_clk_100khzlt6\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__17444\,
            I => \N__17440\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17443\,
            I => \N__17437\
        );

    \I__2319\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17434\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17431\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__17434\,
            I => \N__17428\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__17431\,
            I => \POWERLED.mult1_un138_sum_i_8\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__17428\,
            I => \POWERLED.mult1_un138_sum_i_8\
        );

    \I__2314\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17414\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17414\
        );

    \I__2312\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17414\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__17414\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__2310\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__17405\,
            I => \N__17402\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__17402\,
            I => \POWERLED.count_RNIJEFE_0Z0Z_4\
        );

    \I__2306\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17396\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__17396\,
            I => \N__17392\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__17395\,
            I => \N__17389\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__17392\,
            I => \N__17386\
        );

    \I__2302\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__17386\,
            I => \POWERLED.mult1_un159_sum_i_8\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__17383\,
            I => \POWERLED.mult1_un159_sum_i_8\
        );

    \I__2299\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17375\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__17375\,
            I => \N__17372\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__17369\,
            I => \POWERLED.count_RNIUGSJ_0Z0Z_1\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__17366\,
            I => \N__17362\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17365\,
            I => \N__17351\
        );

    \I__2293\ : InMux
    port map (
            O => \N__17362\,
            I => \N__17351\
        );

    \I__2292\ : InMux
    port map (
            O => \N__17361\,
            I => \N__17351\
        );

    \I__2291\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17351\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__17351\,
            I => \N__17347\
        );

    \I__2289\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17344\
        );

    \I__2288\ : Span4Mux_h
    port map (
            O => \N__17347\,
            I => \N__17341\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__17344\,
            I => \N__17338\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__17341\,
            I => \POWERLED.N_660\
        );

    \I__2285\ : Odrv12
    port map (
            O => \N__17338\,
            I => \POWERLED.N_660\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__17333\,
            I => \POWERLED.count_0_sqmuxa_cascade_\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__17330\,
            I => \N__17327\
        );

    \I__2282\ : InMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__17324\,
            I => \POWERLED.mult1_un103_sum_i_8\
        );

    \I__2280\ : InMux
    port map (
            O => \N__17321\,
            I => \N__17318\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__17318\,
            I => \N__17314\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__17317\,
            I => \N__17310\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__17314\,
            I => \N__17305\
        );

    \I__2276\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17298\
        );

    \I__2275\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17298\
        );

    \I__2274\ : InMux
    port map (
            O => \N__17309\,
            I => \N__17298\
        );

    \I__2273\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17295\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__17305\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__17298\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__17295\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__2269\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17285\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__17285\,
            I => \POWERLED.mult1_un96_sum_i_8\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__17282\,
            I => \N__17279\
        );

    \I__2266\ : InMux
    port map (
            O => \N__17279\,
            I => \N__17276\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__17276\,
            I => \N__17273\
        );

    \I__2264\ : Odrv12
    port map (
            O => \N__17273\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__17270\,
            I => \POWERLED.N_437_cascade_\
        );

    \I__2262\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__17264\,
            I => \N__17260\
        );

    \I__2260\ : InMux
    port map (
            O => \N__17263\,
            I => \N__17257\
        );

    \I__2259\ : Span4Mux_s3_h
    port map (
            O => \N__17260\,
            I => \N__17254\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__17257\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__17254\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__17249\,
            I => \N__17246\
        );

    \I__2255\ : InMux
    port map (
            O => \N__17246\,
            I => \N__17240\
        );

    \I__2254\ : InMux
    port map (
            O => \N__17245\,
            I => \N__17240\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17237\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__17237\,
            I => \N__17234\
        );

    \I__2251\ : Span4Mux_s1_h
    port map (
            O => \N__17234\,
            I => \N__17229\
        );

    \I__2250\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17224\
        );

    \I__2249\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17224\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__17229\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__17224\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__17219\,
            I => \POWERLED.curr_stateZ0Z_0_cascade_\
        );

    \I__2245\ : InMux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__17213\,
            I => \POWERLED.curr_state_1_0\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__17210\,
            I => \N__17207\
        );

    \I__2242\ : InMux
    port map (
            O => \N__17207\,
            I => \N__17204\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__17204\,
            I => \POWERLED.count_0_3\
        );

    \I__2240\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17197\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__17200\,
            I => \N__17194\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__17197\,
            I => \N__17191\
        );

    \I__2237\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17188\
        );

    \I__2236\ : Odrv12
    port map (
            O => \N__17191\,
            I => \POWERLED.mult1_un152_sum_i_8\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__17188\,
            I => \POWERLED.mult1_un152_sum_i_8\
        );

    \I__2234\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__17180\,
            I => \N__17177\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__17174\,
            I => \POWERLED.count_RNIAKSS_0Z0Z_2\
        );

    \I__2230\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17168\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__17168\,
            I => \POWERLED.N_4851_i\
        );

    \I__2228\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17162\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__17162\,
            I => \POWERLED.N_4855_i\
        );

    \I__2226\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17156\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__17156\,
            I => \POWERLED.N_4856_i\
        );

    \I__2224\ : InMux
    port map (
            O => \N__17153\,
            I => \bfn_4_11_0_\
        );

    \I__2223\ : CascadeMux
    port map (
            O => \N__17150\,
            I => \N__17147\
        );

    \I__2222\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17144\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__17141\,
            I => \POWERLED.mult1_un117_sum_i_8\
        );

    \I__2219\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17134\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__17137\,
            I => \N__17130\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__17134\,
            I => \N__17125\
        );

    \I__2216\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17118\
        );

    \I__2215\ : InMux
    port map (
            O => \N__17130\,
            I => \N__17118\
        );

    \I__2214\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17118\
        );

    \I__2213\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17115\
        );

    \I__2212\ : Odrv12
    port map (
            O => \N__17125\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__17118\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__17115\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__2208\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17102\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__17102\,
            I => \POWERLED.mult1_un110_sum_i_8\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__17099\,
            I => \N__17096\
        );

    \I__2205\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17093\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__17093\,
            I => \POWERLED.mult1_un89_sum_i_8\
        );

    \I__2203\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17087\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__17087\,
            I => \N__17083\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__17086\,
            I => \N__17080\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__17083\,
            I => \N__17074\
        );

    \I__2199\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17067\
        );

    \I__2198\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17067\
        );

    \I__2197\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17067\
        );

    \I__2196\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17064\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__17074\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__17067\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__17064\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__2192\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__17054\,
            I => \N__17050\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__17053\,
            I => \N__17047\
        );

    \I__2189\ : Span4Mux_h
    port map (
            O => \N__17050\,
            I => \N__17041\
        );

    \I__2188\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17034\
        );

    \I__2187\ : InMux
    port map (
            O => \N__17046\,
            I => \N__17034\
        );

    \I__2186\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17034\
        );

    \I__2185\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17031\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__17041\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__17034\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__17031\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2181\ : InMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__17018\,
            I => \N__17015\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__17015\,
            I => \POWERLED.count_RNIGTVS_1Z0Z_5\
        );

    \I__2177\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__17009\,
            I => \N__17005\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__17008\,
            I => \N__17002\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__17005\,
            I => \N__16999\
        );

    \I__2173\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__16999\,
            I => \POWERLED.mult1_un131_sum_i_8\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__16996\,
            I => \POWERLED.mult1_un131_sum_i_8\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__16991\,
            I => \N__16988\
        );

    \I__2169\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__16985\,
            I => \POWERLED.count_i_6\
        );

    \I__2167\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__16979\,
            I => \POWERLED.N_4841_i\
        );

    \I__2165\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16973\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__16973\,
            I => \POWERLED.count_i_8\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16967\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__16967\,
            I => \POWERLED.N_4849_i\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__2160\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16958\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__16958\,
            I => \POWERLED.count_i_10\
        );

    \I__2158\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16952\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__16952\,
            I => \POWERLED.count_i_11\
        );

    \I__2156\ : InMux
    port map (
            O => \N__16949\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__2155\ : InMux
    port map (
            O => \N__16946\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__2154\ : InMux
    port map (
            O => \N__16943\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__2153\ : InMux
    port map (
            O => \N__16940\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__16937\,
            I => \N__16934\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16928\
        );

    \I__2150\ : InMux
    port map (
            O => \N__16933\,
            I => \N__16928\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__16928\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2148\ : InMux
    port map (
            O => \N__16925\,
            I => \N__16919\
        );

    \I__2147\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16919\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__16919\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__16916\,
            I => \N__16912\
        );

    \I__2144\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16907\
        );

    \I__2143\ : InMux
    port map (
            O => \N__16912\,
            I => \N__16907\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__16907\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16904\,
            I => \N__16898\
        );

    \I__2140\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16898\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__16898\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2138\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16892\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__16892\,
            I => \POWERLED.N_4842_i\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__16889\,
            I => \N__16886\
        );

    \I__2135\ : InMux
    port map (
            O => \N__16886\,
            I => \N__16883\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__16883\,
            I => \POWERLED.count_i_3\
        );

    \I__2133\ : InMux
    port map (
            O => \N__16880\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__2132\ : InMux
    port map (
            O => \N__16877\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__2131\ : InMux
    port map (
            O => \N__16874\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__2130\ : InMux
    port map (
            O => \N__16871\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__2129\ : InMux
    port map (
            O => \N__16868\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__2128\ : InMux
    port map (
            O => \N__16865\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__2127\ : InMux
    port map (
            O => \N__16862\,
            I => \bfn_4_8_0_\
        );

    \I__2126\ : InMux
    port map (
            O => \N__16859\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__2125\ : InMux
    port map (
            O => \N__16856\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__2124\ : InMux
    port map (
            O => \N__16853\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__2123\ : InMux
    port map (
            O => \N__16850\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__2122\ : InMux
    port map (
            O => \N__16847\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__2121\ : InMux
    port map (
            O => \N__16844\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__2120\ : InMux
    port map (
            O => \N__16841\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__2119\ : InMux
    port map (
            O => \N__16838\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__2118\ : InMux
    port map (
            O => \N__16835\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__2117\ : InMux
    port map (
            O => \N__16832\,
            I => \bfn_4_7_0_\
        );

    \I__2116\ : InMux
    port map (
            O => \N__16829\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__16826\,
            I => \VPP_VDDQ.count_2_1_10_cascade_\
        );

    \I__2114\ : InMux
    port map (
            O => \N__16823\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__2113\ : InMux
    port map (
            O => \N__16820\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__2112\ : InMux
    port map (
            O => \N__16817\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__2111\ : InMux
    port map (
            O => \N__16814\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__2110\ : InMux
    port map (
            O => \N__16811\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__2109\ : InMux
    port map (
            O => \N__16808\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__2108\ : InMux
    port map (
            O => \N__16805\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__2107\ : InMux
    port map (
            O => \N__16802\,
            I => \bfn_4_6_0_\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__16799\,
            I => \VPP_VDDQ.count_2Z0Z_12_cascade_\
        );

    \I__2105\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16793\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__16793\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__2103\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16787\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__16787\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__2101\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16781\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__16781\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__2099\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16775\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__16775\,
            I => \N__16772\
        );

    \I__2097\ : Span12Mux_s10_h
    port map (
            O => \N__16772\,
            I => \N__16765\
        );

    \I__2096\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16756\
        );

    \I__2095\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16756\
        );

    \I__2094\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16756\
        );

    \I__2093\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16756\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__16765\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__16756\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__2090\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16745\
        );

    \I__2089\ : InMux
    port map (
            O => \N__16750\,
            I => \N__16745\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__16745\,
            I => \N__16742\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__16742\,
            I => \N__16738\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__16741\,
            I => \N__16735\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__16738\,
            I => \N__16728\
        );

    \I__2084\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16717\
        );

    \I__2083\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16717\
        );

    \I__2082\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16717\
        );

    \I__2081\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16717\
        );

    \I__2080\ : InMux
    port map (
            O => \N__16731\,
            I => \N__16717\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__16728\,
            I => \VPP_VDDQ_curr_state_1\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__16717\,
            I => \VPP_VDDQ_curr_state_1\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__16712\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\
        );

    \I__2076\ : InMux
    port map (
            O => \N__16709\,
            I => \N__16706\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__16706\,
            I => \N__16703\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__16703\,
            I => \N__16699\
        );

    \I__2073\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16694\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__16699\,
            I => \N__16691\
        );

    \I__2071\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16686\
        );

    \I__2070\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16686\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__16694\,
            I => \N_626\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__16691\,
            I => \N_626\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__16686\,
            I => \N_626\
        );

    \I__2066\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16673\
        );

    \I__2065\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16670\
        );

    \I__2064\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16667\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16664\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16661\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__16670\,
            I => \N__16658\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__16667\,
            I => \N__16655\
        );

    \I__2059\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16652\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__16661\,
            I => \N__16649\
        );

    \I__2057\ : Span12Mux_s1_h
    port map (
            O => \N__16658\,
            I => \N__16646\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__16655\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__16652\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__16649\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__16646\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16633\
        );

    \I__2051\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16630\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16627\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16630\,
            I => \N__16624\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__16627\,
            I => \N__16621\
        );

    \I__2047\ : Span12Mux_s1_v
    port map (
            O => \N__16624\,
            I => \N__16618\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__16621\,
            I => \PCH_PWRGD.N_38_f0\
        );

    \I__2045\ : Odrv12
    port map (
            O => \N__16618\,
            I => \PCH_PWRGD.N_38_f0\
        );

    \I__2044\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16610\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__16610\,
            I => \N__16606\
        );

    \I__2042\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16603\
        );

    \I__2041\ : Span4Mux_s3_v
    port map (
            O => \N__16606\,
            I => \N__16600\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__16603\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__16600\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__16589\,
            I => \VPP_VDDQ.count_2_0_10\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__16586\,
            I => \VPP_VDDQ.count_2_1_14_cascade_\
        );

    \I__2034\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \VPP_VDDQ.count_2_1_4_cascade_\
        );

    \I__2033\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16577\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__16577\,
            I => \VPP_VDDQ.count_2_0_4\
        );

    \I__2031\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16571\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__16571\,
            I => \VPP_VDDQ.count_2_0_5\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__16568\,
            I => \VPP_VDDQ.count_2_1_5_cascade_\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__16565\,
            I => \VPP_VDDQ.count_2_1_12_cascade_\
        );

    \I__2027\ : InMux
    port map (
            O => \N__16562\,
            I => \bfn_2_16_0_\
        );

    \I__2026\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16555\
        );

    \I__2025\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16552\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__16555\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__16552\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__2022\ : CEMux
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__16544\,
            I => \N__16541\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__2019\ : Span4Mux_s1_h
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__16535\,
            I => \VPP_VDDQ.N_92_0\
        );

    \I__2017\ : SRMux
    port map (
            O => \N__16532\,
            I => \N__16527\
        );

    \I__2016\ : SRMux
    port map (
            O => \N__16531\,
            I => \N__16524\
        );

    \I__2015\ : SRMux
    port map (
            O => \N__16530\,
            I => \N__16521\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__16527\,
            I => \N__16518\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__16524\,
            I => \N__16513\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__16521\,
            I => \N__16513\
        );

    \I__2011\ : Span4Mux_v
    port map (
            O => \N__16518\,
            I => \N__16508\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__16513\,
            I => \N__16508\
        );

    \I__2009\ : Span4Mux_s1_h
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__16505\,
            I => \G_30\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__16502\,
            I => \VPP_VDDQ.count_2_1_8_cascade_\
        );

    \I__2006\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__16496\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__16493\,
            I => \VPP_VDDQ.count_2_1_9_cascade_\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16487\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__16487\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16484\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__2000\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16477\
        );

    \I__1999\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16474\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__16477\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__16474\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__1996\ : InMux
    port map (
            O => \N__16469\,
            I => \bfn_2_15_0_\
        );

    \I__1995\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16462\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16459\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__16462\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__16459\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__1991\ : InMux
    port map (
            O => \N__16454\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__1990\ : InMux
    port map (
            O => \N__16451\,
            I => \N__16447\
        );

    \I__1989\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16444\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__16447\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__16444\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__1986\ : InMux
    port map (
            O => \N__16439\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__16436\,
            I => \N__16432\
        );

    \I__1984\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16429\
        );

    \I__1983\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16426\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__16429\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__16426\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__1980\ : InMux
    port map (
            O => \N__16421\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__16418\,
            I => \N__16414\
        );

    \I__1978\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16411\
        );

    \I__1977\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16408\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__16411\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__16408\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__1974\ : InMux
    port map (
            O => \N__16403\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16396\
        );

    \I__1972\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16393\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__16396\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__16393\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16388\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__1968\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16381\
        );

    \I__1967\ : InMux
    port map (
            O => \N__16384\,
            I => \N__16378\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__16381\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__16378\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16373\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \POWERLED.un79_clk_100khz_cascade_\
        );

    \I__1962\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16352\
        );

    \I__1961\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16352\
        );

    \I__1960\ : InMux
    port map (
            O => \N__16365\,
            I => \N__16352\
        );

    \I__1959\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16352\
        );

    \I__1958\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16349\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16344\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16344\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__16352\,
            I => \POWERLED.N_2360_i\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__16349\,
            I => \POWERLED.N_2360_i\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__16344\,
            I => \POWERLED.N_2360_i\
        );

    \I__1952\ : SRMux
    port map (
            O => \N__16337\,
            I => \N__16334\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__1950\ : Span4Mux_s1_h
    port map (
            O => \N__16331\,
            I => \N__16328\
        );

    \I__1949\ : Odrv4
    port map (
            O => \N__16328\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__16325\,
            I => \N__16321\
        );

    \I__1947\ : InMux
    port map (
            O => \N__16324\,
            I => \N__16318\
        );

    \I__1946\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16315\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__16318\,
            I => \N__16310\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__16315\,
            I => \N__16310\
        );

    \I__1943\ : Odrv12
    port map (
            O => \N__16310\,
            I => \VPP_VDDQ.N_64_i\
        );

    \I__1942\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16303\
        );

    \I__1941\ : InMux
    port map (
            O => \N__16306\,
            I => \N__16300\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__16303\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__16300\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__16295\,
            I => \N__16291\
        );

    \I__1937\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16288\
        );

    \I__1936\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16285\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__16288\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__16285\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__1933\ : InMux
    port map (
            O => \N__16280\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__1932\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16273\
        );

    \I__1931\ : InMux
    port map (
            O => \N__16276\,
            I => \N__16270\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__16273\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__16270\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__1928\ : InMux
    port map (
            O => \N__16265\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__1927\ : InMux
    port map (
            O => \N__16262\,
            I => \N__16258\
        );

    \I__1926\ : InMux
    port map (
            O => \N__16261\,
            I => \N__16255\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__16258\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__16255\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__1923\ : InMux
    port map (
            O => \N__16250\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__1922\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16243\
        );

    \I__1921\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16240\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__16243\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__16240\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__1918\ : InMux
    port map (
            O => \N__16235\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__1917\ : InMux
    port map (
            O => \N__16232\,
            I => \N__16228\
        );

    \I__1916\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16225\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__16228\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__16225\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__1913\ : InMux
    port map (
            O => \N__16220\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__1912\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16213\
        );

    \I__1911\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16210\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__16213\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__16210\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__1908\ : InMux
    port map (
            O => \N__16205\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__16202\,
            I => \N__16198\
        );

    \I__1906\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16195\
        );

    \I__1905\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16192\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__16195\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__16192\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__1902\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__16184\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__1900\ : InMux
    port map (
            O => \N__16181\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__1899\ : InMux
    port map (
            O => \N__16178\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__1897\ : InMux
    port map (
            O => \N__16172\,
            I => \N__16163\
        );

    \I__1896\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16163\
        );

    \I__1895\ : InMux
    port map (
            O => \N__16170\,
            I => \N__16163\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__16163\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__16160\,
            I => \POWERLED.count_1_5_cascade_\
        );

    \I__1892\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16150\
        );

    \I__1891\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16150\
        );

    \I__1890\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16147\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__16150\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__16147\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__16142\,
            I => \N__16139\
        );

    \I__1886\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16133\
        );

    \I__1885\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16133\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__16133\,
            I => \POWERLED.count_1_5\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__16130\,
            I => \POWERLED.un79_clk_100khzlto6_0_cascade_\
        );

    \I__1882\ : InMux
    port map (
            O => \N__16127\,
            I => \N__16123\
        );

    \I__1881\ : InMux
    port map (
            O => \N__16126\,
            I => \N__16120\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__16123\,
            I => \POWERLED.un79_clk_100khz\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__16120\,
            I => \POWERLED.un79_clk_100khz\
        );

    \I__1878\ : InMux
    port map (
            O => \N__16115\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__16112\,
            I => \N__16109\
        );

    \I__1876\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16106\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__16106\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__1874\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16100\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__16100\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__1872\ : InMux
    port map (
            O => \N__16097\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__1871\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16091\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__16091\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__1869\ : InMux
    port map (
            O => \N__16088\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__16085\,
            I => \N__16081\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16073\
        );

    \I__1866\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16073\
        );

    \I__1865\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16073\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__16073\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1863\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16067\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__16067\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__1861\ : InMux
    port map (
            O => \N__16064\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__16061\,
            I => \N__16058\
        );

    \I__1859\ : InMux
    port map (
            O => \N__16058\,
            I => \N__16055\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__16055\,
            I => \N__16052\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__16052\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__1856\ : InMux
    port map (
            O => \N__16049\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__1855\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__16043\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__1853\ : InMux
    port map (
            O => \N__16040\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__16037\,
            I => \N__16034\
        );

    \I__1851\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__16031\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__1849\ : InMux
    port map (
            O => \N__16028\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__16025\,
            I => \N__16022\
        );

    \I__1847\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16019\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__16019\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__1845\ : InMux
    port map (
            O => \N__16016\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__1844\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__16010\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__1842\ : InMux
    port map (
            O => \N__16007\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__1841\ : InMux
    port map (
            O => \N__16004\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__1839\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15995\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__15995\,
            I => \POWERLED.mult1_un124_sum_axb_4_l_fx\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15986\
        );

    \I__1836\ : InMux
    port map (
            O => \N__15991\,
            I => \N__15986\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__15986\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__1834\ : InMux
    port map (
            O => \N__15983\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__1833\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15977\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__15977\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__15974\,
            I => \N__15971\
        );

    \I__1830\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15968\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__15968\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__1828\ : InMux
    port map (
            O => \N__15965\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__1827\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15959\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__15959\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__1825\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15953\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__15953\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__1823\ : InMux
    port map (
            O => \N__15950\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__1821\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__15941\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__15938\,
            I => \N_626_cascade_\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__15935\,
            I => \POWERLED.G_30Z0Z_0_cascade_\
        );

    \I__1817\ : InMux
    port map (
            O => \N__15932\,
            I => \N__15926\
        );

    \I__1816\ : InMux
    port map (
            O => \N__15931\,
            I => \N__15926\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__15926\,
            I => \N__15923\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__15923\,
            I => \N__15920\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__15920\,
            I => \VPP_VDDQ_un6_count\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__15917\,
            I => \G_30_cascade_\
        );

    \I__1811\ : InMux
    port map (
            O => \N__15914\,
            I => \N__15911\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__15911\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__1809\ : InMux
    port map (
            O => \N__15908\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__15905\,
            I => \N__15902\
        );

    \I__1807\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15899\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__15899\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__1805\ : InMux
    port map (
            O => \N__15896\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__1804\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15887\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__15887\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__1801\ : InMux
    port map (
            O => \N__15884\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__1800\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15878\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__15878\,
            I => \N__15875\
        );

    \I__1798\ : Odrv12
    port map (
            O => \N__15875\,
            I => \PCH_PWRGD.curr_state_0_0\
        );

    \I__1797\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15869\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__15869\,
            I => \PCH_PWRGD.N_2244_i\
        );

    \I__1795\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15860\
        );

    \I__1794\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15860\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__15860\,
            I => \N__15857\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__15857\,
            I => \N__15854\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__15854\,
            I => vr_ready_vccin
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__15851\,
            I => \PCH_PWRGD.N_2244_i_cascade_\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__15848\,
            I => \PCH_PWRGD.N_655_cascade_\
        );

    \I__1788\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15842\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__15842\,
            I => \PCH_PWRGD.m6_i_i_a2\
        );

    \I__1786\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15835\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__15838\,
            I => \N__15832\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__15835\,
            I => \N__15827\
        );

    \I__1783\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15824\
        );

    \I__1782\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15819\
        );

    \I__1781\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15819\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__15827\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__15824\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__15819\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1777\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15806\
        );

    \I__1776\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15806\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__15806\,
            I => \N__15789\
        );

    \I__1774\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15784\
        );

    \I__1773\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15784\
        );

    \I__1772\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15781\
        );

    \I__1771\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15777\
        );

    \I__1770\ : InMux
    port map (
            O => \N__15801\,
            I => \N__15770\
        );

    \I__1769\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15770\
        );

    \I__1768\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15770\
        );

    \I__1767\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15763\
        );

    \I__1766\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15763\
        );

    \I__1765\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15763\
        );

    \I__1764\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15754\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15754\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15754\
        );

    \I__1761\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15754\
        );

    \I__1760\ : Span4Mux_s1_h
    port map (
            O => \N__15789\,
            I => \N__15747\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__15784\,
            I => \N__15747\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__15781\,
            I => \N__15747\
        );

    \I__1757\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15744\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__15777\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__15770\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__15763\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__15754\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__15747\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__15744\,
            I => \PCH_PWRGD.N_386\
        );

    \I__1750\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15724\
        );

    \I__1749\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15721\
        );

    \I__1748\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15718\
        );

    \I__1747\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15715\
        );

    \I__1746\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15712\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__15724\,
            I => \N__15707\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__15721\,
            I => \N__15707\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__15718\,
            I => \N__15702\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__15715\,
            I => \N__15702\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__15712\,
            I => \N__15699\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__15707\,
            I => \N__15696\
        );

    \I__1739\ : Odrv12
    port map (
            O => \N__15702\,
            I => \PCH_PWRGD.N_2226_i\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__15699\,
            I => \PCH_PWRGD.N_2226_i\
        );

    \I__1737\ : Odrv4
    port map (
            O => \N__15696\,
            I => \PCH_PWRGD.N_2226_i\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__15689\,
            I => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__1735\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15681\
        );

    \I__1734\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15678\
        );

    \I__1733\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15675\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15681\,
            I => \PCH_PWRGD.N_655\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__15678\,
            I => \PCH_PWRGD.N_655\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__15675\,
            I => \PCH_PWRGD.N_655\
        );

    \I__1729\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__15665\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__1727\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__15659\,
            I => \PCH_PWRGD.count_rst_14\
        );

    \I__1725\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15653\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__15653\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__15650\,
            I => \PCH_PWRGD.count_0_sqmuxa_cascade_\
        );

    \I__1722\ : InMux
    port map (
            O => \N__15647\,
            I => \N__15644\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__15644\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__15641\,
            I => \PCH_PWRGD.countZ0Z_6_cascade_\
        );

    \I__1719\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15635\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__15635\,
            I => \PCH_PWRGD.count_1_i_a2_0_0\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__15632\,
            I => \PCH_PWRGD.un2_count_1_axb_1_cascade_\
        );

    \I__1716\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15626\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__15626\,
            I => \N__15622\
        );

    \I__1714\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15619\
        );

    \I__1713\ : Odrv12
    port map (
            O => \N__15622\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__15619\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__1711\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15608\
        );

    \I__1710\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15608\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15608\,
            I => \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\
        );

    \I__1708\ : InMux
    port map (
            O => \N__15605\,
            I => \N__15602\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__15602\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15599\,
            I => \N__15596\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__15596\,
            I => \PCH_PWRGD.un2_count_1_axb_10\
        );

    \I__1704\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15584\
        );

    \I__1703\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15584\
        );

    \I__1702\ : InMux
    port map (
            O => \N__15591\,
            I => \N__15584\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__15584\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15575\
        );

    \I__1699\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15575\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__15575\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__1697\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15566\
        );

    \I__1696\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15566\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__15563\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__15560\,
            I => \PCH_PWRGD.countZ0Z_3_cascade_\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__15554\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__1690\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__15548\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__15545\,
            I => \PCH_PWRGD.countZ0Z_14_cascade_\
        );

    \I__1687\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15538\
        );

    \I__1686\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15535\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__15538\,
            I => \N__15532\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__15535\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__15532\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__15527\,
            I => \PCH_PWRGD.count_1_i_a2_1_0_cascade_\
        );

    \I__1681\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__15518\,
            I => \PCH_PWRGD.count_1_i_a2_2_0\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \N__15512\
        );

    \I__1677\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15506\
        );

    \I__1676\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15506\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__15506\,
            I => \PCH_PWRGD.count_1_i_a2_11_0\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__15503\,
            I => \PCH_PWRGD.count_1_i_a2_11_0_cascade_\
        );

    \I__1673\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15497\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__15497\,
            I => \N__15492\
        );

    \I__1671\ : InMux
    port map (
            O => \N__15496\,
            I => \N__15487\
        );

    \I__1670\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15487\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__15492\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__15487\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__1667\ : InMux
    port map (
            O => \N__15482\,
            I => \N__15476\
        );

    \I__1666\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15476\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__15476\,
            I => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__15473\,
            I => \N__15470\
        );

    \I__1663\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__15467\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__1661\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15455\
        );

    \I__1660\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15455\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15462\,
            I => \N__15455\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__15455\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1657\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15446\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15446\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__15446\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1654\ : InMux
    port map (
            O => \N__15443\,
            I => \N__15440\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__15440\,
            I => \PCH_PWRGD.un2_count_1_axb_2\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__15437\,
            I => \PCH_PWRGD.countZ0Z_11_cascade_\
        );

    \I__1651\ : InMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__15431\,
            I => \PCH_PWRGD.count_1_i_a2_4_0\
        );

    \I__1649\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15425\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__15425\,
            I => \PCH_PWRGD.count_1_i_a2_5_0\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \PCH_PWRGD.count_1_i_a2_3_0_cascade_\
        );

    \I__1646\ : InMux
    port map (
            O => \N__15419\,
            I => \N__15416\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__15416\,
            I => \PCH_PWRGD.count_1_i_a2_6_0\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__15413\,
            I => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__15410\,
            I => \PCH_PWRGD.N_2226_i_cascade_\
        );

    \I__1642\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15404\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__15404\,
            I => \PCH_PWRGD.curr_state_7_0\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__15401\,
            I => \PCH_PWRGD.N_386_cascade_\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__15398\,
            I => \PCH_PWRGD.count_rst_11_cascade_\
        );

    \I__1638\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15390\
        );

    \I__1637\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15387\
        );

    \I__1636\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15384\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__15390\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__15387\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__15384\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1632\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15373\
        );

    \I__1631\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15370\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__15373\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__15370\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__1628\ : InMux
    port map (
            O => \N__15365\,
            I => \HDA_STRAP.un1_count_1_cry_14\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15357\
        );

    \I__1626\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15352\
        );

    \I__1625\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15352\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__15357\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__15352\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__1622\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__15344\,
            I => \HDA_STRAP.un1_count_1_cry_15_THRU_CO\
        );

    \I__1620\ : InMux
    port map (
            O => \N__15341\,
            I => \bfn_2_3_0_\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \N__15330\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__15337\,
            I => \N__15326\
        );

    \I__1617\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15321\
        );

    \I__1616\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15321\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__15334\,
            I => \N__15316\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__15333\,
            I => \N__15313\
        );

    \I__1613\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15309\
        );

    \I__1612\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15306\
        );

    \I__1611\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15303\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__15321\,
            I => \N__15300\
        );

    \I__1609\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15289\
        );

    \I__1608\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15289\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15289\
        );

    \I__1606\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15289\
        );

    \I__1605\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15289\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__15309\,
            I => \N__15284\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__15306\,
            I => \N__15284\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15281\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__15300\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__15289\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__15284\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__15281\,
            I => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \N__15267\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__15271\,
            I => \N__15263\
        );

    \I__1595\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15253\
        );

    \I__1594\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15253\
        );

    \I__1593\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15250\
        );

    \I__1592\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15247\
        );

    \I__1591\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15236\
        );

    \I__1590\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15236\
        );

    \I__1589\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15236\
        );

    \I__1588\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15236\
        );

    \I__1587\ : InMux
    port map (
            O => \N__15258\,
            I => \N__15236\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__15253\,
            I => \N__15233\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__15250\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__15247\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__15236\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__15233\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1581\ : InMux
    port map (
            O => \N__15224\,
            I => \HDA_STRAP.un1_count_1_cry_16\
        );

    \I__1580\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15217\
        );

    \I__1579\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__15217\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__15214\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15205\
        );

    \I__1575\ : InMux
    port map (
            O => \N__15208\,
            I => \N__15202\
        );

    \I__1574\ : InMux
    port map (
            O => \N__15205\,
            I => \N__15199\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__15202\,
            I => \N__15194\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__15199\,
            I => \N__15194\
        );

    \I__1571\ : Span4Mux_s3_v
    port map (
            O => \N__15194\,
            I => \N__15191\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__15191\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1569\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15183\
        );

    \I__1568\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15180\
        );

    \I__1567\ : InMux
    port map (
            O => \N__15186\,
            I => \N__15177\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__15183\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__15180\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__15177\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__15170\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__1562\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15161\
        );

    \I__1561\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15161\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__15161\,
            I => \N__15158\
        );

    \I__1559\ : Span4Mux_h
    port map (
            O => \N__15158\,
            I => \N__15155\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__15155\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__1557\ : InMux
    port map (
            O => \N__15152\,
            I => \N__15149\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__15149\,
            I => \PCH_PWRGD.count_rst_7\
        );

    \I__1555\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15140\
        );

    \I__1554\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15140\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__15140\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__1552\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__15134\,
            I => \N__15129\
        );

    \I__1550\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15124\
        );

    \I__1549\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15124\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__15129\,
            I => \PCH_PWRGD.un2_count_1_axb_7\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__15124\,
            I => \PCH_PWRGD.un2_count_1_axb_7\
        );

    \I__1546\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15116\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__15116\,
            I => \PCH_PWRGD.count_rst_3\
        );

    \I__1544\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__15110\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__1542\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15104\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__15104\,
            I => \N__15100\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__15103\,
            I => \N__15097\
        );

    \I__1539\ : Span12Mux_v
    port map (
            O => \N__15100\,
            I => \N__15093\
        );

    \I__1538\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15090\
        );

    \I__1537\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15087\
        );

    \I__1536\ : Odrv12
    port map (
            O => \N__15093\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__15090\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__15087\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__15080\,
            I => \N__15077\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15073\
        );

    \I__1531\ : InMux
    port map (
            O => \N__15076\,
            I => \N__15070\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__15073\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__15070\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__1528\ : InMux
    port map (
            O => \N__15065\,
            I => \HDA_STRAP.un1_count_1_cry_6\
        );

    \I__1527\ : InMux
    port map (
            O => \N__15062\,
            I => \N__15057\
        );

    \I__1526\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15052\
        );

    \I__1525\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15052\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__15057\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__15052\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__1521\ : InMux
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__15041\,
            I => \HDA_STRAP.un1_count_1_cry_7_THRU_CO\
        );

    \I__1519\ : InMux
    port map (
            O => \N__15038\,
            I => \bfn_2_2_0_\
        );

    \I__1518\ : InMux
    port map (
            O => \N__15035\,
            I => \N__15031\
        );

    \I__1517\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15028\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__15031\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__15028\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__1514\ : InMux
    port map (
            O => \N__15023\,
            I => \HDA_STRAP.un1_count_1_cry_8\
        );

    \I__1513\ : InMux
    port map (
            O => \N__15020\,
            I => \N__15015\
        );

    \I__1512\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15012\
        );

    \I__1511\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15009\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__15015\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__15012\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__15009\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1507\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__14999\,
            I => \HDA_STRAP.un1_count_1_cry_9_THRU_CO\
        );

    \I__1505\ : InMux
    port map (
            O => \N__14996\,
            I => \HDA_STRAP.un1_count_1_cry_9\
        );

    \I__1504\ : InMux
    port map (
            O => \N__14993\,
            I => \N__14988\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14992\,
            I => \N__14985\
        );

    \I__1502\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14982\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__14988\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__14985\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__14982\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__1497\ : InMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__14969\,
            I => \HDA_STRAP.un1_count_1_cry_10_THRU_CO\
        );

    \I__1495\ : InMux
    port map (
            O => \N__14966\,
            I => \HDA_STRAP.un1_count_1_cry_10\
        );

    \I__1494\ : InMux
    port map (
            O => \N__14963\,
            I => \N__14959\
        );

    \I__1493\ : InMux
    port map (
            O => \N__14962\,
            I => \N__14956\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__14959\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__14956\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__1490\ : InMux
    port map (
            O => \N__14951\,
            I => \HDA_STRAP.un1_count_1_cry_11\
        );

    \I__1489\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14944\
        );

    \I__1488\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14941\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__14944\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__14941\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__1485\ : InMux
    port map (
            O => \N__14936\,
            I => \HDA_STRAP.un1_count_1_cry_12\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14933\,
            I => \N__14929\
        );

    \I__1483\ : InMux
    port map (
            O => \N__14932\,
            I => \N__14926\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__14929\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__14926\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__1480\ : InMux
    port map (
            O => \N__14921\,
            I => \HDA_STRAP.un1_count_1_cry_13\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14915\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__14915\,
            I => \N__14912\
        );

    \I__1477\ : Span4Mux_s3_v
    port map (
            O => \N__14912\,
            I => \N__14909\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__14909\,
            I => vpp_ok
        );

    \I__1475\ : IoInMux
    port map (
            O => \N__14906\,
            I => \N__14903\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__14903\,
            I => vddq_en
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \N__14897\
        );

    \I__1472\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14892\
        );

    \I__1471\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14889\
        );

    \I__1470\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14886\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__14892\,
            I => \N__14883\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__14889\,
            I => \N__14878\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__14886\,
            I => \N__14878\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__14883\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__14878\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14870\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__14870\,
            I => \N__14866\
        );

    \I__1462\ : InMux
    port map (
            O => \N__14869\,
            I => \N__14863\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__14866\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__14863\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__1459\ : InMux
    port map (
            O => \N__14858\,
            I => \HDA_STRAP.un1_count_1_cry_0\
        );

    \I__1458\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14851\
        );

    \I__1457\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14848\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__14851\,
            I => \N__14845\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__14848\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__14845\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__1453\ : InMux
    port map (
            O => \N__14840\,
            I => \HDA_STRAP.un1_count_1_cry_1\
        );

    \I__1452\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14833\
        );

    \I__1451\ : InMux
    port map (
            O => \N__14836\,
            I => \N__14830\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__14833\,
            I => \N__14827\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__14830\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__14827\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__1447\ : InMux
    port map (
            O => \N__14822\,
            I => \HDA_STRAP.un1_count_1_cry_2\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__14819\,
            I => \N__14816\
        );

    \I__1445\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14813\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__14813\,
            I => \N__14809\
        );

    \I__1443\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14806\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__14809\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__14806\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__1440\ : InMux
    port map (
            O => \N__14801\,
            I => \HDA_STRAP.un1_count_1_cry_3\
        );

    \I__1439\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14794\
        );

    \I__1438\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14791\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14788\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__14791\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__14788\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__1434\ : InMux
    port map (
            O => \N__14783\,
            I => \HDA_STRAP.un1_count_1_cry_4\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__14780\,
            I => \N__14776\
        );

    \I__1432\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14770\
        );

    \I__1431\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14770\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14775\,
            I => \N__14767\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__14770\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__14767\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__1427\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14759\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__14759\,
            I => \N__14756\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__14756\,
            I => \HDA_STRAP.un1_count_1_cry_5_THRU_CO\
        );

    \I__1424\ : InMux
    port map (
            O => \N__14753\,
            I => \HDA_STRAP.un1_count_1_cry_5\
        );

    \I__1423\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14747\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__14747\,
            I => \POWERLED.N_11\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__14738\,
            I => \POWERLED.g0_2_1\
        );

    \I__1418\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14729\
        );

    \I__1417\ : InMux
    port map (
            O => \N__14734\,
            I => \N__14729\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__14729\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__14726\,
            I => \POWERLED.N_2360_i_cascade_\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__14723\,
            I => \VPP_VDDQ.un6_count_11_cascade_\
        );

    \I__1413\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__14717\,
            I => \VPP_VDDQ.un6_count_9\
        );

    \I__1411\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14711\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__14711\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14705\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__14705\,
            I => \VPP_VDDQ.un6_count_8\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \N__14698\
        );

    \I__1406\ : InMux
    port map (
            O => \N__14701\,
            I => \N__14690\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14690\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14690\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__14690\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__1401\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__1399\ : Odrv4
    port map (
            O => \N__14678\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__1397\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__14666\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__14663\,
            I => \N__14659\
        );

    \I__1393\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14651\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14651\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14651\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__14648\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__14645\,
            I => \POWERLED.g1_i_a4_0_1_cascade_\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__14639\,
            I => \POWERLED.N_12\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__14636\,
            I => \POWERLED.N_5_cascade_\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__14633\,
            I => \POWERLED.pwm_out_en_cascade_\
        );

    \I__1383\ : IoInMux
    port map (
            O => \N__14630\,
            I => \N__14627\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__14624\,
            I => pwrbtn_led
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__14621\,
            I => \N__14617\
        );

    \I__1379\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14609\
        );

    \I__1378\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14609\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14609\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__14609\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__1375\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__14603\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14600\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__1371\ : InMux
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__14591\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__1369\ : InMux
    port map (
            O => \N__14588\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__1368\ : InMux
    port map (
            O => \N__14585\,
            I => \N__14582\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__14582\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__1366\ : InMux
    port map (
            O => \N__14579\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__14576\,
            I => \N__14573\
        );

    \I__1364\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14570\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__14570\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__1362\ : InMux
    port map (
            O => \N__14567\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__1361\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14561\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__14561\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__1359\ : InMux
    port map (
            O => \N__14558\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__1358\ : InMux
    port map (
            O => \N__14555\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__1357\ : InMux
    port map (
            O => \N__14552\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__1356\ : InMux
    port map (
            O => \N__14549\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__1354\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__14540\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__1352\ : InMux
    port map (
            O => \N__14537\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__1351\ : InMux
    port map (
            O => \N__14534\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__1350\ : InMux
    port map (
            O => \N__14531\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__1349\ : InMux
    port map (
            O => \N__14528\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__1348\ : InMux
    port map (
            O => \N__14525\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__1347\ : InMux
    port map (
            O => \N__14522\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__1346\ : InMux
    port map (
            O => \N__14519\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14516\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__14513\,
            I => \N__14509\
        );

    \I__1343\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14501\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14509\,
            I => \N__14501\
        );

    \I__1341\ : InMux
    port map (
            O => \N__14508\,
            I => \N__14501\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__14501\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__1339\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14495\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14495\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__1337\ : InMux
    port map (
            O => \N__14492\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14483\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__14483\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14480\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__1332\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14474\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__14474\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__1330\ : InMux
    port map (
            O => \N__14471\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__14468\,
            I => \N__14465\
        );

    \I__1328\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__14462\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__1326\ : InMux
    port map (
            O => \N__14459\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__1325\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__14453\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__1323\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14444\
        );

    \I__1322\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14444\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__14444\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__14441\,
            I => \PCH_PWRGD.countZ0Z_15_cascade_\
        );

    \I__1319\ : InMux
    port map (
            O => \N__14438\,
            I => \N__14433\
        );

    \I__1318\ : InMux
    port map (
            O => \N__14437\,
            I => \N__14428\
        );

    \I__1317\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14428\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__14433\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__14428\,
            I => \PCH_PWRGD.count_rst_1\
        );

    \I__1314\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14417\
        );

    \I__1313\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14417\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__14417\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__1311\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14411\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__14411\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__1309\ : InMux
    port map (
            O => \N__14408\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__1308\ : InMux
    port map (
            O => \N__14405\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__1307\ : InMux
    port map (
            O => \N__14402\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__1306\ : InMux
    port map (
            O => \N__14399\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14396\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__1304\ : InMux
    port map (
            O => \N__14393\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__1303\ : InMux
    port map (
            O => \N__14390\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14387\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__1301\ : InMux
    port map (
            O => \N__14384\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__1300\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14378\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__14378\,
            I => \PCH_PWRGD.un2_count_1_axb_13\
        );

    \I__1298\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__14372\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14363\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14363\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__14363\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__1293\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14357\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__14357\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__1291\ : InMux
    port map (
            O => \N__14354\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__1290\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14347\
        );

    \I__1289\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14344\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__14347\,
            I => \PCH_PWRGD.un2_count_1_axb_4\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__14344\,
            I => \PCH_PWRGD.un2_count_1_axb_4\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__14339\,
            I => \N__14335\
        );

    \I__1285\ : InMux
    port map (
            O => \N__14338\,
            I => \N__14330\
        );

    \I__1284\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14330\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__14330\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1282\ : InMux
    port map (
            O => \N__14327\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__1281\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14318\
        );

    \I__1280\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14318\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__14318\,
            I => \N__14315\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__14315\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1277\ : InMux
    port map (
            O => \N__14312\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__1276\ : InMux
    port map (
            O => \N__14309\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__1275\ : InMux
    port map (
            O => \N__14306\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__1274\ : InMux
    port map (
            O => \N__14303\,
            I => \N__14300\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__14300\,
            I => \N__14295\
        );

    \I__1272\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14290\
        );

    \I__1271\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14290\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__14295\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__14290\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__14285\,
            I => \N__14281\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14276\
        );

    \I__1266\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14276\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__14276\,
            I => \N__14273\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__14273\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1263\ : InMux
    port map (
            O => \N__14270\,
            I => \PCH_PWRGD.un2_count_1_cry_7\
        );

    \I__1262\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14264\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__14264\,
            I => \N__14260\
        );

    \I__1260\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14257\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__14260\,
            I => \PCH_PWRGD.un2_count_1_axb_9\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__14257\,
            I => \PCH_PWRGD.un2_count_1_axb_9\
        );

    \I__1257\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14246\
        );

    \I__1256\ : InMux
    port map (
            O => \N__14251\,
            I => \N__14246\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__14246\,
            I => \N__14243\
        );

    \I__1254\ : Odrv12
    port map (
            O => \N__14243\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1253\ : InMux
    port map (
            O => \N__14240\,
            I => \bfn_1_7_0_\
        );

    \I__1252\ : InMux
    port map (
            O => \N__14237\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__14234\,
            I => \PCH_PWRGD.count_rst_9_cascade_\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__14231\,
            I => \PCH_PWRGD.countZ0Z_5_cascade_\
        );

    \I__1249\ : InMux
    port map (
            O => \N__14228\,
            I => \N__14225\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__14225\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__14222\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__14219\,
            I => \PCH_PWRGD.un2_count_1_axb_4_cascade_\
        );

    \I__1245\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__14213\,
            I => \PCH_PWRGD.count_rst_10\
        );

    \I__1243\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14204\
        );

    \I__1242\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14204\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__14204\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__1240\ : InMux
    port map (
            O => \N__14201\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \I__1239\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14195\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__14192\,
            I => \HDA_STRAP.un4_count_10\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__14189\,
            I => \HDA_STRAP.un4_count_cascade_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__14183\,
            I => \PCH_PWRGD.count_rst_5\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__14180\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__14177\,
            I => \PCH_PWRGD.un2_count_1_axb_9_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14168\
        );

    \I__1230\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14168\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__14168\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__14165\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__14162\,
            I => \PCH_PWRGD.countZ0Z_8_cascade_\
        );

    \I__1226\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14156\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__14156\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__14153\,
            I => \HDA_STRAP.N_16_cascade_\
        );

    \I__1223\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14147\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__14147\,
            I => \HDA_STRAP.HDA_SDO_ATP_3_0\
        );

    \I__1221\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14140\
        );

    \I__1220\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14137\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__14140\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__14137\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__14132\,
            I => \HDA_STRAP.un4_count_9_cascade_\
        );

    \I__1216\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14126\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__14126\,
            I => \HDA_STRAP.un4_count_12\
        );

    \I__1214\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14120\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__14120\,
            I => \HDA_STRAP.un4_count_11\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__14117\,
            I => \HDA_STRAP.un4_count_13_cascade_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14111\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__14111\,
            I => \PCH_PWRGD.delayed_vccin_okZ0\
        );

    \I__1209\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14105\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__14102\,
            I => \N__14099\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__14099\,
            I => \N__14096\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__14096\,
            I => gpio_fpga_soc_1
        );

    \I__1204\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14090\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__14090\,
            I => \HDA_STRAP.m14_i_0\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__14087\,
            I => \N__14084\
        );

    \I__1201\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14069\
        );

    \I__1200\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14069\
        );

    \I__1199\ : InMux
    port map (
            O => \N__14082\,
            I => \N__14069\
        );

    \I__1198\ : InMux
    port map (
            O => \N__14081\,
            I => \N__14069\
        );

    \I__1197\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14069\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__14069\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__14066\,
            I => \N__14060\
        );

    \I__1194\ : InMux
    port map (
            O => \N__14065\,
            I => \N__14056\
        );

    \I__1193\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14047\
        );

    \I__1192\ : InMux
    port map (
            O => \N__14063\,
            I => \N__14047\
        );

    \I__1191\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14047\
        );

    \I__1190\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14047\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__14056\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__14047\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__14042\,
            I => \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_\
        );

    \I__1186\ : IoInMux
    port map (
            O => \N__14039\,
            I => \N__14036\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__14036\,
            I => \N__14033\
        );

    \I__1184\ : Span12Mux_s0_h
    port map (
            O => \N__14033\,
            I => \N__14030\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__14030\,
            I => hda_sdo_atp
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__14027\,
            I => \N_428_cascade_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_6_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_15_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_8_16_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_2_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_1_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_7\,
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_15\,
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_4_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_4_7_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_2_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_14_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_4_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_4_10_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \N_92_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__18542\,
            GLOBALBUFFEROUTPUT => \N_92_g\
        );

    \N_557_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33621\,
            GLOBALBUFFEROUTPUT => \N_557_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14114\,
            in2 => \_gnd_net_\,
            in3 => \N__30799\,
            lcout => \N_428\,
            ltout => \N_428_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001001"
        )
    port map (
            in0 => \N__14065\,
            in1 => \N__14083\,
            in2 => \N__14027\,
            in3 => \N__14093\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34403\,
            ce => \N__24047\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIJRUK1_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__16636\,
            in1 => \N__16678\,
            in2 => \N__21247\,
            in3 => \N__16613\,
            lcout => \PCH_PWRGD.delayed_vccin_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_0_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100001100"
        )
    port map (
            in0 => \N__14108\,
            in1 => \N__14063\,
            in2 => \N__15272\,
            in3 => \N__14082\,
            lcout => \HDA_STRAP.m14_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100011111000"
        )
    port map (
            in0 => \N__14064\,
            in1 => \N__15270\,
            in2 => \N__14087\,
            in3 => \N__25106\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34403\,
            ce => \N__24047\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_0_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14080\,
            in2 => \_gnd_net_\,
            in3 => \N__14059\,
            lcout => \HDA_STRAP.curr_state_RNIH91AZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIRV1F_2_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001011111"
        )
    port map (
            in0 => \N__14081\,
            in1 => \_gnd_net_\,
            in2 => \N__14066\,
            in3 => \N__14143\,
            lcout => \HDA_STRAP.HDA_SDO_ATP_3_0\,
            ltout => \HDA_STRAP.HDA_SDO_ATP_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14042\,
            in3 => \_gnd_net_\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34403\,
            ce => \N__24047\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIBJB61_7_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14962\,
            in1 => \N__15034\,
            in2 => \N__15080\,
            in3 => \N__14947\,
            lcout => \HDA_STRAP.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDLB61_6_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14932\,
            in1 => \N__15060\,
            in2 => \N__14780\,
            in3 => \N__15376\,
            lcout => \HDA_STRAP.un4_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__14762\,
            in1 => \N__15262\,
            in2 => \N__15334\,
            in3 => \N__14779\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34405\,
            ce => \N__24035\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__15260\,
            in1 => \N__15320\,
            in2 => \N__15047\,
            in3 => \N__15061\,
            lcout => \HDA_STRAP.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34405\,
            ce => \N__24035\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__15020\,
            in1 => \N__15002\,
            in2 => \N__15333\,
            in3 => \N__15261\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34405\,
            ce => \N__24035\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101110000"
        )
    port map (
            in0 => \N__15259\,
            in1 => \N__15319\,
            in2 => \N__14975\,
            in3 => \N__14993\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34405\,
            ce => \N__24035\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_2_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15258\,
            lcout => OPEN,
            ltout => \HDA_STRAP.N_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__14144\,
            in1 => \N__25107\,
            in2 => \N__14153\,
            in3 => \N__14150\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34405\,
            ce => \N__24035\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI2L821_2_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14798\,
            in1 => \N__14837\,
            in2 => \N__14819\,
            in3 => \N__14855\,
            lcout => \HDA_STRAP.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_0_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__14896\,
            in1 => \N__15335\,
            in2 => \N__15338\,
            in3 => \N__15266\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => \N__24039\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI4CB61_17_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__15360\,
            in1 => \N__14873\,
            in2 => \N__14900\,
            in3 => \N__15220\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIH7IR1_10_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14991\,
            in2 => \N__14132\,
            in3 => \N__15018\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB5IA5_2_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14129\,
            in1 => \N__14123\,
            in2 => \N__14117\,
            in3 => \N__14198\,
            lcout => \HDA_STRAP.un4_count\,
            ltout => \HDA_STRAP.un4_count_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__15347\,
            in1 => \N__15336\,
            in2 => \N__14189\,
            in3 => \N__15361\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34513\,
            ce => \N__24039\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOV3T1_0_9_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__14299\,
            in1 => \N__14186\,
            in2 => \N__25572\,
            in3 => \N__14174\,
            lcout => \PCH_PWRGD.count_1_i_a2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNIGD4H1_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__15796\,
            in1 => \N__14251\,
            in2 => \N__25409\,
            in3 => \N__14263\,
            lcout => \PCH_PWRGD.count_rst_5\,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOV3T1_9_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25544\,
            in1 => \_gnd_net_\,
            in2 => \N__14180\,
            in3 => \N__14173\,
            lcout => \PCH_PWRGD.un2_count_1_axb_9\,
            ltout => \PCH_PWRGD.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_9_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__25385\,
            in1 => \N__15811\,
            in2 => \N__14177\,
            in3 => \N__14252\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34727\,
            ce => \N__25566\,
            sr => \N__25405\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNIFB3H1_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__14298\,
            in1 => \N__25380\,
            in2 => \N__14285\,
            in3 => \N__15797\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI6A7E3_8_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14159\,
            in2 => \N__14165\,
            in3 => \N__25543\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => \PCH_PWRGD.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_8_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__14284\,
            in1 => \N__25384\,
            in2 => \N__14162\,
            in3 => \N__15798\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34727\,
            ce => \N__25566\,
            sr => \N__25405\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNIPMNB1_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15208\,
            in1 => \N__15812\,
            in2 => \N__15103\,
            in3 => \N__25406\,
            lcout => \PCH_PWRGD.count_rst_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIC50H1_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__15792\,
            in1 => \N__14323\,
            in2 => \N__25410\,
            in3 => \N__15186\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI014E3_5_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__25539\,
            in1 => \N__14228\,
            in2 => \N__14234\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => \PCH_PWRGD.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_5_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__15794\,
            in1 => \N__25367\,
            in2 => \N__14231\,
            in3 => \N__14324\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34700\,
            ce => \N__25573\,
            sr => \N__25391\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNIB3VG1_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__14350\,
            in1 => \N__25386\,
            in2 => \N__14339\,
            in3 => \N__15793\,
            lcout => \PCH_PWRGD.count_rst_10\,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIJQ3T1_4_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25538\,
            in2 => \N__14222\,
            in3 => \N__14210\,
            lcout => \PCH_PWRGD.un2_count_1_axb_4\,
            ltout => \PCH_PWRGD.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__14338\,
            in1 => \N__25390\,
            in2 => \N__14219\,
            in3 => \N__15795\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34700\,
            ce => \N__25573\,
            sr => \N__25391\
        );

    \PCH_PWRGD.count_RNIJQ3T1_0_4_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__14216\,
            in1 => \N__14209\,
            in2 => \N__25584\,
            in3 => \N__15393\,
            lcout => \PCH_PWRGD.count_1_i_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25621\,
            in2 => \N__25672\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNI9VSG1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25300\,
            in1 => \N__15443\,
            in2 => \_gnd_net_\,
            in3 => \N__14201\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15395\,
            in2 => \_gnd_net_\,
            in3 => \N__14354\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14351\,
            in2 => \_gnd_net_\,
            in3 => \N__14327\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15187\,
            in2 => \_gnd_net_\,
            in3 => \N__14312\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0D_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15647\,
            in2 => \_gnd_net_\,
            in3 => \N__14309\,
            lcout => \PCH_PWRGD.un2_count_1_cry_5_c_RNISK0DZ0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15137\,
            in2 => \_gnd_net_\,
            in3 => \N__14306\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14303\,
            in2 => \_gnd_net_\,
            in3 => \N__14270\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14267\,
            in2 => \_gnd_net_\,
            in3 => \N__14240\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIHF5H1_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25298\,
            in1 => \N__15599\,
            in2 => \_gnd_net_\,
            in3 => \N__14237\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15107\,
            in2 => \_gnd_net_\,
            in3 => \N__14396\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNIQOOB1_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25299\,
            in1 => \N__15541\,
            in2 => \_gnd_net_\,
            in3 => \N__14393\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIRQPB1_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25310\,
            in1 => \N__14381\,
            in2 => \_gnd_net_\,
            in3 => \N__14390\,
            lcout => \PCH_PWRGD.count_rst_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQ7_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15551\,
            in2 => \_gnd_net_\,
            in3 => \N__14387\,
            lcout => \PCH_PWRGD.un2_count_1_cry_13_c_RNIBAQZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNITURB1_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25311\,
            in1 => \N__14360\,
            in2 => \_gnd_net_\,
            in3 => \N__14384\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_0_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18139\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15731\,
            lcout => \PCH_PWRGD.N_38_f0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34740\,
            ce => \N__25582\,
            sr => \N__25373\
        );

    \PCH_PWRGD.count_RNIU7DH3_13_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14450\,
            in1 => \N__14438\,
            in2 => \_gnd_net_\,
            in3 => \N__25549\,
            lcout => \PCH_PWRGD.un2_count_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14436\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34740\,
            ce => \N__25582\,
            sr => \N__25373\
        );

    \PCH_PWRGD.count_RNI2EFH3_15_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14375\,
            in1 => \N__25550\,
            in2 => \_gnd_net_\,
            in3 => \N__14368\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => \PCH_PWRGD.countZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIU7DH3_0_13_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__25551\,
            in1 => \N__14449\,
            in2 => \N__14441\,
            in3 => \N__14437\,
            lcout => \PCH_PWRGD.count_1_i_a2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIS4CH3_12_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14423\,
            in1 => \N__14414\,
            in2 => \_gnd_net_\,
            in3 => \N__25548\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_12_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14422\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34740\,
            ce => \N__25582\,
            sr => \N__25373\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_i_i_a2_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__15686\,
            in1 => \N__15730\,
            in2 => \N__15838\,
            in3 => \N__15803\,
            lcout => \PCH_PWRGD.m6_i_i_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22316\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14508\,
            in2 => \N__20213\,
            in3 => \N__14408\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14498\,
            in2 => \N__14513\,
            in3 => \N__14405\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17046\,
            in2 => \N__14489\,
            in3 => \N__14402\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14477\,
            in2 => \N__17053\,
            in3 => \N__14399\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18583\,
            in1 => \N__14512\,
            in2 => \N__14468\,
            in3 => \N__14519\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14456\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14516\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17045\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22625\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14658\,
            in2 => \N__14546\,
            in3 => \N__14492\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15914\,
            in2 => \N__14663\,
            in3 => \N__14480\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18683\,
            in2 => \N__15905\,
            in3 => \N__14471\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15893\,
            in2 => \N__18693\,
            in3 => \N__14459\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17044\,
            in1 => \N__14662\,
            in2 => \N__16025\,
            in3 => \N__14552\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16013\,
            in2 => \_gnd_net_\,
            in3 => \N__14549\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22586\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22508\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14616\,
            in2 => \N__14675\,
            in3 => \N__14537\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14606\,
            in2 => \N__14621\,
            in3 => \N__14534\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17079\,
            in2 => \N__14597\,
            in3 => \N__14531\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14585\,
            in2 => \N__17086\,
            in3 => \N__14528\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17128\,
            in1 => \N__14620\,
            in2 => \N__14576\,
            in3 => \N__14525\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14522\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17078\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22486\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14697\,
            in2 => \N__14687\,
            in3 => \N__14600\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16070\,
            in2 => \N__14702\,
            in3 => \N__14588\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17309\,
            in2 => \N__16061\,
            in3 => \N__14579\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16046\,
            in2 => \N__17317\,
            in3 => \N__14567\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17077\,
            in1 => \N__14701\,
            in2 => \N__16037\,
            in3 => \N__14558\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14555\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17313\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_1_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101110111011"
        )
    port map (
            in0 => \N__16361\,
            in1 => \N__21245\,
            in2 => \N__24696\,
            in3 => \N__16126\,
            lcout => \POWERLED.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22463\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18695\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNIBLUJ_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__19181\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19379\,
            lcout => OPEN,
            ltout => \POWERLED.g1_i_a4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIM0E82_4_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18917\,
            in1 => \N__16362\,
            in2 => \N__14645\,
            in3 => \N__17462\,
            lcout => \POWERLED.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI9JIT_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__16367\,
            in1 => \_gnd_net_\,
            in2 => \N__17249\,
            in3 => \N__19352\,
            lcout => OPEN,
            ltout => \POWERLED.N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI4GUQ5_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__21246\,
            in1 => \N__14642\,
            in2 => \N__14636\,
            in3 => \N__14750\,
            lcout => OPEN,
            ltout => \POWERLED.pwm_out_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNIV9LA6_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__16365\,
            in1 => \_gnd_net_\,
            in2 => \N__14633\,
            in3 => \N__14735\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNI48JU1_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__16366\,
            in1 => \N__20777\,
            in2 => \_gnd_net_\,
            in3 => \N__17552\,
            lcout => \POWERLED.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001110100010"
        )
    port map (
            in0 => \N__14734\,
            in1 => \N__16364\,
            in2 => \N__14744\,
            in3 => \N__17245\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34717\,
            ce => 'H',
            sr => \N__16337\
        );

    \POWERLED.curr_state_RNI_0_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17267\,
            lcout => \POWERLED.N_2360_i\,
            ltout => \POWERLED.N_2360_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIPOU53_0_5_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14726\,
            in3 => \N__16127\,
            lcout => \POWERLED.N_660\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16465\,
            in1 => \N__16480\,
            in2 => \N__16436\,
            in3 => \N__16306\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14714\,
            in1 => \N__14720\,
            in2 => \N__14723\,
            in3 => \N__14708\,
            lcout => \VPP_VDDQ_un6_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16558\,
            in1 => \N__16399\,
            in2 => \N__16418\,
            in3 => \N__16384\,
            lcout => \VPP_VDDQ.un6_count_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16231\,
            in1 => \N__16246\,
            in2 => \N__16202\,
            in3 => \N__16261\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16216\,
            in1 => \N__16450\,
            in2 => \N__16295\,
            in3 => \N__16276\,
            lcout => \VPP_VDDQ.un6_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14918\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_0_c_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14895\,
            in2 => \N__15337\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_1_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14869\,
            in2 => \_gnd_net_\,
            in3 => \N__14858\,
            lcout => \HDA_STRAP.countZ0Z_1\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_0\,
            carryout => \HDA_STRAP.un1_count_1_cry_1\,
            clk => \N__34463\,
            ce => \N__24038\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14854\,
            in2 => \_gnd_net_\,
            in3 => \N__14840\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_1\,
            carryout => \HDA_STRAP.un1_count_1_cry_2\,
            clk => \N__34463\,
            ce => \N__24038\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14836\,
            in2 => \_gnd_net_\,
            in3 => \N__14822\,
            lcout => \HDA_STRAP.countZ0Z_3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_2\,
            carryout => \HDA_STRAP.un1_count_1_cry_3\,
            clk => \N__34463\,
            ce => \N__24038\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14812\,
            in2 => \_gnd_net_\,
            in3 => \N__14801\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_3\,
            carryout => \HDA_STRAP.un1_count_1_cry_4\,
            clk => \N__34463\,
            ce => \N__24038\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14797\,
            in2 => \_gnd_net_\,
            in3 => \N__14783\,
            lcout => \HDA_STRAP.countZ0Z_5\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_4\,
            carryout => \HDA_STRAP.un1_count_1_cry_5\,
            clk => \N__34463\,
            ce => \N__24038\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14775\,
            in2 => \_gnd_net_\,
            in3 => \N__14753\,
            lcout => \HDA_STRAP.un1_count_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_5\,
            carryout => \HDA_STRAP.un1_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15076\,
            in2 => \_gnd_net_\,
            in3 => \N__15065\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_6\,
            carryout => \HDA_STRAP.un1_count_1_cry_7\,
            clk => \N__34463\,
            ce => \N__24038\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15062\,
            in2 => \_gnd_net_\,
            in3 => \N__15038\,
            lcout => \HDA_STRAP.un1_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15035\,
            in2 => \_gnd_net_\,
            in3 => \N__15023\,
            lcout => \HDA_STRAP.countZ0Z_9\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_8\,
            carryout => \HDA_STRAP.un1_count_1_cry_9\,
            clk => \N__34404\,
            ce => \N__24036\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15019\,
            in2 => \_gnd_net_\,
            in3 => \N__14996\,
            lcout => \HDA_STRAP.un1_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_9\,
            carryout => \HDA_STRAP.un1_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14992\,
            in2 => \_gnd_net_\,
            in3 => \N__14966\,
            lcout => \HDA_STRAP.un1_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_10\,
            carryout => \HDA_STRAP.un1_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14963\,
            in2 => \_gnd_net_\,
            in3 => \N__14951\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_11\,
            carryout => \HDA_STRAP.un1_count_1_cry_12\,
            clk => \N__34404\,
            ce => \N__24036\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14948\,
            in2 => \_gnd_net_\,
            in3 => \N__14936\,
            lcout => \HDA_STRAP.countZ0Z_13\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_12\,
            carryout => \HDA_STRAP.un1_count_1_cry_13\,
            clk => \N__34404\,
            ce => \N__24036\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14933\,
            in2 => \_gnd_net_\,
            in3 => \N__14921\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_13\,
            carryout => \HDA_STRAP.un1_count_1_cry_14\,
            clk => \N__34404\,
            ce => \N__24036\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15377\,
            in2 => \_gnd_net_\,
            in3 => \N__15365\,
            lcout => \HDA_STRAP.countZ0Z_15\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_14\,
            carryout => \HDA_STRAP.un1_count_1_cry_15\,
            clk => \N__34404\,
            ce => \N__24036\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15362\,
            in2 => \_gnd_net_\,
            in3 => \N__15341\,
            lcout => \HDA_STRAP.un1_count_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__15329\,
            in1 => \N__15221\,
            in2 => \N__15271\,
            in3 => \N__15224\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34464\,
            ce => \N__24037\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_11_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__15096\,
            in1 => \N__25392\,
            in2 => \N__15209\,
            in3 => \N__15800\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__25560\,
            sr => \N__25365\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNIE92H1_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__15801\,
            in1 => \N__15167\,
            in2 => \N__25412\,
            in3 => \N__15133\,
            lcout => \PCH_PWRGD.count_rst_7\,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIMT3T1_0_7_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__25561\,
            in1 => \N__15188\,
            in2 => \N__15170\,
            in3 => \N__15146\,
            lcout => \PCH_PWRGD.count_1_i_a2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__15799\,
            in1 => \N__15166\,
            in2 => \N__25411\,
            in3 => \N__15132\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34416\,
            ce => \N__25560\,
            sr => \N__25365\
        );

    \PCH_PWRGD.count_RNIMT3T1_7_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15152\,
            in1 => \N__15145\,
            in2 => \_gnd_net_\,
            in3 => \N__25541\,
            lcout => \PCH_PWRGD.un2_count_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQ1BH3_11_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25540\,
            in1 => \N__15119\,
            in2 => \_gnd_net_\,
            in3 => \N__15113\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => \PCH_PWRGD.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIGN3T1_0_1_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001010000"
        )
    port map (
            in0 => \N__25610\,
            in1 => \N__15629\,
            in2 => \N__15437\,
            in3 => \N__25542\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIHFFK7_1_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15434\,
            in1 => \N__15428\,
            in2 => \N__15422\,
            in3 => \N__15419\,
            lcout => \PCH_PWRGD.count_1_i_a2_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI1TUH1_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15881\,
            in1 => \N__15407\,
            in2 => \_gnd_net_\,
            in3 => \N__24668\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15413\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2226_i\,
            ltout => \PCH_PWRGD.N_2226_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__15839\,
            in1 => \N__16677\,
            in2 => \N__15410\,
            in3 => \N__15780\,
            lcout => \PCH_PWRGD.curr_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI22GO8_1_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__15496\,
            in1 => \N__25663\,
            in2 => \N__15515\,
            in3 => \N__25401\,
            lcout => \PCH_PWRGD.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIHFFK7_0_1_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__25664\,
            in1 => \N__15511\,
            in2 => \_gnd_net_\,
            in3 => \N__15495\,
            lcout => \PCH_PWRGD.N_386\,
            ltout => \PCH_PWRGD.N_386_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNIA1UG1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__15571\,
            in1 => \N__25402\,
            in2 => \N__15401\,
            in3 => \N__15394\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISQ1E3_3_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__25571\,
            in1 => \_gnd_net_\,
            in2 => \N__15398\,
            in3 => \N__15557\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => \PCH_PWRGD.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_3_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15572\,
            in1 => \N__15802\,
            in2 => \N__15560\,
            in3 => \N__25399\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34699\,
            ce => \N__25570\,
            sr => \N__25400\
        );

    \PCH_PWRGD.count_2_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15463\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34540\,
            ce => \N__25562\,
            sr => \N__25366\
        );

    \PCH_PWRGD.count_RNI0BEH3_14_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__15481\,
            in1 => \N__25295\,
            in2 => \N__15473\,
            in3 => \N__25534\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => \PCH_PWRGD.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQN0E3_0_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__25537\,
            in1 => \N__15462\,
            in2 => \N__15545\,
            in3 => \N__15452\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI9P6MA_2_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15542\,
            in1 => \N__15638\,
            in2 => \N__15527\,
            in3 => \N__15524\,
            lcout => \PCH_PWRGD.count_1_i_a2_11_0\,
            ltout => \PCH_PWRGD.count_1_i_a2_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__25296\,
            in1 => \N__25662\,
            in2 => \N__15503\,
            in3 => \N__15500\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34540\,
            ce => \N__25562\,
            sr => \N__25366\
        );

    \PCH_PWRGD.count_14_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__15482\,
            in1 => \N__25297\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34540\,
            ce => \N__25562\,
            sr => \N__25366\
        );

    \PCH_PWRGD.count_RNIQN0E3_2_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25535\,
            in1 => \N__15464\,
            in2 => \_gnd_net_\,
            in3 => \N__15451\,
            lcout => \PCH_PWRGD.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIHOJLA_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15662\,
            in1 => \N__15656\,
            in2 => \_gnd_net_\,
            in3 => \N__25536\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIHI041_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15727\,
            in1 => \N__15684\,
            in2 => \_gnd_net_\,
            in3 => \N__24620\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => \PCH_PWRGD.count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI245E3_6_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__15605\,
            in1 => \N__25467\,
            in2 => \N__15650\,
            in3 => \N__15613\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => \PCH_PWRGD.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIHPOM3_0_10_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__25469\,
            in1 => \N__15591\,
            in2 => \N__15641\,
            in3 => \N__15581\,
            lcout => \PCH_PWRGD.count_1_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIGN3T1_1_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15625\,
            in1 => \N__25606\,
            in2 => \_gnd_net_\,
            in3 => \N__25586\,
            lcout => \PCH_PWRGD.un2_count_1_axb_1\,
            ltout => \PCH_PWRGD.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIHI041_1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__25404\,
            in1 => \_gnd_net_\,
            in2 => \N__15632\,
            in3 => \N__25665\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15614\,
            in2 => \_gnd_net_\,
            in3 => \N__25312\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => \N__25585\,
            sr => \N__25403\
        );

    \PCH_PWRGD.count_RNIHPOM3_10_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__25468\,
            in1 => \N__15593\,
            in2 => \_gnd_net_\,
            in3 => \N__15580\,
            lcout => \PCH_PWRGD.un2_count_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_10_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34650\,
            ce => \N__25585\,
            sr => \N__25403\
        );

    \PCH_PWRGD.curr_state_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__15831\,
            in1 => \N__15728\,
            in2 => \N__16676\,
            in3 => \N__15805\,
            lcout => \PCH_PWRGD.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34551\,
            ce => \N__21206\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI3DJU_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000000"
        )
    port map (
            in0 => \N__15866\,
            in1 => \_gnd_net_\,
            in2 => \N__30810\,
            in3 => \N__15872\,
            lcout => \PCH_PWRGD.N_670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15830\,
            lcout => \PCH_PWRGD.N_2244_i\,
            ltout => \PCH_PWRGD.N_2244_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI3DJU_0_1_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15865\,
            in2 => \N__15851\,
            in3 => \N__30800\,
            lcout => \PCH_PWRGD.N_655\,
            ltout => \PCH_PWRGD.N_655_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_0_a2_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15848\,
            in3 => \N__18124\,
            lcout => \PCH_PWRGD.curr_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI2UUH1_1_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15668\,
            in1 => \N__15845\,
            in2 => \_gnd_net_\,
            in3 => \N__24667\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__15804\,
            in1 => \N__15729\,
            in2 => \N__15689\,
            in3 => \N__15685\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34551\,
            ce => \N__21206\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__16768\,
            in1 => \N__16732\,
            in2 => \_gnd_net_\,
            in3 => \N__16697\,
            lcout => \VPP_VDDQ.N_64_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__15932\,
            in1 => \N__16702\,
            in2 => \N__16741\,
            in3 => \N__16771\,
            lcout => \VPP_VDDQ_curr_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34651\,
            ce => \N__24048\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_0_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21313\,
            in2 => \_gnd_net_\,
            in3 => \N__32021\,
            lcout => \N_626\,
            ltout => \N_626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_30_0_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__16731\,
            in1 => \N__16769\,
            in2 => \N__15938\,
            in3 => \N__24132\,
            lcout => OPEN,
            ltout => \POWERLED.G_30Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_30_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__16770\,
            in1 => \N__16733\,
            in2 => \N__15935\,
            in3 => \N__15931\,
            lcout => \G_30\,
            ltout => \G_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15917\,
            in3 => \N__24133\,
            lcout => \VPP_VDDQ.N_92_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16734\,
            in2 => \_gnd_net_\,
            in3 => \N__16698\,
            lcout => \VPP_VDDQ_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34651\,
            ce => \N__24048\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22585\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25130\,
            in2 => \N__18500\,
            in3 => \N__15908\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15992\,
            in2 => \N__16001\,
            in3 => \N__15896\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25154\,
            in2 => \N__15974\,
            in3 => \N__15884\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15956\,
            in2 => \N__25164\,
            in3 => \N__16016\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18682\,
            in1 => \N__25190\,
            in2 => \N__25207\,
            in3 => \N__16007\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16004\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__15991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25153\,
            lcout => \POWERLED.mult1_un124_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22532\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16080\,
            in2 => \N__17282\,
            in3 => \N__15983\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15980\,
            in2 => \N__16085\,
            in3 => \N__15965\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15962\,
            in2 => \N__17137\,
            in3 => \N__15950\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17133\,
            in2 => \N__15947\,
            in3 => \N__16115\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25152\,
            in1 => \N__16084\,
            in2 => \N__16112\,
            in3 => \N__16097\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16094\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16088\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17129\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22462\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16171\,
            in2 => \N__18515\,
            in3 => \N__16064\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18872\,
            in2 => \N__16175\,
            in3 => \N__16049\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18854\,
            in2 => \N__18767\,
            in3 => \N__16040\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18766\,
            in2 => \N__18833\,
            in3 => \N__16028\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17308\,
            in1 => \N__16170\,
            in2 => \N__18812\,
            in3 => \N__16181\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18788\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16178\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18762\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNISDGE_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19179\,
            in2 => \_gnd_net_\,
            in3 => \N__18915\,
            lcout => \POWERLED.count_1_5\,
            ltout => \POWERLED.count_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGTVS_5_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__24611\,
            in1 => \_gnd_net_\,
            in2 => \N__16160\,
            in3 => \N__16155\,
            lcout => \POWERLED.un1_count_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGTVS_1_5_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \N__17012\,
            in1 => \N__16157\,
            in2 => \N__16142\,
            in3 => \N__24616\,
            lcout => \POWERLED.count_RNIGTVS_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19180\,
            in2 => \_gnd_net_\,
            in3 => \N__18916\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34715\,
            ce => \N__21214\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGTVS_0_5_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__16156\,
            in1 => \N__16138\,
            in2 => \N__24676\,
            in3 => \N__19412\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIPOU53_5_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__20447\,
            in1 => \N__17461\,
            in2 => \N__16130\,
            in3 => \N__17564\,
            lcout => \POWERLED.un79_clk_100khz\,
            ltout => \POWERLED.un79_clk_100khz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__24615\,
            in1 => \_gnd_net_\,
            in2 => \N__16370\,
            in3 => \N__16363\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24156\,
            in1 => \N__16307\,
            in2 => \N__16325\,
            in3 => \N__16324\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_14_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_1_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24152\,
            in1 => \N__16294\,
            in2 => \_gnd_net_\,
            in3 => \N__16280\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_2_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24157\,
            in1 => \N__16277\,
            in2 => \_gnd_net_\,
            in3 => \N__16265\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_3_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24153\,
            in1 => \N__16262\,
            in2 => \_gnd_net_\,
            in3 => \N__16250\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_4_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24158\,
            in1 => \N__16247\,
            in2 => \_gnd_net_\,
            in3 => \N__16235\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_5_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24154\,
            in1 => \N__16232\,
            in2 => \_gnd_net_\,
            in3 => \N__16220\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_6_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24159\,
            in1 => \N__16217\,
            in2 => \_gnd_net_\,
            in3 => \N__16205\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_7_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24155\,
            in1 => \N__16201\,
            in2 => \_gnd_net_\,
            in3 => \N__16484\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__34660\,
            ce => 'H',
            sr => \N__16530\
        );

    \VPP_VDDQ.count_8_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24166\,
            in1 => \N__16481\,
            in2 => \_gnd_net_\,
            in3 => \N__16469\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.count_9_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24162\,
            in1 => \N__16466\,
            in2 => \_gnd_net_\,
            in3 => \N__16454\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.count_10_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24163\,
            in1 => \N__16451\,
            in2 => \_gnd_net_\,
            in3 => \N__16439\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.count_11_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24160\,
            in1 => \N__16435\,
            in2 => \_gnd_net_\,
            in3 => \N__16421\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.count_12_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24164\,
            in1 => \N__16417\,
            in2 => \_gnd_net_\,
            in3 => \N__16403\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.count_13_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24161\,
            in1 => \N__16400\,
            in2 => \_gnd_net_\,
            in3 => \N__16388\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.count_14_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24165\,
            in1 => \N__16385\,
            in2 => \_gnd_net_\,
            in3 => \N__16373\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__34726\,
            ce => 'H',
            sr => \N__16532\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23167\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16559\,
            in2 => \_gnd_net_\,
            in3 => \N__16562\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34718\,
            ce => \N__16547\,
            sr => \N__16531\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21482\,
            in1 => \N__20997\,
            in2 => \N__17734\,
            in3 => \N__21703\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPM861_8_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19979\,
            in2 => \N__16502\,
            in3 => \N__16499\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21485\,
            in1 => \N__21698\,
            in2 => \N__17735\,
            in3 => \N__21000\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34539\,
            ce => \N__20046\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__17717\,
            in1 => \N__21057\,
            in2 => \N__21719\,
            in3 => \N__21486\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34539\,
            ce => \N__20046\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21483\,
            in1 => \N__17716\,
            in2 => \N__21718\,
            in3 => \N__20998\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIRP961_9_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19980\,
            in2 => \N__16493\,
            in3 => \N__16490\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21484\,
            in1 => \N__20999\,
            in2 => \N__17702\,
            in3 => \N__21702\,
            lcout => \VPP_VDDQ.count_2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34539\,
            ce => \N__20046\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21538\,
            in1 => \N__21714\,
            in2 => \N__21063\,
            in3 => \N__17899\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJ48C1_14_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16784\,
            in2 => \N__16586\,
            in3 => \N__20029\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17614\,
            in1 => \N__21536\,
            in2 => \N__21062\,
            in3 => \N__21713\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIHA461_4_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16580\,
            in2 => \N__16583\,
            in3 => \N__20028\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17615\,
            in1 => \N__21537\,
            in2 => \N__21065\,
            in3 => \N__21717\,
            lcout => \VPP_VDDQ.count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34265\,
            ce => \N__20035\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21716\,
            in1 => \N__21540\,
            in2 => \N__17588\,
            in3 => \N__21047\,
            lcout => \VPP_VDDQ.count_2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34265\,
            ce => \N__20035\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21539\,
            in1 => \N__17584\,
            in2 => \N__21064\,
            in3 => \N__21715\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJD561_5_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16574\,
            in2 => \N__16568\,
            in3 => \N__20030\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIH17C1_13_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16790\,
            in1 => \N__20027\,
            in2 => \_gnd_net_\,
            in3 => \N__17840\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21709\,
            in1 => \N__21547\,
            in2 => \N__21059\,
            in3 => \N__17671\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFU5C1_12_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16796\,
            in2 => \N__16565\,
            in3 => \N__20026\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => \VPP_VDDQ.count_2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17885\,
            in1 => \N__17660\,
            in2 => \N__16799\,
            in3 => \N__17915\,
            lcout => \VPP_VDDQ.un9_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21710\,
            in1 => \N__21549\,
            in2 => \N__21060\,
            in3 => \N__17672\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34354\,
            ce => \N__20034\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21548\,
            in1 => \N__21028\,
            in2 => \N__17855\,
            in3 => \N__21712\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34354\,
            ce => \N__20034\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21711\,
            in1 => \N__21550\,
            in2 => \N__21061\,
            in3 => \N__17900\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34354\,
            ce => \N__20034\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100111101001"
        )
    port map (
            in0 => \N__16750\,
            in1 => \N__32880\,
            in2 => \N__24167\,
            in3 => \N__16778\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001111000010"
        )
    port map (
            in0 => \N__32881\,
            in1 => \N__16751\,
            in2 => \N__16712\,
            in3 => \N__16709\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__16679\,
            in1 => \N__16637\,
            in2 => \N__21248\,
            in3 => \N__16609\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21545\,
            in1 => \N__17695\,
            in2 => \N__21058\,
            in3 => \N__21708\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI4TU51_10_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16595\,
            in2 => \N__16826\,
            in3 => \N__20025\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17947\,
            in2 => \N__18173\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18003\,
            in2 => \_gnd_net_\,
            in3 => \N__16823\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18034\,
            in2 => \_gnd_net_\,
            in3 => \N__16820\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17977\,
            in2 => \_gnd_net_\,
            in3 => \N__16817\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17930\,
            in2 => \_gnd_net_\,
            in3 => \N__16814\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18345\,
            in2 => \_gnd_net_\,
            in3 => \N__16811\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17960\,
            in2 => \_gnd_net_\,
            in3 => \N__16808\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__34491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18326\,
            in2 => \_gnd_net_\,
            in3 => \N__16805\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__34491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18287\,
            in2 => \_gnd_net_\,
            in3 => \N__16802\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18301\,
            in2 => \_gnd_net_\,
            in3 => \N__16853\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18314\,
            in2 => \_gnd_net_\,
            in3 => \N__16850\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18275\,
            in2 => \_gnd_net_\,
            in3 => \N__16847\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18250\,
            in2 => \_gnd_net_\,
            in3 => \N__16844\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18236\,
            in2 => \_gnd_net_\,
            in3 => \N__16841\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18263\,
            in2 => \_gnd_net_\,
            in3 => \N__16838\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18224\,
            in2 => \_gnd_net_\,
            in3 => \N__16835\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__34550\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18185\,
            in2 => \_gnd_net_\,
            in3 => \N__16832\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_4_7_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18212\,
            in2 => \_gnd_net_\,
            in3 => \N__16829\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18199\,
            in2 => \_gnd_net_\,
            in3 => \N__16880\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18476\,
            in2 => \_gnd_net_\,
            in3 => \N__16877\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18463\,
            in2 => \_gnd_net_\,
            in3 => \N__16874\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18488\,
            in2 => \_gnd_net_\,
            in3 => \N__16871\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18449\,
            in2 => \_gnd_net_\,
            in3 => \N__16868\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18079\,
            in2 => \_gnd_net_\,
            in3 => \N__16865\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__34495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18065\,
            in2 => \_gnd_net_\,
            in3 => \N__16862\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18092\,
            in2 => \_gnd_net_\,
            in3 => \N__16859\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18104\,
            in2 => \_gnd_net_\,
            in3 => \N__16856\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16904\,
            in2 => \_gnd_net_\,
            in3 => \N__16949\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16915\,
            in2 => \_gnd_net_\,
            in3 => \N__16946\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16937\,
            in3 => \N__16943\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__16925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16940\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16933\,
            in1 => \N__16924\,
            in2 => \N__16916\,
            in3 => \N__16903\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16895\,
            in2 => \N__20135\,
            in3 => \N__19064\,
            lcout => \POWERLED.N_4842_i\,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17378\,
            in2 => \N__17395\,
            in3 => \N__22133\,
            lcout => \POWERLED.mult1_un159_sum_i_8\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17183\,
            in2 => \N__17200\,
            in3 => \N__22241\,
            lcout => \POWERLED.mult1_un152_sum_i_8\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20120\,
            in2 => \N__16889\,
            in3 => \N__18995\,
            lcout => \POWERLED.count_i_3\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17411\,
            in2 => \N__17444\,
            in3 => \N__18595\,
            lcout => \POWERLED.mult1_un138_sum_i_8\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17057\,
            in1 => \N__17024\,
            in2 => \N__17008\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_8\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19411\,
            in1 => \N__18659\,
            in2 => \N__16991\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_6\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16982\,
            in2 => \N__17150\,
            in3 => \N__20762\,
            lcout => \POWERLED.N_4841_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20519\,
            in1 => \N__16976\,
            in2 => \N__17108\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_8\,
            ltout => OPEN,
            carryin => \bfn_4_10_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16970\,
            in2 => \N__17330\,
            in3 => \N__20489\,
            lcout => \POWERLED.N_4849_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17288\,
            in2 => \N__16964\,
            in3 => \N__19280\,
            lcout => \POWERLED.count_i_10\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19250\,
            in1 => \N__16955\,
            in2 => \N__17099\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_11\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18736\,
            in1 => \N__20612\,
            in2 => \N__20629\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20582\,
            in1 => \N__17171\,
            in2 => \N__20276\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4851_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20806\,
            in1 => \N__17165\,
            in2 => \N__18533\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4855_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20843\,
            in1 => \N__17159\,
            in2 => \N__18524\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4856_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17153\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25165\,
            lcout => \POWERLED.mult1_un117_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un110_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18754\,
            lcout => \POWERLED.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17090\,
            lcout => \POWERLED.mult1_un103_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22507\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNIAVUE_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__17263\,
            in1 => \N__17365\,
            in2 => \_gnd_net_\,
            in3 => \N__17232\,
            lcout => OPEN,
            ltout => \POWERLED.N_437_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNICO541_0_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__24555\,
            in1 => \_gnd_net_\,
            in2 => \N__17270\,
            in3 => \N__17216\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => \POWERLED.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17233\,
            in2 => \N__17219\,
            in3 => \N__17361\,
            lcout => \POWERLED.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34680\,
            ce => \N__21211\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010101010"
        )
    port map (
            in0 => \N__18971\,
            in1 => \_gnd_net_\,
            in2 => \N__17366\,
            in3 => \N__24693\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34680\,
            ce => \N__21211\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUHGN_3_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__24692\,
            in1 => \N__17360\,
            in2 => \N__17210\,
            in3 => \N__18970\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIAKSS_0_2_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001111"
        )
    port map (
            in0 => \N__19013\,
            in1 => \N__17201\,
            in2 => \N__17483\,
            in3 => \N__24654\,
            lcout => \POWERLED.count_RNIAKSS_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIAKSS_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24648\,
            in1 => \N__17478\,
            in2 => \_gnd_net_\,
            in3 => \N__19010\,
            lcout => \POWERLED.un1_count_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19012\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34685\,
            ce => \N__21210\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIAKSS_1_2_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110101"
        )
    port map (
            in0 => \N__17482\,
            in1 => \N__19011\,
            in2 => \N__24691\,
            in3 => \N__18990\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIT2CB1_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011010000"
        )
    port map (
            in0 => \N__17422\,
            in1 => \N__24653\,
            in2 => \N__17465\,
            in3 => \N__18945\,
            lcout => \POWERLED.un79_clk_100khzlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_4_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18946\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34685\,
            ce => \N__21210\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIJEFE_4_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17421\,
            in1 => \N__24649\,
            in2 => \_gnd_net_\,
            in3 => \N__18944\,
            lcout => \POWERLED.un1_count_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIJEFE_0_4_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__24655\,
            in1 => \N__17443\,
            in2 => \N__18950\,
            in3 => \N__17423\,
            lcout => \POWERLED.count_RNIJEFE_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUGSJ_0_1_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100110101"
        )
    port map (
            in0 => \N__17504\,
            in1 => \N__17516\,
            in2 => \N__24690\,
            in3 => \N__17399\,
            lcout => \POWERLED.count_RNIUGSJ_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIE5D5_5_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24642\,
            in2 => \_gnd_net_\,
            in3 => \N__17350\,
            lcout => \POWERLED.count_0_sqmuxa\,
            ltout => \POWERLED.count_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIE5D5_0_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__19060\,
            in1 => \_gnd_net_\,
            in2 => \N__17333\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.count_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNITFSJ_0_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17495\,
            in2 => \N__17522\,
            in3 => \N__24643\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => \POWERLED.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIE5D5_1_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19036\,
            in2 => \N__17519\,
            in3 => \N__19141\,
            lcout => \POWERLED.count_1_1\,
            ltout => \POWERLED.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUGSJ_1_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17503\,
            in2 => \N__17510\,
            in3 => \N__24644\,
            lcout => \POWERLED.un1_count_axb_1\,
            ltout => \POWERLED.un1_count_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__19059\,
            in1 => \_gnd_net_\,
            in2 => \N__17507\,
            in3 => \N__19143\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34681\,
            ce => \N__21209\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__19142\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19058\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34681\,
            ce => \N__21209\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19196\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34725\,
            ce => \N__21215\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIALHT_11_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17489\,
            in1 => \N__24688\,
            in2 => \_gnd_net_\,
            in3 => \N__19218\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19225\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34725\,
            ce => \N__21215\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19087\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34725\,
            ce => \N__21215\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGUKT_14_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17573\,
            in1 => \N__24689\,
            in2 => \_gnd_net_\,
            in3 => \N__19192\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => \POWERLED.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19245\,
            in1 => \N__19272\,
            in2 => \N__17567\,
            in3 => \N__20823\,
            lcout => \POWERLED.un79_clk_100khzlto15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI1Q9V_10_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19418\,
            in1 => \N__24687\,
            in2 => \_gnd_net_\,
            in3 => \N__19434\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNIOF011_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__24666\,
            in1 => \N__19439\,
            in2 => \N__20485\,
            in3 => \N__19226\,
            lcout => \POWERLED.g1_i_o4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNII1MT_15_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__24665\,
            in1 => \_gnd_net_\,
            in2 => \N__19091\,
            in3 => \N__17540\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21490\,
            in1 => \N__17630\,
            in2 => \N__21694\,
            in3 => \N__21008\,
            lcout => \VPP_VDDQ.count_2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34254\,
            ce => \N__20040\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17629\,
            in1 => \N__21487\,
            in2 => \N__21052\,
            in3 => \N__21636\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID4261_2_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17534\,
            in2 => \N__17528\,
            in3 => \N__19952\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => \VPP_VDDQ.count_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_2_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19295\,
            in1 => \N__17603\,
            in2 => \N__17525\,
            in3 => \N__17747\,
            lcout => \VPP_VDDQ.un9_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21489\,
            in1 => \N__21004\,
            in2 => \N__21693\,
            in3 => \N__17866\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34254\,
            ce => \N__20040\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17867\,
            in1 => \N__21491\,
            in2 => \N__21054\,
            in3 => \N__21644\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIL79C1_15_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20041\,
            in1 => \_gnd_net_\,
            in2 => \N__17645\,
            in3 => \N__17642\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__19316\,
            in1 => \N__21488\,
            in2 => \N__21053\,
            in3 => \N__21643\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34254\,
            ce => \N__20040\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19621\,
            in2 => \N__19604\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17636\,
            in2 => \_gnd_net_\,
            in3 => \N__17621\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19294\,
            in2 => \_gnd_net_\,
            in3 => \N__17618\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19522\,
            in2 => \_gnd_net_\,
            in3 => \N__17606\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17599\,
            in2 => \_gnd_net_\,
            in3 => \N__17576\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19463\,
            in2 => \_gnd_net_\,
            in3 => \N__17753\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17783\,
            in2 => \_gnd_net_\,
            in3 => \N__17750\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17746\,
            in2 => \_gnd_net_\,
            in3 => \N__17720\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17812\,
            in2 => \_gnd_net_\,
            in3 => \N__17705\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17833\,
            in2 => \_gnd_net_\,
            in3 => \N__17684\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19871\,
            in2 => \_gnd_net_\,
            in3 => \N__17681\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17678\,
            in2 => \_gnd_net_\,
            in3 => \N__17663\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17659\,
            in2 => \_gnd_net_\,
            in3 => \N__17648\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17911\,
            in2 => \_gnd_net_\,
            in3 => \N__17888\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17884\,
            in2 => \_gnd_net_\,
            in3 => \N__17870\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21551\,
            in1 => \N__21646\,
            in2 => \N__21051\,
            in3 => \N__17851\,
            lcout => \VPP_VDDQ.count_2_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_1_7_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17834\,
            in1 => \N__17798\,
            in2 => \N__17822\,
            in3 => \N__19870\,
            lcout => \VPP_VDDQ.un9_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_0_7_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010011"
        )
    port map (
            in0 => \N__17792\,
            in1 => \N__17813\,
            in2 => \N__20039\,
            in3 => \N__17762\,
            lcout => \VPP_VDDQ.un9_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21705\,
            in1 => \N__21542\,
            in2 => \N__21055\,
            in3 => \N__17774\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => \VPP_VDDQ.count_2_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_7_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20009\,
            in1 => \_gnd_net_\,
            in2 => \N__17786\,
            in3 => \N__17761\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21706\,
            in1 => \N__21544\,
            in2 => \N__21056\,
            in3 => \N__17773\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34489\,
            ce => \N__20047\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21541\,
            in1 => \N__19599\,
            in2 => \N__21048\,
            in3 => \N__21704\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIT1QU_0_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18047\,
            in2 => \N__18053\,
            in3 => \N__20008\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21543\,
            in1 => \N__21015\,
            in2 => \N__18050\,
            in3 => \N__21707\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34489\,
            ce => \N__20047\,
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18033\,
            in1 => \N__17973\,
            in2 => \N__18004\,
            in3 => \N__18161\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__18035\,
            in1 => \N__29841\,
            in2 => \_gnd_net_\,
            in3 => \N__18041\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18017\,
            in1 => \N__17929\,
            in2 => \_gnd_net_\,
            in3 => \N__29846\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__18162\,
            in1 => \_gnd_net_\,
            in2 => \N__17948\,
            in3 => \N__29844\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__18011\,
            in1 => \_gnd_net_\,
            in2 => \N__18005\,
            in3 => \N__29845\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000010010"
        )
    port map (
            in0 => \N__17984\,
            in1 => \N__29842\,
            in2 => \N__17978\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17959\,
            in1 => \N__17943\,
            in2 => \N__18347\,
            in3 => \N__17928\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__18346\,
            in1 => \N__29843\,
            in2 => \_gnd_net_\,
            in3 => \N__18353\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18325\,
            in1 => \N__18313\,
            in2 => \N__18302\,
            in3 => \N__18286\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18274\,
            in1 => \N__18262\,
            in2 => \N__18251\,
            in3 => \N__18235\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18223\,
            in1 => \N__18211\,
            in2 => \N__18200\,
            in3 => \N__18184\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__29847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18172\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNII6BQ1_0_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001100"
        )
    port map (
            in0 => \N__25319\,
            in1 => \N__33661\,
            in2 => \N__18146\,
            in3 => \N__18125\,
            lcout => \PCH_PWRGD.curr_state_RNII6BQ1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18103\,
            in1 => \N__18091\,
            in2 => \N__18080\,
            in3 => \N__18064\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18487\,
            in1 => \N__18475\,
            in2 => \N__18464\,
            in3 => \N__18448\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22349\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18567\,
            in2 => \N__22256\,
            in3 => \N__18437\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18434\,
            in2 => \N__18572\,
            in3 => \N__18422\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18419\,
            in2 => \N__18608\,
            in3 => \N__18407\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18607\,
            in2 => \N__18404\,
            in3 => \N__18389\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21882\,
            in1 => \N__18571\,
            in2 => \N__18386\,
            in3 => \N__18371\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18368\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18356\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.VCCST_EN_i_1_i_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35131\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_12_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24505\,
            in2 => \_gnd_net_\,
            in3 => \N__29886\,
            lcout => \G_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24506\,
            in2 => \_gnd_net_\,
            in3 => \N__29887\,
            lcout => suswarn_n,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34701\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20421\,
            lcout => \POWERLED.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22742\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20684\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22397\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22427\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22531\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22396\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18618\,
            in2 => \N__18653\,
            in3 => \N__18641\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20195\,
            in2 => \N__18623\,
            in3 => \N__18638\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20296\,
            in2 => \N__20186\,
            in3 => \N__18635\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20174\,
            in2 => \N__20300\,
            in3 => \N__18632\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18730\,
            in1 => \N__18622\,
            in2 => \N__20165\,
            in3 => \N__18629\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__20312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18626\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20295\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22423\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18705\,
            in2 => \N__18884\,
            in3 => \N__18863\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18860\,
            in2 => \N__18710\,
            in3 => \N__18845\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18732\,
            in2 => \N__18842\,
            in3 => \N__18821\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18818\,
            in2 => \N__18737\,
            in3 => \N__18800\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18753\,
            in1 => \N__18709\,
            in2 => \N__18797\,
            in3 => \N__18779\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__18776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18770\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18731\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19057\,
            in2 => \N__19037\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIP7DE_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19144\,
            in1 => \_gnd_net_\,
            in2 => \N__19022\,
            in3 => \N__18998\,
            lcout => \POWERLED.count_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18994\,
            in3 => \N__18962\,
            lcout => \POWERLED.un1_count_cry_2_c_RNICZ0Z419\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2\,
            carryout => \POWERLED.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNIEQUS_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19145\,
            in1 => \_gnd_net_\,
            in2 => \N__18959\,
            in3 => \N__18932\,
            lcout => \POWERLED.count_1_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3\,
            carryout => \POWERLED.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18929\,
            in3 => \N__18896\,
            lcout => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNITFHE_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19146\,
            in1 => \_gnd_net_\,
            in2 => \N__19410\,
            in3 => \N__18893\,
            lcout => \POWERLED.count_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIUHIE_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19160\,
            in1 => \_gnd_net_\,
            in2 => \N__20754\,
            in3 => \N__18890\,
            lcout => \POWERLED.count_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIVJJE_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19147\,
            in1 => \_gnd_net_\,
            in2 => \N__20518\,
            in3 => \N__18887\,
            lcout => \POWERLED.count_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNI0MKE_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19172\,
            in1 => \_gnd_net_\,
            in2 => \N__20483\,
            in3 => \N__19283\,
            lcout => \POWERLED.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNI1OLE_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19161\,
            in1 => \_gnd_net_\,
            in2 => \N__19276\,
            in3 => \N__19253\,
            lcout => \POWERLED.count_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNI9ITC_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19173\,
            in1 => \_gnd_net_\,
            in2 => \N__19249\,
            in3 => \N__19205\,
            lcout => \POWERLED.count_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNIAKUC_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19162\,
            in1 => \_gnd_net_\,
            in2 => \N__19073\,
            in3 => \N__19202\,
            lcout => \POWERLED.count_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNIBMVC_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19174\,
            in1 => \_gnd_net_\,
            in2 => \N__20578\,
            in3 => \N__19199\,
            lcout => \POWERLED.count_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNICO0D_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__19163\,
            in1 => \_gnd_net_\,
            in2 => \N__20802\,
            in3 => \N__19184\,
            lcout => \POWERLED.count_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIDQ1D_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19175\,
            in1 => \N__20841\,
            in2 => \_gnd_net_\,
            in3 => \N__19094\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIDQ1DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICOIT_12_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20559\,
            in1 => \N__24664\,
            in2 => \_gnd_net_\,
            in3 => \N__20534\,
            lcout => \POWERLED.un1_count_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIO94T_9_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__24663\,
            in1 => \_gnd_net_\,
            in2 => \N__19457\,
            in3 => \N__19445\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19456\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34686\,
            ce => \N__21208\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19435\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34686\,
            ce => \N__21208\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNII01T_6_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19358\,
            in1 => \N__24661\,
            in2 => \_gnd_net_\,
            in3 => \N__19377\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34686\,
            ce => \N__21208\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIM63T_8_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24662\,
            in1 => \N__19325\,
            in2 => \_gnd_net_\,
            in3 => \N__19347\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19348\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34724\,
            ce => \N__21213\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__21371\,
            in1 => \N__21426\,
            in2 => \N__21349\,
            in3 => \N__21237\,
            lcout => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21480\,
            in1 => \N__19315\,
            in2 => \N__20981\,
            in3 => \N__21645\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIF7361_3_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19304\,
            in1 => \_gnd_net_\,
            in2 => \N__19298\,
            in3 => \N__19953\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__19543\,
            in1 => \N__21344\,
            in2 => \N__19820\,
            in3 => \N__19840\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34062\,
            ce => 'H',
            sr => \N__19859\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNI6JOT1_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__19841\,
            in1 => \N__19819\,
            in2 => \N__21350\,
            in3 => \N__19544\,
            lcout => OPEN,
            ltout => \VPP_VDDQ_delayed_vddq_ok_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_PWRGD_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19535\,
            in3 => \N__25114\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21428\,
            in1 => \N__19492\,
            in2 => \N__20957\,
            in3 => \N__21648\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34264\,
            ce => \N__20042\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI38QU_0_6_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110101"
        )
    port map (
            in0 => \N__19472\,
            in1 => \N__19481\,
            in2 => \N__20048\,
            in3 => \N__19526\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIOUR33_1_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19574\,
            in1 => \N__19511\,
            in2 => \N__19505\,
            in3 => \N__19502\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => \VPP_VDDQ.N_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__19493\,
            in1 => \N__20895\,
            in2 => \N__19484\,
            in3 => \N__21427\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => \VPP_VDDQ.count_2_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI38QU_6_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19934\,
            in2 => \N__19475\,
            in3 => \N__19471\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrgd_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19762\,
            in1 => \N__19739\,
            in2 => \N__19670\,
            in3 => \N__19720\,
            lcout => rsmrst_pwrgd_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_SUSn_RNIN4K9_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19669\,
            lcout => v33a_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19595\,
            in2 => \_gnd_net_\,
            in3 => \N__19622\,
            lcout => \VPP_VDDQ.count_2_RNIZ0Z_1\,
            ltout => \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_1_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21518\,
            in1 => \N__20986\,
            in2 => \N__19628\,
            in3 => \N__21632\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => \VPP_VDDQ.count_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU2QU_1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__19960\,
            in1 => \_gnd_net_\,
            in2 => \N__19625\,
            in3 => \N__19561\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__19562\,
            in1 => \N__19610\,
            in2 => \N__19603\,
            in3 => \N__20024\,
            lcout => \VPP_VDDQ.un9_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21633\,
            in1 => \N__21522\,
            in2 => \N__21049\,
            in3 => \N__19568\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34198\,
            ce => \N__20023\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__19552\,
            in1 => \N__20987\,
            in2 => \N__21546\,
            in3 => \N__21634\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34198\,
            ce => \N__20023\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21635\,
            in1 => \N__19553\,
            in2 => \N__21050\,
            in3 => \N__21523\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIDR4C1_11_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19959\,
            in2 => \N__19880\,
            in3 => \N__19877\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19834\,
            lcout => \VPP_VDDQ.N_60_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20982\,
            lcout => \VPP_VDDQ.curr_state_2_RNIZ0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111111"
        )
    port map (
            in0 => \N__21516\,
            in1 => \N__21306\,
            in2 => \N__19844\,
            in3 => \N__24630\,
            lcout => \VPP_VDDQ.N_60\,
            ltout => \VPP_VDDQ.N_60_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNINI731_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21517\,
            in2 => \N__19823\,
            in3 => \N__21238\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19805\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19796\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19787\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19778\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20108\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20099\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20087\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20075\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20060\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25852\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30417\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20148\,
            in2 => \N__20057\,
            in3 => \N__22121\,
            lcout => \G_2161\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22037\,
            in2 => \N__20153\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22122\,
            in2 => \N__22019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21992\,
            in2 => \N__22129\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20152\,
            in2 => \N__22196\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__22154\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20138\,
            lcout => \POWERLED.mult1_un166_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22236\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23822\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34426\,
            ce => \N__34002\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_52_and_i_o3_0_a2_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35443\,
            in1 => \N__32541\,
            in2 => \_gnd_net_\,
            in3 => \N__35097\,
            lcout => \POWERLED.N_600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21883\,
            lcout => \POWERLED.mult1_un145_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5QAN_0_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__35442\,
            in1 => \N__32408\,
            in2 => \_gnd_net_\,
            in3 => \N__29314\,
            lcout => \POWERLED.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22621\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22700\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20422\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22718\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22738\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20201\,
            in2 => \N__20329\,
            in3 => \N__20189\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20325\,
            in2 => \N__20255\,
            in3 => \N__20177\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20417\,
            in2 => \N__20243\,
            in3 => \N__20168\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20231\,
            in2 => \N__20423\,
            in3 => \N__20156\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20294\,
            in1 => \N__20222\,
            in2 => \N__20330\,
            in3 => \N__20306\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20438\,
            in3 => \N__20303\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => \POWERLED.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20279\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22714\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20264\,
            in2 => \N__20650\,
            in3 => \N__20246\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20646\,
            in2 => \N__20384\,
            in3 => \N__20234\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20372\,
            in2 => \N__20680\,
            in3 => \N__20225\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20676\,
            in2 => \N__20363\,
            in3 => \N__20216\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20416\,
            in1 => \N__20351\,
            in2 => \N__20651\,
            in3 => \N__20429\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20342\,
            in3 => \N__20426\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22666\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22696\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20390\,
            in2 => \N__22801\,
            in3 => \N__20375\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22797\,
            in2 => \N__21146\,
            in3 => \N__20366\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22900\,
            in2 => \N__21131\,
            in3 => \N__20354\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21116\,
            in2 => \N__22904\,
            in3 => \N__20345\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__20672\,
            in1 => \N__21104\,
            in2 => \N__22802\,
            in3 => \N__20333\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21092\,
            in2 => \_gnd_net_\,
            in3 => \N__20687\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => \POWERLED.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20654\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICOIT_0_12_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__20561\,
            in1 => \N__20633\,
            in2 => \N__20543\,
            in3 => \N__24641\,
            lcout => \POWERLED.count_RNICOIT_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20542\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34557\,
            ce => \N__21207\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_13_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20594\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34557\,
            ce => \N__21207\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIERJT_13_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20600\,
            in1 => \N__24639\,
            in2 => \_gnd_net_\,
            in3 => \N__20590\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => \POWERLED.countZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICOIT_1_12_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__24640\,
            in1 => \N__20560\,
            in2 => \N__20546\,
            in3 => \N__20535\,
            lcout => \POWERLED.un79_clk_100khzlto15_3\,
            ltout => \POWERLED.un79_clk_100khzlto15_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICOIT_5_12_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20517\,
            in1 => \N__20484\,
            in2 => \N__20450\,
            in3 => \N__20747\,
            lcout => \POWERLED.un79_clk_100khzlto15_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICOIT_4_12_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__20849\,
            in1 => \N__20842\,
            in2 => \N__20755\,
            in3 => \N__20807\,
            lcout => \POWERLED.g1_i_o4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIK32T_7_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20717\,
            in1 => \N__24631\,
            in2 => \_gnd_net_\,
            in3 => \N__20725\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34553\,
            ce => \N__21212\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI12AS_8_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__30291\,
            in1 => \N__32483\,
            in2 => \_gnd_net_\,
            in3 => \N__32960\,
            lcout => \POWERLED.un1_clk_100khz_32_and_i_0_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6SKJ1_0_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32484\,
            in1 => \N__20708\,
            in2 => \_gnd_net_\,
            in3 => \N__30290\,
            lcout => \POWERLED.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI4MHI4_4_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23870\,
            in1 => \N__33986\,
            in2 => \_gnd_net_\,
            in3 => \N__23846\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINE7B4_0_10_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__33988\,
            in1 => \_gnd_net_\,
            in2 => \N__26651\,
            in3 => \N__26696\,
            lcout => \POWERLED.un1_count_clk_2_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8SJI4_6_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20699\,
            in1 => \N__33987\,
            in2 => \_gnd_net_\,
            in3 => \N__23821\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22670\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_15_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22817\,
            in3 => \N__21134\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22844\,
            in2 => \N__22826\,
            in3 => \N__21119\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23147\,
            in2 => \N__22976\,
            in3 => \N__21107\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23148\,
            in2 => \N__22955\,
            in3 => \N__21095\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22898\,
            in1 => \N__22934\,
            in2 => \N__21077\,
            in3 => \N__21083\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21080\,
            lcout => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__22932\,
            in1 => \N__22933\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__21274\,
            in1 => \N__21372\,
            in2 => \N__21348\,
            in3 => \N__21425\,
            lcout => \VPP_VDDQ.N_53\,
            ltout => \VPP_VDDQ.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__24695\,
            in1 => \_gnd_net_\,
            in2 => \N__21068\,
            in3 => \N__21254\,
            lcout => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1\,
            ltout => \VPP_VDDQ.curr_state_2_RNIUIRHZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_a2_1_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21722\,
            in3 => \N__21647\,
            lcout => \VPP_VDDQ.N_664\,
            ltout => \VPP_VDDQ.N_664_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_0_0_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__21374\,
            in1 => \N__21481\,
            in2 => \N__21557\,
            in3 => \N__21337\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.m4_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21266\,
            in2 => \N__21554\,
            in3 => \N__24694\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_0_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__21373\,
            in1 => \N__21336\,
            in2 => \N__21278\,
            in3 => \N__21275\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34061\,
            ce => \N__21199\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_1_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21260\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34061\,
            ce => \N__21199\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_m0_0_0_a2_2_0_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__35474\,
            in1 => \N__32656\,
            in2 => \_gnd_net_\,
            in3 => \N__24675\,
            lcout => \POWERLED.N_627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI4MLK1_1_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23041\,
            in1 => \N__23257\,
            in2 => \N__23078\,
            in3 => \N__23059\,
            lcout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIVSS4_11_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23212\,
            in2 => \_gnd_net_\,
            in3 => \N__23227\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI5BM11_10_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23242\,
            in1 => \N__23272\,
            in2 => \N__21149\,
            in3 => \N__23023\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIST215_10_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24338\,
            in1 => \N__21833\,
            in2 => \N__21827\,
            in3 => \N__21824\,
            lcout => \RSMRST_PWRGD.N_662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNISRRR_15_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23182\,
            in1 => \N__23197\,
            in2 => \N__23093\,
            in3 => \N__23287\,
            lcout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30140\,
            in2 => \_gnd_net_\,
            in3 => \N__23422\,
            lcout => \POWERLED.N_613\,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21861\,
            in2 => \N__22073\,
            in3 => \N__21818\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21815\,
            in2 => \N__21866\,
            in3 => \N__21800\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21895\,
            in2 => \N__21797\,
            in3 => \N__21779\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21776\,
            in2 => \N__21899\,
            in3 => \N__21761\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22212\,
            in1 => \N__21865\,
            in2 => \N__21758\,
            in3 => \N__21740\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21737\,
            in2 => \_gnd_net_\,
            in3 => \N__21902\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21894\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__21851\,
            in1 => \N__27551\,
            in2 => \N__23342\,
            in3 => \N__33589\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34293\,
            ce => 'H',
            sr => \N__31539\
        );

    \POWERLED.dutycycle_RNIA8C49_2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__21850\,
            in2 => \N__33643\,
            in3 => \N__23338\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => \POWERLED.dutycycleZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_2_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33122\,
            in2 => \N__21842\,
            in3 => \N__32270\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110000111"
        )
    port map (
            in0 => \N__31407\,
            in1 => \N__25835\,
            in2 => \N__21839\,
            in3 => \N__31025\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_2_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21836\,
            in3 => \N__30150\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__31408\,
            in1 => \N__25836\,
            in2 => \N__30175\,
            in3 => \N__31026\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011111"
        )
    port map (
            in0 => \N__31024\,
            in1 => \_gnd_net_\,
            in2 => \N__25867\,
            in3 => \N__31406\,
            lcout => \POWERLED.un1_dutycycle_53_axb_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIER938_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__33600\,
            in1 => \N__21958\,
            in2 => \N__21971\,
            in3 => \N__23368\,
            lcout => \POWERLED.dutycycle\,
            ltout => \POWERLED.dutycycle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__27339\,
            in1 => \N__33358\,
            in2 => \N__21974\,
            in3 => \N__27415\,
            lcout => \POWERLED.dutycycle_1_0_0\,
            ltout => \POWERLED.dutycycle_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111100001000"
        )
    port map (
            in0 => \N__33602\,
            in1 => \N__23369\,
            in2 => \N__21962\,
            in3 => \N__21959\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34245\,
            ce => 'H',
            sr => \N__31538\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111011"
        )
    port map (
            in0 => \N__27340\,
            in1 => \N__33359\,
            in2 => \N__27421\,
            in3 => \N__25778\,
            lcout => \POWERLED.dutycycle_1_0_1\,
            ltout => \POWERLED.dutycycle_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNII6848_1_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111011001100"
        )
    port map (
            in0 => \N__33601\,
            in1 => \N__21928\,
            in2 => \N__21950\,
            in3 => \N__21944\,
            lcout => \dutycycle_RNII6848_0_1\,
            ltout => \dutycycle_RNII6848_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITL8S5_1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111111"
        )
    port map (
            in0 => \N__23359\,
            in1 => \N__30712\,
            in2 => \N__21947\,
            in3 => \N__33739\,
            lcout => \POWERLED.dutycycle_eena_0\,
            ltout => \POWERLED.dutycycle_eena_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__21938\,
            in1 => \N__21929\,
            in2 => \N__21932\,
            in3 => \N__33603\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34245\,
            ce => 'H',
            sr => \N__31538\
        );

    \POWERLED.func_state_RNI4R67A_1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__22082\,
            in1 => \N__24413\,
            in2 => \N__21920\,
            in3 => \N__29247\,
            lcout => \POWERLED.N_13_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_2_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111011101"
        )
    port map (
            in0 => \N__31017\,
            in1 => \N__22289\,
            in2 => \N__30204\,
            in3 => \N__30630\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m1_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__22288\,
            in1 => \N__27341\,
            in2 => \N__21905\,
            in3 => \N__29559\,
            lcout => \POWERLED_un1_dutycycle_172_m1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__25848\,
            in1 => \N__23423\,
            in2 => \N__30400\,
            in3 => \N__33108\,
            lcout => OPEN,
            ltout => \POWERLED.N_672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_5_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35576\,
            in2 => \N__22058\,
            in3 => \N__31016\,
            lcout => \dutycycle_RNI_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__30629\,
            in1 => \N__22055\,
            in2 => \N__29572\,
            in3 => \N__23480\,
            lcout => OPEN,
            ltout => \dutycycle_RNI_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNINCRN3_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__22054\,
            in1 => \N__22046\,
            in2 => \N__22040\,
            in3 => \N__25711\,
            lcout => \G_11_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_1_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25872\,
            in2 => \_gnd_net_\,
            in3 => \N__35642\,
            lcout => \N_50\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22179\,
            in2 => \N__22100\,
            in3 => \N__22031\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22028\,
            in2 => \N__22184\,
            in3 => \N__22010\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22232\,
            in2 => \N__22007\,
            in3 => \N__21986\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21983\,
            in2 => \N__22240\,
            in3 => \N__22187\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22120\,
            in1 => \N__22183\,
            in2 => \N__22169\,
            in3 => \N__22148\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__22145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22136\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30194\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_141_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29945\,
            in3 => \N__29848\,
            lcout => \G_141\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000100"
        )
    port map (
            in0 => \N__22091\,
            in1 => \N__33124\,
            in2 => \N__22552\,
            in3 => \N__32272\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIT53D6_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22262\,
            in2 => \_gnd_net_\,
            in3 => \N__29849\,
            lcout => \POWERLED.g0_7_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__30395\,
            in1 => \N__31409\,
            in2 => \_gnd_net_\,
            in3 => \N__25868\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22345\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_rep1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29872\,
            in3 => \N__29928\,
            lcout => \SUSWARN_N_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34425\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_0_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__25869\,
            in1 => \N__22274\,
            in2 => \N__35575\,
            in3 => \N__30396\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32959\,
            in1 => \N__23513\,
            in2 => \N__25907\,
            in3 => \N__28508\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_0_a2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_14_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__34969\,
            in1 => \N__22273\,
            in2 => \N__22277\,
            in3 => \N__22355\,
            lcout => \POWERLED.N_612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__32274\,
            in1 => \N__31400\,
            in2 => \_gnd_net_\,
            in3 => \N__32846\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \N__26228\,
            in1 => \N__23609\,
            in2 => \N__26108\,
            in3 => \N__23579\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32847\,
            in1 => \N__31386\,
            in2 => \_gnd_net_\,
            in3 => \N__32275\,
            lcout => \POWERLED.N_604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1O2V5_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30882\,
            in1 => \N__29939\,
            in2 => \N__32590\,
            in3 => \N__26918\,
            lcout => \POWERLED.func_state_RNI1O2V5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22309\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_8_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101011111"
        )
    port map (
            in0 => \N__31410\,
            in1 => \_gnd_net_\,
            in2 => \N__31252\,
            in3 => \N__31820\,
            lcout => OPEN,
            ltout => \POWERLED.N_9_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100001000"
        )
    port map (
            in0 => \N__33144\,
            in1 => \N__31224\,
            in2 => \N__22376\,
            in3 => \N__32831\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__31225\,
            in1 => \N__28529\,
            in2 => \N__22373\,
            in3 => \N__31821\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI14KO1_8_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__27661\,
            in1 => \N__22370\,
            in2 => \N__31254\,
            in3 => \N__31892\,
            lcout => \POWERLED.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI02AS_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27660\,
            in2 => \N__27814\,
            in3 => \N__32529\,
            lcout => \POWERLED.N_421\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_6_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011000100"
        )
    port map (
            in0 => \N__23552\,
            in1 => \N__33123\,
            in2 => \N__31826\,
            in3 => \N__32830\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_6\,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__32832\,
            in1 => \N__31230\,
            in2 => \N__22358\,
            in3 => \N__28202\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_10_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33173\,
            lcout => \POWERLED.un2_count_clk_17_0_0_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32276\,
            in2 => \N__30416\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_53_axb_0\,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30394\,
            in2 => \N__22328\,
            in3 => \N__22292\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22637\,
            in2 => \N__30195\,
            in3 => \N__22604\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22601\,
            in2 => \N__30206\,
            in3 => \N__22568\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22565\,
            in2 => \N__22553\,
            in3 => \N__22511\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31027\,
            in2 => \N__30926\,
            in3 => \N__22490\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31028\,
            in2 => \N__23435\,
            in3 => \N__22466\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28309\,
            in2 => \N__23681\,
            in3 => \N__22442\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28198\,
            in2 => \N__22439\,
            in3 => \N__22409\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22406\,
            in2 => \N__28525\,
            in3 => \N__22379\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26242\,
            in2 => \N__26171\,
            in3 => \N__22721\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34934\,
            in2 => \N__26087\,
            in3 => \N__22703\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31107\,
            in2 => \N__23693\,
            in3 => \N__22685\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26237\,
            in2 => \N__22682\,
            in3 => \N__22652\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34936\,
            in2 => \N__23666\,
            in3 => \N__22649\,
            lcout => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31085\,
            in2 => \N__23738\,
            in3 => \N__22646\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31108\,
            in2 => \N__22784\,
            in3 => \N__22643\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22640\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23002\,
            lcout => \POWERLED.un1_dutycycle_53_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22899\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34935\,
            in2 => \_gnd_net_\,
            in3 => \N__23750\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIC2MI4_8_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22775\,
            in1 => \N__33955\,
            in2 => \_gnd_net_\,
            in3 => \N__23944\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23945\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34552\,
            ce => \N__33933\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDTBQ11_7_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28589\,
            in1 => \N__29461\,
            in2 => \_gnd_net_\,
            in3 => \N__28613\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIF0DQ11_8_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__29462\,
            in1 => \_gnd_net_\,
            in2 => \N__28550\,
            in3 => \N__28574\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22768\,
            in2 => \N__22760\,
            in3 => \N__22873\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__22769\,
            in1 => \_gnd_net_\,
            in2 => \N__22877\,
            in3 => \N__22758\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22759\,
            in3 => \N__22872\,
            lcout => \POWERLED.mult1_un47_sum_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23006\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22853\,
            in3 => \N__22988\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22985\,
            in3 => \N__22967\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23163\,
            in2 => \N__22964\,
            in3 => \N__22946\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22943\,
            in2 => \N__23168\,
            in3 => \N__22919\,
            lcout => \POWERLED.mult1_un47_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_5\,
            carryout => \POWERLED.mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22916\,
            in3 => \N__22907\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22871\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__22842\,
            in1 => \N__22843\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26691\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34655\,
            ce => \N__33992\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24138\,
            in1 => \N__23092\,
            in2 => \N__24323\,
            in3 => \N__24322\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_1_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24134\,
            in1 => \N__23077\,
            in2 => \_gnd_net_\,
            in3 => \N__23063\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_2_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24139\,
            in1 => \N__23060\,
            in2 => \_gnd_net_\,
            in3 => \N__23048\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_3_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24135\,
            in1 => \N__24350\,
            in2 => \_gnd_net_\,
            in3 => \N__23045\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_4_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24140\,
            in1 => \N__23042\,
            in2 => \_gnd_net_\,
            in3 => \N__23030\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_5_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24136\,
            in1 => \N__24377\,
            in2 => \_gnd_net_\,
            in3 => \N__23027\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_6_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24141\,
            in1 => \N__23024\,
            in2 => \_gnd_net_\,
            in3 => \N__23012\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_7_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24137\,
            in1 => \N__24364\,
            in2 => \_gnd_net_\,
            in3 => \N__23009\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__34063\,
            ce => 'H',
            sr => \N__24186\
        );

    \RSMRST_PWRGD.count_8_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24148\,
            in1 => \N__23273\,
            in2 => \_gnd_net_\,
            in3 => \N__23261\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.count_9_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24144\,
            in1 => \N__23258\,
            in2 => \_gnd_net_\,
            in3 => \N__23246\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.count_10_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24145\,
            in1 => \N__23243\,
            in2 => \_gnd_net_\,
            in3 => \N__23231\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.count_11_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24142\,
            in1 => \N__23228\,
            in2 => \_gnd_net_\,
            in3 => \N__23216\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.count_12_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24146\,
            in1 => \N__23213\,
            in2 => \_gnd_net_\,
            in3 => \N__23201\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.count_13_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24143\,
            in1 => \N__23198\,
            in2 => \_gnd_net_\,
            in3 => \N__23186\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.count_14_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__24147\,
            in1 => \N__23183\,
            in2 => \_gnd_net_\,
            in3 => \N__23171\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__34286\,
            ce => 'H',
            sr => \N__24193\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23134\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23288\,
            in2 => \_gnd_net_\,
            in3 => \N__23291\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34333\,
            ce => \N__23957\,
            sr => \N__24194\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIHIN01_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000101"
        )
    port map (
            in0 => \N__25754\,
            in1 => \N__29714\,
            in2 => \N__35495\,
            in3 => \N__30559\,
            lcout => \POWERLED.N_452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.slp_s3n_signal_i_0_o2_2_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35491\,
            in2 => \_gnd_net_\,
            in3 => \N__30853\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24260\,
            in2 => \N__24302\,
            in3 => \N__29119\,
            lcout => \RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34465\,
            ce => \N__24040\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100000"
        )
    port map (
            in0 => \N__24261\,
            in1 => \N__24283\,
            in2 => \N__29130\,
            in3 => \_gnd_net_\,
            lcout => \RSMRSTn_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34465\,
            ce => \N__24040\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep2_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24262\,
            in2 => \N__24303\,
            in3 => \N__29123\,
            lcout => \RSMRSTn_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34465\,
            ce => \N__24040\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__24263\,
            in1 => \N__24284\,
            in2 => \N__29131\,
            in3 => \N__24219\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34465\,
            ce => \N__24040\,
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNI0RLU1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__32385\,
            in1 => \N__27873\,
            in2 => \N__27799\,
            in3 => \N__23329\,
            lcout => \COUNTER.tmp_0_fast_RNI0RLUZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOI5P1_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__23306\,
            in1 => \N__30033\,
            in2 => \N__23318\,
            in3 => \N__29679\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI81IE3_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__30710\,
            in1 => \_gnd_net_\,
            in2 => \N__23276\,
            in3 => \N__24877\,
            lcout => \POWERLED.N_413_N\,
            ltout => \POWERLED.N_413_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITL8S5_0_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100111011"
        )
    port map (
            in0 => \N__30390\,
            in1 => \N__33738\,
            in2 => \N__23372\,
            in3 => \N__30711\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_215_i_0_o2_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__32386\,
            in1 => \N__27874\,
            in2 => \N__27798\,
            in3 => \N__23328\,
            lcout => \POWERLED.N_430\,
            ltout => \POWERLED.N_430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITL8S5_2_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101011111"
        )
    port map (
            in0 => \N__23360\,
            in1 => \N__30709\,
            in2 => \N__23345\,
            in3 => \N__27101\,
            lcout => \POWERLED.dutycycle_eena_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_en_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__24669\,
            in1 => \N__28055\,
            in2 => \_gnd_net_\,
            in3 => \N__29873\,
            lcout => \POWERLED.func_state_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__23330\,
            in1 => \_gnd_net_\,
            in2 => \N__29888\,
            in3 => \_gnd_net_\,
            lcout => \SUSWARN_N_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_0_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001111"
        )
    port map (
            in0 => \N__24922\,
            in1 => \N__27338\,
            in2 => \N__35641\,
            in3 => \N__24718\,
            lcout => \POWERLED.un1_count_off_1_sqmuxa_8_m0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_7_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011110101111"
        )
    port map (
            in0 => \N__30002\,
            in1 => \N__24940\,
            in2 => \N__30658\,
            in3 => \N__24923\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m1_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMQ0F_1_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__27677\,
            in1 => \_gnd_net_\,
            in2 => \N__23309\,
            in3 => \N__31953\,
            lcout => \POWERLED.un1_count_off_1_sqmuxa_8_m1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNILKMD2_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23300\,
            in3 => \N__30729\,
            lcout => \N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30358\,
            in1 => \N__30997\,
            in2 => \N__33056\,
            in3 => \N__25822\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_0\,
            ltout => \POWERLED.dutycycle_RNI_6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__30625\,
            in1 => \_gnd_net_\,
            in2 => \N__23399\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_10Z0Z_0\,
            ltout => \POWERLED.dutycycle_RNI_10Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__27396\,
            in1 => \N__24929\,
            in2 => \N__23396\,
            in3 => \N__24717\,
            lcout => \POWERLED.N_676\,
            ltout => \POWERLED.N_676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI99TE_1_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32598\,
            in1 => \N__35085\,
            in2 => \N__23393\,
            in3 => \N__27676\,
            lcout => \POWERLED.N_492\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__35635\,
            in1 => \N__23449\,
            in2 => \N__29681\,
            in3 => \N__30054\,
            lcout => \POWERLED.dutycycle_RNI_13Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNILKMD2_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23560\,
            in1 => \N__25710\,
            in2 => \_gnd_net_\,
            in3 => \N__35633\,
            lcout => \G_11_i_a10_0_1\,
            ltout => \G_11_i_a10_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNI2Q8O5_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__25709\,
            in1 => \N__30089\,
            in2 => \N__23390\,
            in3 => \N__23378\,
            lcout => OPEN,
            ltout => \N_9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKJI1H_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23387\,
            in1 => \N__23486\,
            in2 => \N__23381\,
            in3 => \N__24989\,
            lcout => \POWERLED.g0_i_o4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__35634\,
            in1 => \N__23448\,
            in2 => \N__29680\,
            in3 => \N__30053\,
            lcout => \N_8_3\,
            ltout => \N_8_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIBFNS2_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__27437\,
            in1 => \N__23495\,
            in2 => \N__23489\,
            in3 => \N__25874\,
            lcout => \POWERLED.N_10_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__35636\,
            in1 => \N__23450\,
            in2 => \_gnd_net_\,
            in3 => \N__30055\,
            lcout => \POWERLED.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000001"
        )
    port map (
            in0 => \N__24958\,
            in1 => \N__25875\,
            in2 => \N__23564\,
            in3 => \N__35637\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__23474\,
            in1 => \N__24844\,
            in2 => \N__25010\,
            in3 => \N__23464\,
            lcout => \POWERLED.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34584\,
            ce => 'H',
            sr => \N__31543\
        );

    \POWERLED.dutycycle_RNIH61711_5_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001010"
        )
    port map (
            in0 => \N__24845\,
            in1 => \N__23473\,
            in2 => \N__23465\,
            in3 => \N__25000\,
            lcout => \POWERLED.dutycycleZ1Z_5\,
            ltout => \POWERLED.dutycycleZ1Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33089\,
            in1 => \N__30420\,
            in2 => \N__23453\,
            in3 => \N__25871\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__23421\,
            in1 => \N__30419\,
            in2 => \N__33145\,
            in3 => \N__25870\,
            lcout => \POWERLED.N_546\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001000"
        )
    port map (
            in0 => \N__32257\,
            in1 => \N__31415\,
            in2 => \N__31258\,
            in3 => \N__32849\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__30984\,
            in1 => \N__33088\,
            in2 => \N__23438\,
            in3 => \N__31811\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__30418\,
            in1 => \N__33128\,
            in2 => \_gnd_net_\,
            in3 => \N__23420\,
            lcout => \N_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_3_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101011101"
        )
    port map (
            in0 => \N__31414\,
            in1 => \N__33087\,
            in2 => \N__32271\,
            in3 => \N__31245\,
            lcout => \POWERLED.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__23537\,
            in1 => \N__26036\,
            in2 => \N__23531\,
            in3 => \N__29531\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34592\,
            ce => 'H',
            sr => \N__31556\
        );

    \POWERLED.dutycycle_RNI99TE_13_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__32591\,
            in1 => \N__23512\,
            in2 => \_gnd_net_\,
            in3 => \N__35126\,
            lcout => OPEN,
            ltout => \POWERLED.N_598_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI9B7B1_13_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000000010"
        )
    port map (
            in0 => \N__31887\,
            in1 => \N__27683\,
            in2 => \N__23543\,
            in3 => \N__26227\,
            lcout => OPEN,
            ltout => \POWERLED.N_450_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5FJ65_13_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010100010"
        )
    port map (
            in0 => \N__33544\,
            in1 => \N__33802\,
            in2 => \N__23540\,
            in3 => \N__30832\,
            lcout => \POWERLED.dutycycle_RNI5FJ65Z0Z_13\,
            ltout => \POWERLED.dutycycle_RNI5FJ65Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIT3QT5_13_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__23527\,
            in1 => \N__26035\,
            in2 => \N__23519\,
            in3 => \N__29530\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => \POWERLED.dutycycleZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_13_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23516\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2336_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIT70K5_8_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__23501\,
            in1 => \N__33795\,
            in2 => \N__30833\,
            in3 => \N__33543\,
            lcout => \POWERLED.dutycycle_RNIT70K5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__26050\,
            in1 => \N__28436\,
            in2 => \N__33642\,
            in3 => \N__23603\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34582\,
            ce => 'H',
            sr => \N__31589\
        );

    \POWERLED.dutycycle_RNI_6_8_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__26119\,
            in1 => \N__31217\,
            in2 => \N__32853\,
            in3 => \N__27724\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__28181\,
            in1 => \_gnd_net_\,
            in2 => \N__31809\,
            in3 => \N__28495\,
            lcout => OPEN,
            ltout => \POWERLED.un1_m2_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_8_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__32837\,
            in1 => \N__23789\,
            in2 => \N__23612\,
            in3 => \N__31219\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIGQPC6_12_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33582\,
            in1 => \N__23602\,
            in2 => \N__26051\,
            in3 => \N__28435\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => \POWERLED.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28180\,
            in2 => \N__23594\,
            in3 => \N__31769\,
            lcout => \POWERLED.un1_dutycycle_53_56_a1_2\,
            ltout => \POWERLED.un1_dutycycle_53_56_a1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_8_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__31218\,
            in1 => \N__27725\,
            in2 => \N__23591\,
            in3 => \N__32836\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_3Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_8_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23790\,
            in2 => \N__23588\,
            in3 => \N__23585\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM3TC6_15_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__23572\,
            in1 => \N__29508\,
            in2 => \N__33455\,
            in3 => \N__25930\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__25931\,
            in1 => \N__33451\,
            in2 => \N__29538\,
            in3 => \N__23573\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__31569\
        );

    \POWERLED.dutycycle_8_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__23642\,
            in1 => \N__29510\,
            in2 => \N__23654\,
            in3 => \N__25732\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34678\,
            ce => 'H',
            sr => \N__31569\
        );

    \POWERLED.dutycycle_RNI_3_10_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33134\,
            in1 => \N__31402\,
            in2 => \N__32957\,
            in3 => \N__28278\,
            lcout => \POWERLED.g0_9_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_10_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__33133\,
            in1 => \N__31215\,
            in2 => \N__28298\,
            in3 => \N__32942\,
            lcout => \POWERLED.N_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIT1OR5_8_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__29509\,
            in1 => \N__23650\,
            in2 => \N__25733\,
            in3 => \N__23641\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => \POWERLED.dutycycleZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_8_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23630\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_8\,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33132\,
            in2 => \N__23627\,
            in3 => \N__31401\,
            lcout => \POWERLED.N_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__33136\,
            in1 => \N__31404\,
            in2 => \N__31253\,
            in3 => \N__32273\,
            lcout => OPEN,
            ltout => \POWERLED.N_6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28166\,
            in1 => \N__31756\,
            in2 => \N__23624\,
            in3 => \N__32845\,
            lcout => OPEN,
            ltout => \POWERLED.N_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__23672\,
            in1 => \N__23621\,
            in2 => \N__23615\,
            in3 => \N__26315\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_15Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__28167\,
            in1 => \N__31086\,
            in2 => \N__23696\,
            in3 => \N__28511\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_6_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33135\,
            in2 => \N__31798\,
            in3 => \N__31121\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_10_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__28284\,
            in1 => \N__33137\,
            in2 => \N__23684\,
            in3 => \N__32844\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHDMC5_10_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110101"
        )
    port map (
            in0 => \N__33817\,
            in1 => \N__28214\,
            in2 => \N__27755\,
            in3 => \N__33437\,
            lcout => \POWERLED.dutycycle_RNIHDMC5Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32258\,
            in2 => \_gnd_net_\,
            in3 => \N__31226\,
            lcout => \POWERLED.N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000111100"
        )
    port map (
            in0 => \N__34937\,
            in1 => \N__26233\,
            in2 => \N__25922\,
            in3 => \N__23768\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__25949\,
            in1 => \N__23762\,
            in2 => \N__29571\,
            in3 => \N__28087\,
            lcout => \POWERLED.dutycycleZ1Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34676\,
            ce => 'H',
            sr => \N__31570\
        );

    \POWERLED.dutycycle_RNI_7_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32854\,
            in3 => \N__25899\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_12_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_13_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__25918\,
            in1 => \N__26232\,
            in2 => \N__23657\,
            in3 => \N__23792\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_8_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001001100"
        )
    port map (
            in0 => \N__23791\,
            in1 => \N__25900\,
            in2 => \N__32855\,
            in3 => \N__31244\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIK0SC6_14_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__23761\,
            in1 => \N__29555\,
            in2 => \N__28088\,
            in3 => \N__25948\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => \POWERLED.dutycycleZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_15_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__31109\,
            in1 => \_gnd_net_\,
            in2 => \N__23753\,
            in3 => \N__23749\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI4QQA4_13_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23729\,
            in1 => \N__33956\,
            in2 => \_gnd_net_\,
            in3 => \N__23908\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23909\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34656\,
            ce => \N__33935\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIFIL44_1_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__27149\,
            in1 => \N__28022\,
            in2 => \N__33669\,
            in3 => \N__23723\,
            lcout => \POWERLED.count_clk_en\,
            ltout => \POWERLED.count_clk_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI0GFI4_2_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23861\,
            in1 => \_gnd_net_\,
            in2 => \N__23711\,
            in3 => \N__23708\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23860\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34656\,
            ce => \N__33935\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23887\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34656\,
            ce => \N__33935\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI80TA4_15_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23888\,
            in1 => \N__23702\,
            in2 => \_gnd_net_\,
            in3 => \N__33957\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23842\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34656\,
            ce => \N__33935\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28676\,
            in2 => \N__34880\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34815\,
            in1 => \N__26477\,
            in2 => \_gnd_net_\,
            in3 => \N__23852\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34809\,
            in1 => \N__26342\,
            in2 => \_gnd_net_\,
            in3 => \N__23849\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34812\,
            in1 => \N__26507\,
            in2 => \_gnd_net_\,
            in3 => \N__23828\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34810\,
            in1 => \N__26763\,
            in2 => \_gnd_net_\,
            in3 => \N__23825\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34813\,
            in1 => \N__26529\,
            in2 => \_gnd_net_\,
            in3 => \N__23798\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34811\,
            in1 => \N__26406\,
            in2 => \_gnd_net_\,
            in3 => \N__23795\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34814\,
            in1 => \N__26542\,
            in2 => \_gnd_net_\,
            in3 => \N__23936\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34830\,
            in1 => \N__26749\,
            in2 => \_gnd_net_\,
            in3 => \N__23933\,
            lcout => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_8_16_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34832\,
            in1 => \N__23930\,
            in2 => \_gnd_net_\,
            in3 => \N__23918\,
            lcout => \POWERLED.count_clk_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28363\,
            in2 => \_gnd_net_\,
            in3 => \N__23915\,
            lcout => \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10\,
            carryout => \POWERLED.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34833\,
            in1 => \N__26579\,
            in2 => \_gnd_net_\,
            in3 => \N__23912\,
            lcout => \POWERLED.count_clk_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11\,
            carryout => \POWERLED.un1_count_clk_2_cry_12_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34831\,
            in1 => \N__26710\,
            in2 => \_gnd_net_\,
            in3 => \N__23897\,
            lcout => \POWERLED.count_clk_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNI6TRA4_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__34834\,
            in1 => \N__23876\,
            in2 => \_gnd_net_\,
            in3 => \N__23894\,
            lcout => \POWERLED.count_clk_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__34835\,
            in2 => \_gnd_net_\,
            in3 => \N__23891\,
            lcout => \POWERLED.count_clk_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIUMD84_0_14_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33978\,
            in1 => \N__26797\,
            in2 => \_gnd_net_\,
            in3 => \N__26571\,
            lcout => \POWERLED.un1_count_clk_2_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIN0RE1_3_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24376\,
            in1 => \N__24304\,
            in2 => \N__24365\,
            in3 => \N__24349\,
            lcout => \RSMRST_PWRGD.un1_curr_state_0_sqmuxa_0_i_a2_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24307\,
            in1 => \N__29116\,
            in2 => \_gnd_net_\,
            in3 => \N__24245\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.RSMRSTn_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__24247\,
            in1 => \_gnd_net_\,
            in2 => \N__24326\,
            in3 => \N__24221\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34399\,
            ce => \N__24028\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__24305\,
            in1 => \N__29118\,
            in2 => \_gnd_net_\,
            in3 => \N__24243\,
            lcout => \RSMRST_PWRGD.N_264_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__24246\,
            in1 => \N__29115\,
            in2 => \_gnd_net_\,
            in3 => \N__24308\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34399\,
            ce => \N__24028\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_0_1_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__24306\,
            in1 => \N__29117\,
            in2 => \_gnd_net_\,
            in3 => \N__24242\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_555_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__G_14_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__24244\,
            in1 => \N__24220\,
            in2 => \N__24197\,
            in3 => \N__24130\,
            lcout => \RSMRST_PWRGD.G_14\,
            ltout => \RSMRST_PWRGD.G_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__24131\,
            in1 => \_gnd_net_\,
            in2 => \N__23960\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_92_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIB4D36_1_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__35472\,
            in1 => \N__32676\,
            in2 => \N__26907\,
            in3 => \N__29186\,
            lcout => \POWERLED.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIOTGO_10_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__32394\,
            in1 => \N__30742\,
            in2 => \N__30577\,
            in3 => \N__29261\,
            lcout => \POWERLED.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_0_0_o2_0_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__35470\,
            in1 => \N__32674\,
            in2 => \_gnd_net_\,
            in3 => \N__27806\,
            lcout => \POWERLED.dutycycle_1_0_iv_0_0_o2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_18_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27807\,
            in1 => \N__35473\,
            in2 => \N__32681\,
            in3 => \N__32395\,
            lcout => OPEN,
            ltout => \POWERLED.N_423_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI7KPT2_1_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000000000"
        )
    port map (
            in0 => \N__30561\,
            in1 => \N__27316\,
            in2 => \N__24401\,
            in3 => \N__33369\,
            lcout => \POWERLED.N_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__32675\,
            in1 => \N__35471\,
            in2 => \_gnd_net_\,
            in3 => \N__29294\,
            lcout => OPEN,
            ltout => \POWERLED.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJ2SL7_1_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__29961\,
            in1 => \N__30277\,
            in2 => \N__24398\,
            in3 => \N__24395\,
            lcout => OPEN,
            ltout => \POWERLED.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICVMGB_1_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__24389\,
            in1 => \N__32003\,
            in2 => \N__24383\,
            in3 => \N__29889\,
            lcout => \POWERLED.g0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDNS62_1_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__29185\,
            in1 => \N__27317\,
            in2 => \N__28067\,
            in3 => \N__30560\,
            lcout => OPEN,
            ltout => \POWERLED.N_541_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6NN75_1_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__24797\,
            in1 => \N__33776\,
            in2 => \N__24380\,
            in3 => \N__24806\,
            lcout => \POWERLED.N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__24737\,
            in1 => \N__24752\,
            in2 => \N__24776\,
            in3 => \N__24782\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIP4521_1_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__24683\,
            in1 => \N__35049\,
            in2 => \N__27896\,
            in3 => \N__33364\,
            lcout => \POWERLED.N_542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8KQ72_0_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__24791\,
            in1 => \N__24824\,
            in2 => \_gnd_net_\,
            in3 => \N__29885\,
            lcout => \POWERLED.g2\,
            ltout => \POWERLED.g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIGC9OO_0_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__24763\,
            in1 => \N__24751\,
            in2 => \N__24740\,
            in3 => \N__24736\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => \POWERLED.func_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24722\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2291_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27389\,
            in1 => \N__24928\,
            in2 => \_gnd_net_\,
            in3 => \N__24719\,
            lcout => \POWERLED.func_state_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_430_i_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__32352\,
            in1 => \N__24698\,
            in2 => \N__27895\,
            in3 => \N__35050\,
            lcout => \POWERLED.N_430_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_7_o3_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35481\,
            in2 => \_gnd_net_\,
            in3 => \N__27797\,
            lcout => OPEN,
            ltout => \POWERLED.N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1PE62_1_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__27332\,
            in1 => \N__33366\,
            in2 => \N__24416\,
            in3 => \N__30539\,
            lcout => \POWERLED.N_16_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8H551_9_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110011"
        )
    port map (
            in0 => \N__32657\,
            in1 => \N__35480\,
            in2 => \N__32384\,
            in3 => \N__31822\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_e_N_3L4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_9_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111010"
        )
    port map (
            in0 => \N__31823\,
            in1 => \N__33368\,
            in2 => \N__24827\,
            in3 => \N__30271\,
            lcout => \POWERLED.dutycycle_RNI6SKJ1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.g0_8_0_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__32658\,
            in1 => \N__29960\,
            in2 => \N__35490\,
            in3 => \N__30260\,
            lcout => \POWERLED.g0_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33367\,
            in2 => \_gnd_net_\,
            in3 => \N__30540\,
            lcout => \POWERLED.N_435\,
            ltout => \POWERLED.N_435_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_1_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__33365\,
            in1 => \N__24924\,
            in2 => \N__24818\,
            in3 => \N__24815\,
            lcout => \POWERLED.func_state_1_m2s2_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__33361\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29262\,
            lcout => \POWERLED.func_state_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27348\,
            in1 => \N__27985\,
            in2 => \N__30644\,
            in3 => \N__33363\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_m1_0_a2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__32655\,
            in1 => \N__35450\,
            in2 => \N__32402\,
            in3 => \N__30264\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_0_a2_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_215_i_0_o2_0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35449\,
            in1 => \N__32654\,
            in2 => \N__35144\,
            in3 => \N__32387\,
            lcout => OPEN,
            ltout => \POWERLED.N_423_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRQ4D3_0_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100101111"
        )
    port map (
            in0 => \N__30576\,
            in1 => \N__27347\,
            in2 => \N__24800\,
            in3 => \N__28056\,
            lcout => \POWERLED.N_688\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDNFD1_1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__29710\,
            in1 => \N__33360\,
            in2 => \N__27886\,
            in3 => \N__30574\,
            lcout => \POWERLED.N_545\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.VCCST_EN_i_0_o2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__32653\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30854\,
            lcout => \VCCST_EN_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRKB61_1_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001010"
        )
    port map (
            in0 => \N__35213\,
            in1 => \N__33362\,
            in2 => \N__30797\,
            in3 => \N__30575\,
            lcout => \POWERLED.N_252_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_6_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000101"
        )
    port map (
            in0 => \N__33052\,
            in1 => \N__24944\,
            in2 => \N__33371\,
            in3 => \N__24921\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_51_and_i_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI12AS_6_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__30275\,
            in2 => \N__24881\,
            in3 => \N__33051\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_13_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI9S7D5_6_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011111111"
        )
    port map (
            in0 => \N__27254\,
            in1 => \N__24878\,
            in2 => \N__24863\,
            in3 => \N__33735\,
            lcout => \POWERLED.dutycycle_eena_13\,
            ltout => \POWERLED.dutycycle_eena_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIH1T5A_6_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__25052\,
            in1 => \N__25036\,
            in2 => \N__24860\,
            in3 => \N__33634\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNIIFNR3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__24833\,
            in1 => \N__24857\,
            in2 => \_gnd_net_\,
            in3 => \N__33736\,
            lcout => \POWERLED.dutycycle_set_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI12AS_1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__32634\,
            in1 => \N__33349\,
            in2 => \_gnd_net_\,
            in3 => \N__30276\,
            lcout => \POWERLED.func_state_RNI12ASZ0Z_1\,
            ltout => \POWERLED.func_state_RNI12ASZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHOR3_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27116\,
            in2 => \N__25055\,
            in3 => \N__33737\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3\,
            ltout => \POWERLED.un1_dutycycle_94_cry_5_c_RNIJHORZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__25046\,
            in1 => \N__25037\,
            in2 => \N__25040\,
            in3 => \N__33635\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34451\,
            ce => 'H',
            sr => \N__31563\
        );

    \POWERLED.dutycycle_RNI_1_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__30415\,
            in1 => \N__27269\,
            in2 => \N__25880\,
            in3 => \N__25028\,
            lcout => \POWERLED.N_2363_0\,
            ltout => \POWERLED.N_2363_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25022\,
            in3 => \N__35625\,
            lcout => \POWERLED.N_12_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNILKMD2_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__30311\,
            in1 => \N__25712\,
            in2 => \_gnd_net_\,
            in3 => \N__25876\,
            lcout => OPEN,
            ltout => \G_11_i_a10_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO453C_5_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__29624\,
            in1 => \N__25019\,
            in2 => \N__25013\,
            in3 => \N__25682\,
            lcout => \POWERLED.g2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_RNIGTMK4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25708\,
            in1 => \N__24983\,
            in2 => \N__24977\,
            in3 => \N__29623\,
            lcout => \N_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_17_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29641\,
            in2 => \_gnd_net_\,
            in3 => \N__29672\,
            lcout => \N_7\,
            ltout => \N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__24976\,
            in1 => \N__30310\,
            in2 => \N__24962\,
            in3 => \N__24959\,
            lcout => OPEN,
            ltout => \POWERLED.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI87EE7_5_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__29777\,
            in1 => \N__27436\,
            in2 => \N__25715\,
            in3 => \N__25707\,
            lcout => \POWERLED.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__25676\,
            in1 => \N__25631\,
            in2 => \_gnd_net_\,
            in3 => \N__25407\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34585\,
            ce => \N__25583\,
            sr => \N__25408\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25175\,
            in2 => \_gnd_net_\,
            in3 => \N__25214\,
            lcout => \POWERLED.mult1_un124_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25174\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNI8LV32_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25118\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27703\,
            lcout => \POWERLED.func_state_RNI_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30052\,
            lcout => \POWERLED.N_435_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30424\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25873\,
            in2 => \N__26005\,
            in3 => \N__25766\,
            lcout => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25983\,
            in2 => \N__30205\,
            in3 => \N__25763\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29570\,
            in1 => \N__32250\,
            in2 => \N__26006\,
            in3 => \N__25760\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25987\,
            in2 => \N__31405\,
            in3 => \N__25757\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25989\,
            in2 => \N__30996\,
            in3 => \N__25742\,
            lcout => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33106\,
            in2 => \N__26007\,
            in3 => \N__25739\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25988\,
            in2 => \N__32822\,
            in3 => \N__25736\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26008\,
            in2 => \N__31234\,
            in3 => \N__25721\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29568\,
            in1 => \N__26019\,
            in2 => \N__31807\,
            in3 => \N__25718\,
            lcout => \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29567\,
            in1 => \N__26010\,
            in2 => \N__28308\,
            in3 => \N__26057\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPE_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29569\,
            in1 => \N__26020\,
            in2 => \N__28179\,
            in3 => \N__26054\,
            lcout => \POWERLED.un1_dutycycle_94_cry_10_c_RNIKFPEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQE_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__29566\,
            in1 => \N__26009\,
            in2 => \N__28509\,
            in3 => \N__26039\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNILHQEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26021\,
            in2 => \N__26238\,
            in3 => \N__26024\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26011\,
            in2 => \N__34970\,
            in3 => \N__25937\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__31104\,
            in1 => \N__30068\,
            in2 => \_gnd_net_\,
            in3 => \N__25934\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_12_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__28272\,
            in1 => \N__28163\,
            in2 => \N__28510\,
            in3 => \N__26156\,
            lcout => \POWERLED.un1_dutycycle_53_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__28325\,
            in1 => \N__33658\,
            in2 => \N__26150\,
            in3 => \N__26137\,
            lcout => \POWERLED.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34596\,
            ce => 'H',
            sr => \N__31568\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31810\,
            in3 => \N__28162\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31773\,
            in2 => \N__28183\,
            in3 => \N__32940\,
            lcout => \POWERLED.un1_dutycycle_53_59_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6G5Q6_11_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33657\,
            in1 => \N__26146\,
            in2 => \N__26138\,
            in3 => \N__28324\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__31216\,
            in1 => \N__28491\,
            in2 => \N__26126\,
            in3 => \N__31774\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_12_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__32941\,
            in1 => \N__26093\,
            in2 => \N__26123\,
            in3 => \N__26120\,
            lcout => \POWERLED.un1_dutycycle_53_8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28271\,
            in2 => \N__28182\,
            in3 => \N__28490\,
            lcout => \POWERLED.un1_dutycycle_53_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28280\,
            in1 => \N__28165\,
            in2 => \N__34967\,
            in3 => \N__26063\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__31403\,
            in1 => \N__33107\,
            in2 => \N__32958\,
            in3 => \N__31750\,
            lcout => OPEN,
            ltout => \POWERLED.G_7_i_a5_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_10_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__28279\,
            in1 => \N__32690\,
            in2 => \N__26075\,
            in3 => \N__31220\,
            lcout => OPEN,
            ltout => \POWERLED.N_16_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_9_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__26072\,
            in1 => \N__31751\,
            in2 => \N__26066\,
            in3 => \N__26348\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITRJC6_10_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__26284\,
            in1 => \N__26269\,
            in2 => \N__26302\,
            in3 => \N__33659\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => \POWERLED.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100000"
        )
    port map (
            in0 => \N__28164\,
            in1 => \N__31752\,
            in2 => \N__26318\,
            in3 => \N__26309\,
            lcout => \POWERLED.g0_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_9_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32848\,
            in2 => \N__31797\,
            in3 => \N__32946\,
            lcout => \POWERLED.g0_9_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__26303\,
            in1 => \N__33660\,
            in2 => \N__26273\,
            in3 => \N__26285\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34708\,
            ce => 'H',
            sr => \N__31585\
        );

    \POWERLED.dutycycle_RNI_0_8_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111000000"
        )
    port map (
            in0 => \N__27740\,
            in1 => \N__32852\,
            in2 => \N__31796\,
            in3 => \N__31243\,
            lcout => \POWERLED.un1_dutycycle_53_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHDMC5_9_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111011"
        )
    port map (
            in0 => \N__26261\,
            in1 => \N__33818\,
            in2 => \N__31646\,
            in3 => \N__33436\,
            lcout => \POWERLED.dutycycle_RNIHDMC5Z0Z_9\,
            ltout => \POWERLED.dutycycle_RNIHDMC5Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_9_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__26393\,
            in1 => \N__26383\,
            in2 => \N__26246\,
            in3 => \N__33673\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34742\,
            ce => 'H',
            sr => \N__31580\
        );

    \POWERLED.dutycycle_RNI_1_10_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28274\,
            in2 => \_gnd_net_\,
            in3 => \N__31746\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_41_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000111100"
        )
    port map (
            in0 => \N__26243\,
            in1 => \N__26180\,
            in2 => \N__26174\,
            in3 => \N__31427\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKUPA6_9_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33672\,
            in1 => \N__26392\,
            in2 => \N__26384\,
            in3 => \N__26369\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_10_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28273\,
            in1 => \N__32850\,
            in2 => \N__26363\,
            in3 => \N__31242\,
            lcout => OPEN,
            ltout => \POWERLED.N_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__32851\,
            in1 => \N__31742\,
            in2 => \N__26360\,
            in3 => \N__26357\,
            lcout => \POWERLED.G_7_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINSEUC_7_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__26462\,
            in1 => \N__26408\,
            in2 => \_gnd_net_\,
            in3 => \N__26450\,
            lcout => \POWERLED.count_clk_RNINSEUCZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34737\,
            ce => \N__33936\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2JGI4_3_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26557\,
            in1 => \N__33944\,
            in2 => \_gnd_net_\,
            in3 => \N__26328\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => \POWERLED.count_clkZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__26476\,
            in1 => \N__26549\,
            in2 => \N__26336\,
            in3 => \N__26506\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_168_0_0_o2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINSEUC_6_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__26531\,
            in1 => \N__26407\,
            in2 => \N__26333\,
            in3 => \N__26449\,
            lcout => \count_clk_RNINSEUC_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2JGI4_0_3_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101100"
        )
    port map (
            in0 => \N__26330\,
            in1 => \N__26558\,
            in2 => \N__33985\,
            in3 => \N__26548\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2JGI4_1_3_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__26530\,
            in1 => \N__26505\,
            in2 => \N__26480\,
            in3 => \N__26475\,
            lcout => \POWERLED.N_625\,
            ltout => \POWERLED.N_625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINSEUC_1_10_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__26735\,
            in1 => \_gnd_net_\,
            in2 => \N__26456\,
            in3 => \N__26621\,
            lcout => \POWERLED.N_668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26417\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__33934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIE5NI4_9_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33917\,
            in1 => \N__26432\,
            in2 => \_gnd_net_\,
            in3 => \N__26440\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => \POWERLED.count_clkZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINSEUC_0_10_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__26764\,
            in1 => \N__26617\,
            in2 => \N__26453\,
            in3 => \N__28674\,
            lcout => \POWERLED.count_clk_RNINSEUC_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26441\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__33934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI6PII4_5_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26426\,
            in1 => \N__33915\,
            in2 => \_gnd_net_\,
            in3 => \N__26416\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAVKI4_7_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__33916\,
            in1 => \N__26720\,
            in2 => \_gnd_net_\,
            in3 => \N__26728\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => \POWERLED.count_clkZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__26765\,
            in1 => \N__26750\,
            in2 => \N__26738\,
            in3 => \N__28675\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_a2_8_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26729\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34677\,
            ce => \N__33934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2NPA4_12_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101100"
        )
    port map (
            in0 => \N__26591\,
            in1 => \N__26714\,
            in2 => \N__33997\,
            in3 => \N__26600\,
            lcout => \POWERLED.un2_count_clk_17_0_o2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26590\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34738\,
            ce => \N__34004\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINE7B4_10_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101100"
        )
    port map (
            in0 => \N__26692\,
            in1 => \N__26672\,
            in2 => \N__33998\,
            in3 => \N__26650\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_o2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNINSEUC_10_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26630\,
            in1 => \N__26606\,
            in2 => \N__26624\,
            in3 => \N__28364\,
            lcout => \POWERLED.count_clk_RNINSEUCZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIUMD84_14_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__33977\,
            in1 => \N__26798\,
            in2 => \N__34879\,
            in3 => \N__26573\,
            lcout => \POWERLED.un2_count_clk_17_0_o2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2NPA4_0_12_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__26599\,
            in1 => \N__33970\,
            in2 => \_gnd_net_\,
            in3 => \N__26589\,
            lcout => \POWERLED.un1_count_clk_2_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26572\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34738\,
            ce => \N__34004\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34423\,
            ce => \N__29412\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIH3EQ11_9_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29446\,
            in1 => \N__26786\,
            in2 => \_gnd_net_\,
            in3 => \N__26845\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => \POWERLED.count_offZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_10_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26980\,
            in1 => \N__28699\,
            in2 => \N__26780\,
            in3 => \N__26827\,
            lcout => \POWERLED.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIQDJO11_10_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29447\,
            in1 => \N__26777\,
            in2 => \_gnd_net_\,
            in3 => \N__26812\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34423\,
            ce => \N__29412\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI5O1N11_12_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29448\,
            in1 => \N__26771\,
            in2 => \_gnd_net_\,
            in3 => \N__26965\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26966\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34423\,
            ce => \N__29412\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI9U3N11_14_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28619\,
            in1 => \_gnd_net_\,
            in2 => \N__29460\,
            in3 => \N__28636\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28838\,
            in2 => \N__28964\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNI3666G_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28926\,
            in1 => \_gnd_net_\,
            in2 => \N__28748\,
            in3 => \N__26876\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27014\,
            in2 => \_gnd_net_\,
            in3 => \N__26873\,
            lcout => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27005\,
            in3 => \N__26870\,
            lcout => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNI6C96G_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28929\,
            in1 => \_gnd_net_\,
            in2 => \N__28763\,
            in3 => \N__26867\,
            lcout => \POWERLED.count_off_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNI7EA6G_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28927\,
            in1 => \_gnd_net_\,
            in2 => \N__28772\,
            in3 => \N__26864\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNI8GB6G_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28930\,
            in1 => \_gnd_net_\,
            in2 => \N__27236\,
            in3 => \N__26861\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNI9IC6G_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28928\,
            in1 => \_gnd_net_\,
            in2 => \N__27203\,
            in3 => \N__26858\,
            lcout => \POWERLED.count_off_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNIAKD6G_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__28931\,
            in1 => \N__26855\,
            in2 => \_gnd_net_\,
            in3 => \N__26834\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNIBME6G_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28922\,
            in1 => \_gnd_net_\,
            in2 => \N__26831\,
            in3 => \N__26801\,
            lcout => \POWERLED.count_off_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNIJSR4G_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28932\,
            in1 => \_gnd_net_\,
            in2 => \N__28700\,
            in3 => \N__26987\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNIKUS4G_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28923\,
            in1 => \_gnd_net_\,
            in2 => \N__26984\,
            in3 => \N__26954\,
            lcout => \POWERLED.count_off_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNIL0U4G_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28933\,
            in1 => \_gnd_net_\,
            in2 => \N__29042\,
            in3 => \N__26951\,
            lcout => \POWERLED.count_off_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNIM2V4G_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__28924\,
            in1 => \_gnd_net_\,
            in2 => \N__29033\,
            in3 => \N__26948\,
            lcout => \POWERLED.count_off_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIN405G_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__29009\,
            in1 => \N__28925\,
            in2 => \_gnd_net_\,
            in3 => \N__26945\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNIN405GZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBH2F5_1_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101010"
        )
    port map (
            in0 => \N__27092\,
            in1 => \N__26942\,
            in2 => \N__26930\,
            in3 => \N__33287\,
            lcout => OPEN,
            ltout => \POWERLED.N_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIVO7PG_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111011"
        )
    port map (
            in0 => \N__29327\,
            in1 => \N__26917\,
            in2 => \N__26885\,
            in3 => \N__27155\,
            lcout => \POWERLED.func_state_1_m2_1\,
            ltout => \POWERLED.func_state_1_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIFFPVI_1_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__27061\,
            in1 => \N__31954\,
            in2 => \N__26882\,
            in3 => \N__27082\,
            lcout => \POWERLED.func_state\,
            ltout => \POWERLED.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_2_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__30197\,
            in1 => \_gnd_net_\,
            in2 => \N__26879\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_426_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001010001000"
        )
    port map (
            in0 => \N__27944\,
            in1 => \N__33288\,
            in2 => \N__29260\,
            in3 => \N__27416\,
            lcout => \POWERLED.un1_func_state25_6_0_0_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIT3R01_10_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__29703\,
            in1 => \N__29241\,
            in2 => \N__30798\,
            in3 => \N__30640\,
            lcout => \POWERLED.N_562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__27062\,
            in1 => \N__31955\,
            in2 => \N__27086\,
            in3 => \N__27068\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34398\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_0_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__32668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35444\,
            lcout => \N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27026\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28917\,
            lcout => \POWERLED.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34573\,
            ce => \N__29389\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__28916\,
            in1 => \_gnd_net_\,
            in2 => \N__27047\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34573\,
            ce => \N__29389\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI7K8Q11_4_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__27053\,
            in1 => \N__28915\,
            in2 => \N__29413\,
            in3 => \N__27043\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI5H7Q11_3_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__27032\,
            in1 => \N__29385\,
            in2 => \N__28934\,
            in3 => \N__27025\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => \POWERLED.count_offZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_3_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27001\,
            in1 => \N__27235\,
            in2 => \N__27206\,
            in3 => \N__27202\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_10_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28730\,
            in1 => \N__27176\,
            in2 => \N__27164\,
            in3 => \N__28982\,
            lcout => \POWERLED.count_off_RNI_0Z0Z_10\,
            ltout => \POWERLED.count_off_RNI_0Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI8AQH_10_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27161\,
            in3 => \N__29697\,
            lcout => \POWERLED.count_off_RNI8AQHZ0Z_10\,
            ltout => \POWERLED.count_off_RNI8AQHZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIU30A4_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__30101\,
            in1 => \_gnd_net_\,
            in2 => \N__27158\,
            in3 => \N__29144\,
            lcout => \POWERLED.func_state_1_m2_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__33293\,
            in1 => \N__29240\,
            in2 => \N__27353\,
            in3 => \N__30631\,
            lcout => \POWERLED.N_494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIA61DE_10_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__27868\,
            in1 => \N__35111\,
            in2 => \N__27943\,
            in3 => \N__28384\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICU5NF_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011101100"
        )
    port map (
            in0 => \N__33292\,
            in1 => \N__27275\,
            in2 => \N__27134\,
            in3 => \N__27420\,
            lcout => \POWERLED.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__30632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32376\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_i_i_m2_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIIKO01_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110111011"
        )
    port map (
            in0 => \N__35379\,
            in1 => \N__27131\,
            in2 => \N__27119\,
            in3 => \N__29969\,
            lcout => \POWERLED.N_453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMQ0F_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__31996\,
            in1 => \N__27682\,
            in2 => \N__30660\,
            in3 => \N__31035\,
            lcout => \POWERLED.N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__33294\,
            in1 => \N__27869\,
            in2 => \N__27422\,
            in3 => \N__30639\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2O4A1_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27986\,
            in1 => \N__29189\,
            in2 => \N__30659\,
            in3 => \N__27352\,
            lcout => \POWERLED.N_490\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_3_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31352\,
            in1 => \N__30070\,
            in2 => \N__35568\,
            in3 => \N__32215\,
            lcout => \POWERLED.g1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2MQD_5_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__31018\,
            in1 => \N__35377\,
            in2 => \N__27681\,
            in3 => \N__30661\,
            lcout => \POWERLED.un1_dutycycle_172_m0_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__35378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29318\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNI2MQDZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIDASB1_6_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__30794\,
            in1 => \N__27242\,
            in2 => \N__27257\,
            in3 => \N__27611\,
            lcout => \POWERLED.dutycycle_eena_13_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_6_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33299\,
            in2 => \_gnd_net_\,
            in3 => \N__33143\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110100"
        )
    port map (
            in0 => \N__33300\,
            in1 => \N__32105\,
            in2 => \N__32249\,
            in3 => \N__30283\,
            lcout => \POWERLED.dutycycle_RNI6SKJ1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9S7D5_1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110011"
        )
    port map (
            in0 => \N__27532\,
            in1 => \N__33803\,
            in2 => \N__27587\,
            in3 => \N__33402\,
            lcout => \POWERLED.func_state_RNI9S7D5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIJ17U4_1_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__33403\,
            in1 => \N__27533\,
            in2 => \N__29603\,
            in3 => \N__33804\,
            lcout => \POWERLED.func_state_RNIJ17U4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNILC2B6_4_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__27490\,
            in1 => \N__27509\,
            in2 => \N__33671\,
            in3 => \N__27500\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNIFPUF_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__27518\,
            in1 => \N__35118\,
            in2 => \N__32647\,
            in3 => \N__27655\,
            lcout => \POWERLED.dutycycle_e_1_4\,
            ltout => \POWERLED.dutycycle_e_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33651\,
            in1 => \N__27491\,
            in2 => \N__27503\,
            in3 => \N__27499\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34741\,
            ce => 'H',
            sr => \N__31567\
        );

    \POWERLED.dutycycle_7_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__27464\,
            in1 => \N__27470\,
            in2 => \N__33670\,
            in3 => \N__27449\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34741\,
            ce => 'H',
            sr => \N__31567\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNIIV1G_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__27656\,
            in1 => \N__35119\,
            in2 => \N__32646\,
            in3 => \N__27479\,
            lcout => \POWERLED.dutycycle_e_1_7\,
            ltout => \POWERLED.dutycycle_e_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHG6Q6_7_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33644\,
            in1 => \N__27463\,
            in2 => \N__27452\,
            in3 => \N__27448\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => \POWERLED.dutycycleZ1Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101011111"
        )
    port map (
            in0 => \N__31340\,
            in1 => \_gnd_net_\,
            in2 => \N__27440\,
            in3 => \N__32192\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_25_0_tz_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__33142\,
            in1 => \N__31341\,
            in2 => \N__27728\,
            in3 => \N__31808\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2MQD_7_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__32773\,
            in1 => \N__35344\,
            in2 => \_gnd_net_\,
            in3 => \N__33298\,
            lcout => \POWERLED.dutycycle_RNI2MQDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__33297\,
            in1 => \N__29263\,
            in2 => \N__27707\,
            in3 => \N__30657\,
            lcout => \POWERLED.N_2075_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMQ0F_7_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__32063\,
            in1 => \N__32578\,
            in2 => \N__32821\,
            in3 => \N__30901\,
            lcout => \POWERLED.un1_clk_100khz_36_and_i_0_a2_1_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35345\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33289\,
            lcout => \POWERLED.func_state_RNI2MQDZ0Z_1\,
            ltout => \POWERLED.func_state_RNI2MQDZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_8_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27617\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.func_state_RNI_8Z0Z_1\,
            ltout => \POWERLED.func_state_RNI_8Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMQ0F_0_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__32579\,
            in1 => \N__30899\,
            in2 => \N__27614\,
            in3 => \N__35541\,
            lcout => \POWERLED.func_state_RNIMQ0F_0Z0Z_1\,
            ltout => \POWERLED.func_state_RNIMQ0F_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEBSB1_7_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__27602\,
            in1 => \_gnd_net_\,
            in2 => \N__27596\,
            in3 => \N__27593\,
            lcout => \POWERLED.dutycycle_RNIEBSB1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIS27B2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__27575\,
            in1 => \N__32062\,
            in2 => \N__28010\,
            in3 => \N__27563\,
            lcout => \POWERLED.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3T8L1_0_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__30809\,
            in1 => \N__28073\,
            in2 => \N__32407\,
            in3 => \N__28066\,
            lcout => \POWERLED.count_clk_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_0_0_o2_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__35325\,
            in1 => \N__32524\,
            in2 => \_gnd_net_\,
            in3 => \N__35142\,
            lcout => \POWERLED.N_443\,
            ltout => \POWERLED.N_443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIH37EG_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__27998\,
            in1 => \N__27821\,
            in2 => \N__27989\,
            in3 => \N__27902\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIS94QD_1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__27891\,
            in1 => \N__33290\,
            in2 => \N__27981\,
            in3 => \N__27927\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__33291\,
            in1 => \N__27890\,
            in2 => \N__35551\,
            in3 => \N__29264\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI02AS_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__32523\,
            in1 => \N__27815\,
            in2 => \_gnd_net_\,
            in3 => \N__35533\,
            lcout => \POWERLED.N_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_10_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__35340\,
            in1 => \N__35207\,
            in2 => \N__30296\,
            in3 => \N__28303\,
            lcout => OPEN,
            ltout => \POWERLED.N_506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_0_10_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__28302\,
            in1 => \_gnd_net_\,
            in2 => \N__27758\,
            in3 => \N__33301\,
            lcout => \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100111111"
        )
    port map (
            in0 => \N__32228\,
            in1 => \N__31387\,
            in2 => \N__33146\,
            in3 => \N__32813\,
            lcout => \POWERLED.g0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_11_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__28201\,
            in1 => \N__31869\,
            in2 => \N__32026\,
            in3 => \N__32085\,
            lcout => OPEN,
            ltout => \POWERLED.N_514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHDMC5_11_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011101"
        )
    port map (
            in0 => \N__33819\,
            in1 => \N__28103\,
            in2 => \N__28328\,
            in3 => \N__33435\,
            lcout => \POWERLED.dutycycle_RNIHDMC5Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_10_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100000000"
        )
    port map (
            in0 => \N__28304\,
            in1 => \N__31868\,
            in2 => \N__32025\,
            in3 => \N__32084\,
            lcout => \POWERLED.N_508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_11_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000110000"
        )
    port map (
            in0 => \N__30295\,
            in1 => \N__28200\,
            in2 => \N__35390\,
            in3 => \N__35208\,
            lcout => OPEN,
            ltout => \POWERLED.N_512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6SKJ1_0_11_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33302\,
            in2 => \N__28205\,
            in3 => \N__28199\,
            lcout => \POWERLED.dutycycle_RNI6SKJ1_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3T8L1_14_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__33295\,
            in1 => \N__34886\,
            in2 => \N__34968\,
            in3 => \N__33434\,
            lcout => \POWERLED.un1_clk_100khz_47_and_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_14_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000110000"
        )
    port map (
            in0 => \N__34959\,
            in1 => \N__31886\,
            in2 => \N__32093\,
            in3 => \N__32014\,
            lcout => OPEN,
            ltout => \POWERLED.N_526_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQ8KL5_14_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__33666\,
            in1 => \N__33821\,
            in2 => \N__28097\,
            in3 => \N__28094\,
            lcout => \POWERLED.dutycycle_en_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE3861_12_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__28527\,
            in1 => \N__35324\,
            in2 => \N__35148\,
            in3 => \N__35209\,
            lcout => OPEN,
            ltout => \POWERLED.N_518_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE3861_0_12_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__33296\,
            in1 => \_gnd_net_\,
            in2 => \N__28532\,
            in3 => \N__28526\,
            lcout => \POWERLED.dutycycle_RNIE3861_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_12_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000110000"
        )
    port map (
            in0 => \N__28528\,
            in1 => \N__31885\,
            in2 => \N__32092\,
            in3 => \N__32013\,
            lcout => OPEN,
            ltout => \POWERLED.N_520_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIPK9V4_12_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111011"
        )
    port map (
            in0 => \N__28445\,
            in1 => \N__33820\,
            in2 => \N__28439\,
            in3 => \N__33433\,
            lcout => \POWERLED.dutycycle_RNIPK9V4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIB15N11_15_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29458\,
            in1 => \N__28403\,
            in2 => \_gnd_net_\,
            in3 => \N__28420\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28421\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34720\,
            ce => \N__29459\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIUQMRH_1_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__32528\,
            in1 => \N__35272\,
            in2 => \N__28397\,
            in3 => \N__28373\,
            lcout => \POWERLED.func_state_RNIUQMRH_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI0KOA4_11_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__34783\,
            in1 => \N__28348\,
            in2 => \N__28337\,
            in3 => \N__33983\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34784\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34739\,
            ce => \N__33996\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34865\,
            in2 => \_gnd_net_\,
            in3 => \N__34786\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI92UF4_0_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34754\,
            in2 => \N__28685\,
            in3 => \N__33982\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => \POWERLED.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28665\,
            in2 => \N__28682\,
            in3 => \N__34782\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIA3UF4_1_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28646\,
            in2 => \N__28679\,
            in3 => \N__33984\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => \POWERLED.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34864\,
            in2 => \N__28649\,
            in3 => \N__34785\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34739\,
            ce => \N__33996\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28715\,
            lcout => \POWERLED.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__29411\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29057\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__29411\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28640\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__29411\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28603\,
            lcout => \POWERLED.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__29411\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28564\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34424\,
            ce => \N__29411\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34583\,
            ce => \N__29452\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI3E6Q11_2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28808\,
            in2 => \N__29435\,
            in3 => \N__28816\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34583\,
            ce => \N__29452\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI9N9Q11_5_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29406\,
            in1 => \N__28793\,
            in2 => \_gnd_net_\,
            in3 => \N__28801\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34583\,
            ce => \N__29452\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIBQAQ11_6_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29407\,
            in1 => \N__28787\,
            in2 => \_gnd_net_\,
            in3 => \N__28780\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => \POWERLED.count_offZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_1_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__28762\,
            in1 => \N__28747\,
            in2 => \N__28733\,
            in3 => \N__28833\,
            lcout => \POWERLED.un34_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI3L0N11_11_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__28721\,
            in1 => \_gnd_net_\,
            in2 => \N__29436\,
            in3 => \N__28711\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28940\,
            in2 => \_gnd_net_\,
            in3 => \N__28920\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34532\,
            ce => \N__29369\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI7R2N11_13_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29402\,
            in1 => \N__29066\,
            in2 => \_gnd_net_\,
            in3 => \N__29053\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => \POWERLED.count_offZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28961\,
            in1 => \N__29032\,
            in2 => \N__29012\,
            in3 => \N__29008\,
            lcout => \POWERLED.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__28919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28962\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34532\,
            ce => \N__29369\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNICU5NF_0_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__28963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28918\,
            lcout => OPEN,
            ltout => \POWERLED.count_off_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIA46B11_0_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28973\,
            in2 => \N__28967\,
            in3 => \N__29368\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => \POWERLED.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28943\,
            in3 => \N__28837\,
            lcout => \POWERLED.count_off_RNIZ0Z_1\,
            ltout => \POWERLED.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIB56B11_1_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__28921\,
            in1 => \N__28847\,
            in2 => \N__28841\,
            in3 => \N__29367\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__35447\,
            in1 => \N__32307\,
            in2 => \_gnd_net_\,
            in3 => \N__30616\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_0_a6_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_1_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__31987\,
            in1 => \N__33280\,
            in2 => \N__29594\,
            in3 => \N__29246\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_o_N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__29591\,
            in1 => \N__29582\,
            in2 => \N__29576\,
            in3 => \N__29138\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI31IBH_0_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__29573\,
            in1 => \N__29310\,
            in2 => \N__29465\,
            in3 => \N__33668\,
            lcout => \POWERLED.func_state_RNI31IBHZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIGCDO1_1_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__35446\,
            in1 => \N__32670\,
            in2 => \N__29273\,
            in3 => \N__29187\,
            lcout => \POWERLED.N_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__32669\,
            in1 => \N__35445\,
            in2 => \N__35135\,
            in3 => \N__29309\,
            lcout => \POWERLED.func_state_RNIBVNSZ0Z_0\,
            ltout => \POWERLED.func_state_RNIBVNSZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBQDR2_1_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__29245\,
            in1 => \N__29188\,
            in2 => \N__29147\,
            in3 => \N__33794\,
            lcout => \POWERLED.func_state_1_m0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a6_3_2_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__32308\,
            in1 => \N__35448\,
            in2 => \N__32680\,
            in3 => \N__35110\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35561\,
            in2 => \_gnd_net_\,
            in3 => \N__32244\,
            lcout => \POWERLED.G_11_i_o10_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_1_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__30796\,
            in1 => \N__29132\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \VCCIN_PWRGD.un10_outputZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29765\,
            in1 => \N__29759\,
            in2 => \N__29747\,
            in3 => \N__29744\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_0_o2_2_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__32375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29968\,
            lcout => \POWERLED.N_253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMQ0F_4_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110110011"
        )
    port map (
            in0 => \N__32652\,
            in1 => \N__31411\,
            in2 => \N__30905\,
            in3 => \N__35557\,
            lcout => \POWERLED.dutycycle_e_N_6L11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29995\,
            lcout => \POWERLED.func_state_RNI_6Z0Z_1\,
            ltout => \POWERLED.func_state_RNI_6Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_18_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29645\,
            in1 => \_gnd_net_\,
            in2 => \N__29630\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.N_2361_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIR8072_5_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000110101"
        )
    port map (
            in0 => \N__31046\,
            in1 => \N__30082\,
            in2 => \N__29627\,
            in3 => \N__30107\,
            lcout => \N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2MQD_4_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__35457\,
            in1 => \N__31412\,
            in2 => \_gnd_net_\,
            in3 => \N__33345\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI2MQDZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOGRS_4_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29612\,
            in2 => \N__29606\,
            in3 => \N__32082\,
            lcout => \POWERLED.dutycycle_RNIOGRSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__30069\,
            in1 => \N__31413\,
            in2 => \N__30434\,
            in3 => \N__30425\,
            lcout => \N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI3O4A1_2_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32651\,
            in1 => \N__30289\,
            in2 => \N__35476\,
            in3 => \N__30196\,
            lcout => \POWERLED.N_488\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_0_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32649\,
            in1 => \N__35127\,
            in2 => \N__35475\,
            in3 => \N__30662\,
            lcout => \POWERLED.N_540_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOGRS_5_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31020\,
            in1 => \N__29975\,
            in2 => \_gnd_net_\,
            in3 => \N__30900\,
            lcout => \POWERLED_un1_dutycycle_172_m0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30071\,
            in2 => \_gnd_net_\,
            in3 => \N__35540\,
            lcout => \POWERLED.func_state_RNI_4Z0Z_1\,
            ltout => \POWERLED.func_state_RNI_4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5DLR_5_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__31019\,
            in1 => \N__29984\,
            in2 => \N__29978\,
            in3 => \N__32648\,
            lcout => \POWERLED.dutycycle_RNI5DLRZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI7ABC3_5_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100111111"
        )
    port map (
            in0 => \N__31052\,
            in1 => \N__29958\,
            in2 => \N__29894\,
            in3 => \N__33793\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI7ABC3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNITNMH4_5_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011111100"
        )
    port map (
            in0 => \N__29959\,
            in1 => \N__30795\,
            in2 => \N__29897\,
            in3 => \N__29893\,
            lcout => \POWERLED.g2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_32_and_i_0_o2_0_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__32650\,
            in1 => \N__32377\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6RAN_5_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111110"
        )
    port map (
            in0 => \N__30663\,
            in1 => \N__35175\,
            in2 => \N__33377\,
            in3 => \N__31044\,
            lcout => \POWERLED.g1_1cf0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__32208\,
            in1 => \N__31347\,
            in2 => \_gnd_net_\,
            in3 => \N__32772\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_5_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__31348\,
            in1 => \N__31045\,
            in2 => \N__30929\,
            in3 => \N__31259\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6RAN_1_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__35176\,
            in1 => \N__33372\,
            in2 => \N__30664\,
            in3 => \N__30465\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_32_and_i_0cf0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIRKB61_0_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__30466\,
            in1 => \N__35403\,
            in2 => \N__30908\,
            in3 => \N__30898\,
            lcout => \POWERLED.un1_clk_100khz_32_and_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNILP0F_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__33376\,
            in1 => \N__30790\,
            in2 => \N__30665\,
            in3 => \N__30467\,
            lcout => \POWERLED.func_state_RNILP0FZ0Z_1\,
            ltout => \POWERLED.func_state_RNILP0FZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIHDMC5_3_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111111"
        )
    port map (
            in0 => \N__30440\,
            in1 => \N__30449\,
            in2 => \N__30443\,
            in3 => \N__33789\,
            lcout => \POWERLED.dutycycle_RNIHDMC5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100000000"
        )
    port map (
            in0 => \N__31997\,
            in1 => \N__31891\,
            in2 => \N__32248\,
            in3 => \N__32081\,
            lcout => \POWERLED.N_523\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8CJA6_3_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__31618\,
            in1 => \N__31627\,
            in2 => \N__31601\,
            in3 => \N__33662\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => \POWERLED.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_3_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__31812\,
            in1 => \N__32769\,
            in2 => \N__31631\,
            in3 => \N__31255\,
            lcout => \POWERLED.N_12_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__31600\,
            in1 => \N__31628\,
            in2 => \N__33674\,
            in3 => \N__31619\,
            lcout => \POWERLED.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34719\,
            ce => 'H',
            sr => \N__31581\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32193\,
            in2 => \_gnd_net_\,
            in3 => \N__31256\,
            lcout => OPEN,
            ltout => \POWERLED.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_6_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100111111"
        )
    port map (
            in0 => \N__32771\,
            in1 => \N__33115\,
            in2 => \N__31439\,
            in3 => \N__31813\,
            lcout => OPEN,
            ltout => \POWERLED.g0_7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_4_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110001"
        )
    port map (
            in0 => \N__31346\,
            in1 => \N__31436\,
            in2 => \N__31430\,
            in3 => \N__32900\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_3_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010111"
        )
    port map (
            in0 => \N__31345\,
            in1 => \N__32770\,
            in2 => \N__32237\,
            in3 => \N__31257\,
            lcout => \POWERLED.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE3861_15_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__31106\,
            in1 => \N__35458\,
            in2 => \N__35206\,
            in3 => \N__35143\,
            lcout => \POWERLED.N_527\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31105\,
            lcout => \POWERLED.N_2341_i\,
            ltout => \POWERLED.N_2341_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_15_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000100010"
        )
    port map (
            in0 => \N__32064\,
            in1 => \N__31864\,
            in2 => \N__33824\,
            in3 => \N__32007\,
            lcout => OPEN,
            ltout => \POWERLED.N_529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQ8KL5_1_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__33152\,
            in1 => \N__33811\,
            in2 => \N__33677\,
            in3 => \N__33667\,
            lcout => \POWERLED.dutycycle_en_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI3T8L1_1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__33432\,
            in1 => \N__33370\,
            in2 => \N__33182\,
            in3 => \N__33169\,
            lcout => \POWERLED.un1_clk_100khz_48_and_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011111111"
        )
    port map (
            in0 => \N__33141\,
            in1 => \N__32814\,
            in2 => \N__31825\,
            in3 => \N__32953\,
            lcout => \POWERLED.g0_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__32008\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32894\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_3_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32229\,
            in2 => \_gnd_net_\,
            in3 => \N__32812\,
            lcout => \POWERLED.G_7_i_o5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI8H551_3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110011"
        )
    port map (
            in0 => \N__32645\,
            in1 => \N__35409\,
            in2 => \N__32406\,
            in3 => \N__32230\,
            lcout => \POWERLED.dutycycle_e_N_3L4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIMSAB1_9_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001010"
        )
    port map (
            in0 => \N__32083\,
            in1 => \N__32012\,
            in2 => \N__31884\,
            in3 => \N__31824\,
            lcout => \POWERLED.N_505\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_6_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35629\,
            lcout => \POWERLED.N_412_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE3861_14_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__35351\,
            in1 => \N__35194\,
            in2 => \N__35153\,
            in3 => \N__34960\,
            lcout => \POWERLED.N_524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34872\,
            in2 => \_gnd_net_\,
            in3 => \N__34808\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__34716\,
            ce => \N__34003\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
