-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 13 2022 16:56:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : in std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : in std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : in std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__37129\ : std_logic;
signal \N__37128\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37118\ : std_logic;
signal \N__37117\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37091\ : std_logic;
signal \N__37090\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37073\ : std_logic;
signal \N__37072\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37055\ : std_logic;
signal \N__37054\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37046\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37036\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37027\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37009\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37001\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36992\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36983\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36973\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36965\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36963\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36946\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36937\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36928\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36919\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36892\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36884\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36866\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36857\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36848\ : std_logic;
signal \N__36847\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36820\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36818\ : std_logic;
signal \N__36817\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36802\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36793\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36783\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36778\ : std_logic;
signal \N__36775\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36772\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36765\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36760\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36732\ : std_logic;
signal \N__36727\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36706\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36699\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36693\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36663\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36660\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36656\ : std_logic;
signal \N__36655\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36629\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36622\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36619\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36617\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36615\ : std_logic;
signal \N__36614\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36608\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36605\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36601\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36593\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36590\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36585\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36583\ : std_logic;
signal \N__36582\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36404\ : std_logic;
signal \N__36403\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36400\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36376\ : std_logic;
signal \N__36373\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36360\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36357\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36352\ : std_logic;
signal \N__36349\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36343\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36292\ : std_logic;
signal \N__36289\ : std_logic;
signal \N__36286\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36270\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36266\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36232\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36226\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36211\ : std_logic;
signal \N__36208\ : std_logic;
signal \N__36205\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36194\ : std_logic;
signal \N__36191\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36187\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36146\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36133\ : std_logic;
signal \N__36130\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36128\ : std_logic;
signal \N__36125\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36119\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36037\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36031\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36028\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35984\ : std_logic;
signal \N__35975\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35969\ : std_logic;
signal \N__35966\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35932\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35929\ : std_logic;
signal \N__35926\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35924\ : std_logic;
signal \N__35923\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35918\ : std_logic;
signal \N__35917\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35893\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35891\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35887\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35870\ : std_logic;
signal \N__35867\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35837\ : std_logic;
signal \N__35834\ : std_logic;
signal \N__35831\ : std_logic;
signal \N__35828\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35816\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35797\ : std_logic;
signal \N__35794\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35782\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35764\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35746\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35744\ : std_logic;
signal \N__35741\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35731\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35715\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35684\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35654\ : std_logic;
signal \N__35653\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35647\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35630\ : std_logic;
signal \N__35627\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35593\ : std_logic;
signal \N__35590\ : std_logic;
signal \N__35587\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35571\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35566\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35548\ : std_logic;
signal \N__35545\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35526\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35517\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35488\ : std_logic;
signal \N__35485\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35447\ : std_logic;
signal \N__35444\ : std_logic;
signal \N__35443\ : std_logic;
signal \N__35440\ : std_logic;
signal \N__35435\ : std_logic;
signal \N__35432\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35419\ : std_logic;
signal \N__35416\ : std_logic;
signal \N__35413\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35404\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35389\ : std_logic;
signal \N__35386\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35382\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35378\ : std_logic;
signal \N__35377\ : std_logic;
signal \N__35374\ : std_logic;
signal \N__35369\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35328\ : std_logic;
signal \N__35323\ : std_logic;
signal \N__35320\ : std_logic;
signal \N__35317\ : std_logic;
signal \N__35314\ : std_logic;
signal \N__35311\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35299\ : std_logic;
signal \N__35296\ : std_logic;
signal \N__35293\ : std_logic;
signal \N__35290\ : std_logic;
signal \N__35287\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35281\ : std_logic;
signal \N__35278\ : std_logic;
signal \N__35275\ : std_logic;
signal \N__35272\ : std_logic;
signal \N__35269\ : std_logic;
signal \N__35266\ : std_logic;
signal \N__35263\ : std_logic;
signal \N__35260\ : std_logic;
signal \N__35257\ : std_logic;
signal \N__35254\ : std_logic;
signal \N__35251\ : std_logic;
signal \N__35248\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35213\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35175\ : std_logic;
signal \N__35172\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35080\ : std_logic;
signal \N__35077\ : std_logic;
signal \N__35074\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35068\ : std_logic;
signal \N__35065\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35058\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35046\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35043\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35039\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35024\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35016\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35003\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34990\ : std_logic;
signal \N__34987\ : std_logic;
signal \N__34984\ : std_logic;
signal \N__34981\ : std_logic;
signal \N__34978\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34955\ : std_logic;
signal \N__34952\ : std_logic;
signal \N__34949\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34921\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34912\ : std_logic;
signal \N__34909\ : std_logic;
signal \N__34906\ : std_logic;
signal \N__34903\ : std_logic;
signal \N__34900\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34892\ : std_logic;
signal \N__34889\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34883\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34871\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34854\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34834\ : std_logic;
signal \N__34831\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34819\ : std_logic;
signal \N__34816\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34810\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34798\ : std_logic;
signal \N__34795\ : std_logic;
signal \N__34792\ : std_logic;
signal \N__34789\ : std_logic;
signal \N__34786\ : std_logic;
signal \N__34783\ : std_logic;
signal \N__34780\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34753\ : std_logic;
signal \N__34750\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34738\ : std_logic;
signal \N__34735\ : std_logic;
signal \N__34732\ : std_logic;
signal \N__34729\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34721\ : std_logic;
signal \N__34718\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34711\ : std_logic;
signal \N__34702\ : std_logic;
signal \N__34697\ : std_logic;
signal \N__34694\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34675\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34669\ : std_logic;
signal \N__34666\ : std_logic;
signal \N__34663\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34661\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34607\ : std_logic;
signal \N__34600\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34591\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34582\ : std_logic;
signal \N__34579\ : std_logic;
signal \N__34576\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34558\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34549\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34523\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34513\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34501\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34495\ : std_logic;
signal \N__34492\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34477\ : std_logic;
signal \N__34474\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34468\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34459\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34441\ : std_logic;
signal \N__34438\ : std_logic;
signal \N__34437\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34423\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34410\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34378\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34325\ : std_logic;
signal \N__34322\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34316\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34288\ : std_logic;
signal \N__34285\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34279\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34270\ : std_logic;
signal \N__34267\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34249\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34242\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34214\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34198\ : std_logic;
signal \N__34195\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34177\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34171\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34144\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34108\ : std_logic;
signal \N__34105\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34078\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34073\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34054\ : std_logic;
signal \N__34051\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34018\ : std_logic;
signal \N__34015\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33955\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33904\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33892\ : std_logic;
signal \N__33889\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33883\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33870\ : std_logic;
signal \N__33867\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33859\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33847\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33814\ : std_logic;
signal \N__33811\ : std_logic;
signal \N__33808\ : std_logic;
signal \N__33805\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33797\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33785\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33782\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33771\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33746\ : std_logic;
signal \N__33743\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33735\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33653\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33647\ : std_logic;
signal \N__33644\ : std_logic;
signal \N__33641\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33633\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33629\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33625\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33617\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33604\ : std_logic;
signal \N__33601\ : std_logic;
signal \N__33598\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33596\ : std_logic;
signal \N__33595\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33566\ : std_logic;
signal \N__33563\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33544\ : std_logic;
signal \N__33529\ : std_logic;
signal \N__33526\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33487\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33457\ : std_logic;
signal \N__33454\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33448\ : std_logic;
signal \N__33445\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33424\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33352\ : std_logic;
signal \N__33349\ : std_logic;
signal \N__33346\ : std_logic;
signal \N__33343\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33329\ : std_logic;
signal \N__33326\ : std_logic;
signal \N__33323\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33320\ : std_logic;
signal \N__33317\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33205\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33199\ : std_logic;
signal \N__33196\ : std_logic;
signal \N__33193\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33113\ : std_logic;
signal \N__33110\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33086\ : std_logic;
signal \N__33083\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33050\ : std_logic;
signal \N__33047\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33028\ : std_logic;
signal \N__33025\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33014\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33001\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32969\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32955\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32944\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32939\ : std_logic;
signal \N__32936\ : std_logic;
signal \N__32933\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32923\ : std_logic;
signal \N__32920\ : std_logic;
signal \N__32917\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32869\ : std_logic;
signal \N__32866\ : std_logic;
signal \N__32863\ : std_logic;
signal \N__32860\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32841\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32837\ : std_logic;
signal \N__32834\ : std_logic;
signal \N__32831\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32795\ : std_logic;
signal \N__32788\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32776\ : std_logic;
signal \N__32773\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32760\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32731\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32725\ : std_logic;
signal \N__32722\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32700\ : std_logic;
signal \N__32695\ : std_logic;
signal \N__32692\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32670\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32657\ : std_logic;
signal \N__32654\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32648\ : std_logic;
signal \N__32645\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32587\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32578\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32570\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32530\ : std_logic;
signal \N__32521\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32519\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32498\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32475\ : std_logic;
signal \N__32472\ : std_logic;
signal \N__32469\ : std_logic;
signal \N__32468\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32456\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32446\ : std_logic;
signal \N__32443\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32438\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32417\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32407\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32393\ : std_logic;
signal \N__32390\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32374\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32365\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32354\ : std_logic;
signal \N__32351\ : std_logic;
signal \N__32348\ : std_logic;
signal \N__32345\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32332\ : std_logic;
signal \N__32329\ : std_logic;
signal \N__32326\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32254\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32248\ : std_logic;
signal \N__32245\ : std_logic;
signal \N__32242\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32236\ : std_logic;
signal \N__32233\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32174\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32150\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32143\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32141\ : std_logic;
signal \N__32140\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32135\ : std_logic;
signal \N__32132\ : std_logic;
signal \N__32129\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32093\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32090\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32015\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31999\ : std_logic;
signal \N__31996\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31977\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31969\ : std_logic;
signal \N__31966\ : std_logic;
signal \N__31963\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31940\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31927\ : std_logic;
signal \N__31924\ : std_logic;
signal \N__31921\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31913\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31910\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31907\ : std_logic;
signal \N__31900\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31865\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31849\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31823\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31813\ : std_logic;
signal \N__31810\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31774\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31762\ : std_logic;
signal \N__31759\ : std_logic;
signal \N__31756\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31706\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31690\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31681\ : std_logic;
signal \N__31678\ : std_logic;
signal \N__31673\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31595\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31543\ : std_logic;
signal \N__31540\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31519\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31511\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31493\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31481\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31466\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31432\ : std_logic;
signal \N__31429\ : std_logic;
signal \N__31426\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31371\ : std_logic;
signal \N__31368\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31362\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31354\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31285\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31279\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31247\ : std_logic;
signal \N__31244\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31192\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31132\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31085\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31059\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31013\ : std_logic;
signal \N__31010\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30982\ : std_logic;
signal \N__30981\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30979\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30976\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30973\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30958\ : std_logic;
signal \N__30957\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30952\ : std_logic;
signal \N__30951\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30887\ : std_logic;
signal \N__30884\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30855\ : std_logic;
signal \N__30854\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30845\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30842\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30821\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30815\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30812\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30715\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30710\ : std_logic;
signal \N__30709\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30697\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30665\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30661\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30655\ : std_logic;
signal \N__30644\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30634\ : std_logic;
signal \N__30629\ : std_logic;
signal \N__30626\ : std_logic;
signal \N__30617\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30587\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30562\ : std_logic;
signal \N__30559\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30536\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30521\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30457\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30445\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30437\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30416\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30398\ : std_logic;
signal \N__30395\ : std_logic;
signal \N__30392\ : std_logic;
signal \N__30389\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30370\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30352\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30343\ : std_logic;
signal \N__30340\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30331\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30314\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30287\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30283\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30266\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30249\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30230\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30190\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30130\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30124\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30088\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30086\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30070\ : std_logic;
signal \N__30067\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30051\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30031\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30025\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29992\ : std_logic;
signal \N__29989\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29956\ : std_logic;
signal \N__29953\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29947\ : std_logic;
signal \N__29944\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29906\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29839\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29836\ : std_logic;
signal \N__29833\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29806\ : std_logic;
signal \N__29803\ : std_logic;
signal \N__29800\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29774\ : std_logic;
signal \N__29771\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29761\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29746\ : std_logic;
signal \N__29743\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29732\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29726\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29713\ : std_logic;
signal \N__29710\ : std_logic;
signal \N__29707\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29560\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29542\ : std_logic;
signal \N__29539\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29534\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29506\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29495\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29446\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29426\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29400\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29379\ : std_logic;
signal \N__29376\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29330\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29323\ : std_logic;
signal \N__29320\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29230\ : std_logic;
signal \N__29227\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29201\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29164\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29116\ : std_logic;
signal \N__29115\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29101\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29088\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29068\ : std_logic;
signal \N__29065\ : std_logic;
signal \N__29062\ : std_logic;
signal \N__29059\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29053\ : std_logic;
signal \N__29050\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29047\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29015\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28960\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28939\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28918\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28872\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28837\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28822\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28814\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28754\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28744\ : std_logic;
signal \N__28741\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28696\ : std_logic;
signal \N__28693\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28687\ : std_logic;
signal \N__28684\ : std_logic;
signal \N__28681\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28666\ : std_logic;
signal \N__28663\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28579\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28522\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28513\ : std_logic;
signal \N__28510\ : std_logic;
signal \N__28507\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28499\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28459\ : std_logic;
signal \N__28456\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28447\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28442\ : std_logic;
signal \N__28439\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28426\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28396\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28342\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28309\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28201\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28139\ : std_logic;
signal \N__28136\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28126\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28120\ : std_logic;
signal \N__28117\ : std_logic;
signal \N__28114\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28084\ : std_logic;
signal \N__28081\ : std_logic;
signal \N__28078\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28045\ : std_logic;
signal \N__28042\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28019\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28009\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27975\ : std_logic;
signal \N__27972\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27958\ : std_logic;
signal \N__27955\ : std_logic;
signal \N__27952\ : std_logic;
signal \N__27949\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27910\ : std_logic;
signal \N__27907\ : std_logic;
signal \N__27904\ : std_logic;
signal \N__27903\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27865\ : std_logic;
signal \N__27862\ : std_logic;
signal \N__27859\ : std_logic;
signal \N__27856\ : std_logic;
signal \N__27853\ : std_logic;
signal \N__27850\ : std_logic;
signal \N__27849\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27820\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27759\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27692\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27671\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27663\ : std_logic;
signal \N__27660\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27657\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27617\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27575\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27502\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27460\ : std_logic;
signal \N__27457\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27452\ : std_logic;
signal \N__27451\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27335\ : std_logic;
signal \N__27332\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27292\ : std_logic;
signal \N__27289\ : std_logic;
signal \N__27286\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27123\ : std_logic;
signal \N__27120\ : std_logic;
signal \N__27117\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27109\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27105\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27100\ : std_logic;
signal \N__27097\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27092\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27078\ : std_logic;
signal \N__27075\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27054\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27034\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26943\ : std_logic;
signal \N__26942\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26876\ : std_logic;
signal \N__26873\ : std_logic;
signal \N__26870\ : std_logic;
signal \N__26867\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26848\ : std_logic;
signal \N__26845\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26834\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26830\ : std_logic;
signal \N__26827\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26801\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26791\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26517\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26436\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26347\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26341\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26305\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26206\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26103\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25885\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25758\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25708\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25525\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25511\ : std_logic;
signal \N__25508\ : std_logic;
signal \N__25505\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25462\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25390\ : std_logic;
signal \N__25387\ : std_logic;
signal \N__25384\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25375\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25305\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25285\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25251\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25231\ : std_logic;
signal \N__25228\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25219\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25192\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25069\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25003\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24994\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24988\ : std_logic;
signal \N__24985\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24845\ : std_logic;
signal \N__24842\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24826\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24778\ : std_logic;
signal \N__24775\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24735\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24717\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24682\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24643\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24640\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24587\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24400\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24395\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24389\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24371\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24290\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24233\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23900\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23835\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23453\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22867\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22701\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22207\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21669\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21442\ : std_logic;
signal \N__21439\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21372\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20919\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20750\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20556\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20212\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20081\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20039\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19861\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19273\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19145\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18907\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18514\ : std_logic;
signal \N__18511\ : std_logic;
signal \N__18508\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18329\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17867\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17553\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15238\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15208\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14857\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \b2v_inst16.count_rst_0_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst16.count_4_11\ : std_logic;
signal \b2v_inst16.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst16.count_4_8\ : std_logic;
signal \b2v_inst16.count_rst_8_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst16.count_4_3\ : std_logic;
signal \b2v_inst16.countZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst16.count_rst_14\ : std_logic;
signal \b2v_inst16.count_4_9\ : std_logic;
signal \b2v_inst16.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst16.count_4_7\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_1\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_2\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_5\ : std_logic;
signal \b2v_inst16.countZ0Z_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_6\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8\ : std_logic;
signal \b2v_inst16.countZ0Z_9\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_8_THRU_CO\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_9\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_10\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_11\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_12\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_13\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_14\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgd_en\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgdZ0\ : std_logic;
signal \b2v_inst16.delayed_vddq_pwrgd_en_cascade_\ : std_logic;
signal b2v_inst16_un2_vpp_en_0_i : std_logic;
signal \b2v_inst200.count_enZ0\ : std_logic;
signal \b2v_inst16.count_rst_7\ : std_logic;
signal \b2v_inst16.count_en_cascade_\ : std_logic;
signal \b2v_inst16.count_4_2\ : std_logic;
signal \b2v_inst11.g3_cascade_\ : std_logic;
signal \b2v_inst11.g1_0_1_cascade_\ : std_logic;
signal \b2v_inst11.N_7_3_0_cascade_\ : std_logic;
signal \b2v_inst11.g2_1_0_0_cascade_\ : std_logic;
signal \b2v_inst11.g2_2_0\ : std_logic;
signal \b2v_inst11.g2_1_0\ : std_logic;
signal \b2v_inst11.g0_12_0\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\ : std_logic;
signal \b2v_inst11.N_379_cascade_\ : std_logic;
signal \SLP_S3n_ibuf_RNIF6NLZ0\ : std_logic;
signal \b2v_inst11.N_379\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2\ : std_logic;
signal \b2v_inst11.count_clk_RNIVS8U1Z0Z_14\ : std_logic;
signal \b2v_inst11.N_428\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_0\ : std_logic;
signal \b2v_inst11.N_175\ : std_logic;
signal \b2v_inst11.N_175_cascade_\ : std_logic;
signal \b2v_inst11.N_190\ : std_logic;
signal \b2v_inst11.N_190_cascade_\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o3_0_4\ : std_logic;
signal \b2v_inst11.count_clk_en_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_13\ : std_logic;
signal \b2v_inst11.count_clk_0_15\ : std_logic;
signal \b2v_inst11.count_clk_0_12\ : std_logic;
signal \b2v_inst11.count_clk_0_10\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_o2_4\ : std_logic;
signal \b2v_inst11.count_clk_0_11\ : std_logic;
signal \b2v_inst11.count_clk_0_4\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_1\ : std_logic;
signal \b2v_inst20.counter_1_cry_2\ : std_logic;
signal \b2v_inst20.counter_1_cry_3\ : std_logic;
signal \b2v_inst20.counter_1_cry_4\ : std_logic;
signal \b2v_inst20.counter_1_cry_5\ : std_logic;
signal \b2v_inst20.counter_1_cry_6\ : std_logic;
signal \b2v_inst20.counter_1_cry_7\ : std_logic;
signal \b2v_inst20.counter_1_cry_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_9\ : std_logic;
signal \b2v_inst20.counter_1_cry_10\ : std_logic;
signal \b2v_inst20.counter_1_cry_11\ : std_logic;
signal \b2v_inst20.counter_1_cry_12\ : std_logic;
signal \b2v_inst20.counter_1_cry_13\ : std_logic;
signal \b2v_inst20.counter_1_cry_14\ : std_logic;
signal \b2v_inst20.counter_1_cry_15\ : std_logic;
signal \b2v_inst20.counter_1_cry_16\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_17\ : std_logic;
signal \b2v_inst20.counter_1_cry_18\ : std_logic;
signal \b2v_inst20.counter_1_cry_19\ : std_logic;
signal \b2v_inst20.counter_1_cry_20\ : std_logic;
signal \b2v_inst20.counter_1_cry_21\ : std_logic;
signal \b2v_inst20.counter_1_cry_22\ : std_logic;
signal \b2v_inst20.counter_1_cry_23\ : std_logic;
signal \b2v_inst20.counter_1_cry_24\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \b2v_inst20.counter_1_cry_25\ : std_logic;
signal \b2v_inst20.counter_1_cry_26\ : std_logic;
signal \b2v_inst20.counter_1_cry_27\ : std_logic;
signal \b2v_inst20.counter_1_cry_28\ : std_logic;
signal \b2v_inst20.counter_1_cry_29\ : std_logic;
signal \b2v_inst20.counter_1_cry_30\ : std_logic;
signal \b2v_inst16.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_8\ : std_logic;
signal \b2v_inst16.N_416_cascade_\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst16.count_rst_13\ : std_logic;
signal \b2v_inst16.count_rst_5\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst16.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst16.count_4_5\ : std_logic;
signal \b2v_inst16.countZ0Z_5\ : std_logic;
signal \b2v_inst16.count_rst\ : std_logic;
signal \b2v_inst16.count_4_10\ : std_logic;
signal \b2v_inst16.count_rst_11\ : std_logic;
signal \b2v_inst16.count_4_6\ : std_logic;
signal \b2v_inst16.count_rst_4\ : std_logic;
signal \b2v_inst16.count_4_15\ : std_logic;
signal \b2v_inst16.count_4_14\ : std_logic;
signal \b2v_inst16.count_rst_3\ : std_logic;
signal \b2v_inst16.countZ0Z_14\ : std_logic;
signal \b2v_inst16.countZ0Z_3\ : std_logic;
signal \b2v_inst16.countZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_13\ : std_logic;
signal \b2v_inst16.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_4\ : std_logic;
signal \b2v_inst16.un4_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst16.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst16.count_4_4\ : std_logic;
signal \b2v_inst16.count_rst_2\ : std_logic;
signal \b2v_inst16.count_4_13\ : std_logic;
signal \b2v_inst16.un4_count_1_axb_1_cascade_\ : std_logic;
signal \b2v_inst16.un4_count_1_axb_1\ : std_logic;
signal \b2v_inst16.countZ0Z_6\ : std_logic;
signal \b2v_inst16.countZ0Z_12\ : std_logic;
signal \b2v_inst16.countZ0Z_10\ : std_logic;
signal \b2v_inst16.countZ0Z_2\ : std_logic;
signal \b2v_inst16.count_4_1\ : std_logic;
signal \b2v_inst16.count_rst_6\ : std_logic;
signal \b2v_inst16.countZ0Z_15\ : std_logic;
signal \b2v_inst16.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst16.countZ0Z_11\ : std_logic;
signal \b2v_inst16.count_4_i_a3_8_0\ : std_logic;
signal \b2v_inst16.count_4_i_a3_10_0\ : std_logic;
signal \b2v_inst16.count_4_i_a3_7_0_cascade_\ : std_logic;
signal \b2v_inst16.count_4_i_a3_9_0\ : std_logic;
signal \b2v_inst16.N_414\ : std_logic;
signal \b2v_inst16.countZ0Z_0\ : std_logic;
signal \b2v_inst16.N_414_cascade_\ : std_logic;
signal \b2v_inst16.count_4_0\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_1\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_off_0_1\ : std_logic;
signal \b2v_inst11.count_off_0_0\ : std_logic;
signal \b2v_inst11.count_off_0_10\ : std_logic;
signal \b2v_inst16.N_1440\ : std_logic;
signal \b2v_inst16.curr_state_RNI3B692Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst16.N_416\ : std_logic;
signal \b2v_inst16.curr_state_7_0_1_cascade_\ : std_logic;
signal \b2v_inst16.curr_state_2_1\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst16.curr_state_2_0\ : std_logic;
signal \b2v_inst16.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst16.curr_state_RNI3B692Z0Z_0\ : std_logic;
signal \b2v_inst16.N_268\ : std_logic;
signal \b2v_inst16.N_268_cascade_\ : std_logic;
signal \b2v_inst16.N_26\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_a3_0_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNINPGR_2Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.g0_20_1\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNIVS8U1Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_329_N\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_1_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI_1Z0Z_0\ : std_logic;
signal \N_236_0\ : std_logic;
signal \b2v_inst11.g1_0_0_1\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_331_N\ : std_logic;
signal \b2v_inst11.count_clk_en_1\ : std_logic;
signal \b2v_inst11.N_328\ : std_logic;
signal \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1\ : std_logic;
signal \b2v_inst11.N_340\ : std_logic;
signal \b2v_inst11.func_state_1_ss0_i_0_o3_1\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI_1Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_4_i_a3_0_1\ : std_logic;
signal \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_0_1\ : std_logic;
signal \b2v_inst11.count_clk_0_0\ : std_logic;
signal \b2v_inst11.count_clk_0_7\ : std_logic;
signal \b2v_inst11.N_168_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNICGI84_0_0_cascade_\ : std_logic;
signal \b2v_inst11.count_clk_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst11.func_state_RNIVS8U1_0Z0Z_0\ : std_logic;
signal \b2v_inst11.count_clk_0_14\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_2\ : std_logic;
signal \b2v_inst11.un1_count_clk_1_sqmuxa_0_3\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_1\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_0\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_7\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_6\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_cZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8\ : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_10\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_11\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_10_cZ0\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_12\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_11\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_13\ : std_logic;
signal \b2v_inst11.count_clk_1_13\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_12\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_14\ : std_logic;
signal \b2v_inst11.count_clk_1_14\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_13\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_15\ : std_logic;
signal \b2v_inst11.func_state_RNICGI84_0_0\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_14\ : std_logic;
signal \b2v_inst11.count_clk_1_15\ : std_logic;
signal \b2v_inst20.counterZ0Z_11\ : std_logic;
signal \b2v_inst20.counterZ0Z_9\ : std_logic;
signal \b2v_inst20.counterZ0Z_10\ : std_logic;
signal \b2v_inst20.counterZ0Z_8\ : std_logic;
signal \b2v_inst20.counterZ0Z_15\ : std_logic;
signal \b2v_inst20.counterZ0Z_14\ : std_logic;
signal \b2v_inst20.counterZ0Z_13\ : std_logic;
signal \b2v_inst20.counterZ0Z_12\ : std_logic;
signal \b2v_inst20.counterZ0Z_19\ : std_logic;
signal \b2v_inst20.counterZ0Z_17\ : std_logic;
signal \b2v_inst20.counterZ0Z_18\ : std_logic;
signal \b2v_inst20.counterZ0Z_16\ : std_logic;
signal \b2v_inst20.counterZ0Z_23\ : std_logic;
signal \b2v_inst20.counterZ0Z_21\ : std_logic;
signal \b2v_inst20.counterZ0Z_22\ : std_logic;
signal \b2v_inst20.counterZ0Z_20\ : std_logic;
signal \VPP_OK_c\ : std_logic;
signal \VDDQ_EN_c\ : std_logic;
signal \bfn_2_15_0_\ : std_logic;
signal \b2v_inst20.un4_counter_0\ : std_logic;
signal \b2v_inst20.un4_counter_2_and\ : std_logic;
signal \b2v_inst20.un4_counter_1\ : std_logic;
signal \b2v_inst20.un4_counter_3_and\ : std_logic;
signal \b2v_inst20.un4_counter_2\ : std_logic;
signal \b2v_inst20.un4_counter_4_and\ : std_logic;
signal \b2v_inst20.un4_counter_3\ : std_logic;
signal \b2v_inst20.un4_counter_5_and\ : std_logic;
signal \b2v_inst20.un4_counter_4\ : std_logic;
signal \b2v_inst20.un4_counter_5\ : std_logic;
signal \b2v_inst20.un4_counter_6\ : std_logic;
signal b2v_inst20_un4_counter_7 : std_logic;
signal \bfn_2_16_0_\ : std_logic;
signal \b2v_inst20.counterZ0Z_31\ : std_logic;
signal \b2v_inst20.counterZ0Z_29\ : std_logic;
signal \b2v_inst20.counterZ0Z_30\ : std_logic;
signal \b2v_inst20.counterZ0Z_28\ : std_logic;
signal \b2v_inst20.un4_counter_7_and\ : std_logic;
signal \b2v_inst20.counterZ0Z_27\ : std_logic;
signal \b2v_inst20.counterZ0Z_25\ : std_logic;
signal \b2v_inst20.counterZ0Z_26\ : std_logic;
signal \b2v_inst20.counterZ0Z_24\ : std_logic;
signal \b2v_inst20.un4_counter_6_and\ : std_logic;
signal \b2v_inst200.count_3_1\ : std_logic;
signal \b2v_inst200.count_3_2\ : std_logic;
signal \b2v_inst200.count_3_3\ : std_logic;
signal \b2v_inst200.count_3_12\ : std_logic;
signal \b2v_inst200.count_3_4\ : std_logic;
signal \b2v_inst200.count_3_5\ : std_logic;
signal \b2v_inst200.count_3_7\ : std_logic;
signal \b2v_inst11.count_off_0_15\ : std_logic;
signal \b2v_inst11.count_off_0_13\ : std_logic;
signal \b2v_inst11.count_offZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.count_off_0_8\ : std_logic;
signal \b2v_inst11.count_offZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.count_offZ0Z_0\ : std_logic;
signal \bfn_4_4_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6\ : std_logic;
signal \b2v_inst11.count_offZ0Z_8\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_7\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11\ : std_logic;
signal \b2v_inst11.count_offZ0Z_13\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_12\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13\ : std_logic;
signal \b2v_inst11.count_offZ0Z_15\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_11\ : std_logic;
signal \b2v_inst11.count_off_1_11\ : std_logic;
signal \b2v_inst11.count_off_1_11_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\ : std_logic;
signal \b2v_inst11.count_off_0_12\ : std_logic;
signal \b2v_inst11.count_offZ0Z_12\ : std_logic;
signal \b2v_inst11.count_offZ0Z_10\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_5\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_4_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_11\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_11\ : std_logic;
signal \b2v_inst11.g4_cascade_\ : std_logic;
signal \b2v_inst11.g0_17_N_3L3_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIVGS13Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNI24DD8Z0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_RNIVGS13Z0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.N_160_i_cascade_\ : std_logic;
signal \b2v_inst11.g1_0_sx\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI608H1_0Z0Z_1\ : std_logic;
signal \b2v_inst11.N_354_cascade_\ : std_logic;
signal b2v_inst11_g0_i_m2_i_a6_3_2 : std_logic;
signal \b2v_inst11.N_159_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m0_0_1_1_0_cascade_\ : std_logic;
signal \b2v_inst11.un1_func_state25_6_0_o_N_313_N\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_sx_cascade_\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1\ : std_logic;
signal \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.N_337\ : std_logic;
signal \b2v_inst11.func_state_1_m2s2_i_0_cascade_\ : std_logic;
signal \b2v_inst11.N_338\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.N_231_N\ : std_logic;
signal \b2v_inst11.N_306_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI_1Z0Z_1\ : std_logic;
signal \b2v_inst11.func_state_1_m2_am_1_1_cascade_\ : std_logic;
signal \b2v_inst11.count_off_RNIZ0Z_9\ : std_logic;
signal \b2v_inst11.func_state_RNIR5S85Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.func_state_cascade_\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.N_160_i\ : std_logic;
signal \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\ : std_logic;
signal \b2v_inst11.func_state_1_m0_0_1_0\ : std_logic;
signal \b2v_inst11.func_state_1_m2_1_0_cascade_\ : std_logic;
signal \b2v_inst11.N_76\ : std_logic;
signal \b2v_inst11.func_state_1_m2_0\ : std_logic;
signal \func_state_RNIVS8U1_4_1\ : std_logic;
signal \b2v_inst11.func_stateZ0Z_1\ : std_logic;
signal \b2v_inst11.count_clk_enZ0Z_0\ : std_logic;
signal \VCCST_EN_i_0_o3_0_cascade_\ : std_logic;
signal \b2v_inst11.func_state_1_m2_1\ : std_logic;
signal \func_state_RNI6BE8E_0_1_cascade_\ : std_logic;
signal \b2v_inst11.count_0_7\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_3\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_6\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_8\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_2\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_9\ : std_logic;
signal \b2v_inst11.count_clkZ0Z_9\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_3\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_5\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_6\ : std_logic;
signal \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\ : std_logic;
signal \b2v_inst11.count_clk_0_8\ : std_logic;
signal \b2v_inst11.count_clk_en\ : std_logic;
signal \b2v_inst20.un4_counter_0_and\ : std_logic;
signal \b2v_inst11.N_381_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_\ : std_logic;
signal \b2v_inst11.N_381_0\ : std_logic;
signal \N_15_i_0_a4_0_1\ : std_logic;
signal \b2v_inst20.counter_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_3\ : std_logic;
signal \b2v_inst20.counterZ0Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\ : std_logic;
signal \b2v_inst20.counter_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_4\ : std_logic;
signal \b2v_inst20.counter_1_cry_4_THRU_CO\ : std_logic;
signal \delayed_vccin_vccinaux_ok_RNI8L1J7_0\ : std_logic;
signal \b2v_inst20.counter_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_2\ : std_logic;
signal \bfn_5_1_0_\ : std_logic;
signal \b2v_inst200.countZ0Z_1\ : std_logic;
signal \b2v_inst200.count_RNIC03N_5Z0Z_0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1_cy\ : std_logic;
signal \b2v_inst200.countZ0Z_2\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst200.countZ0Z_3\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst200.countZ0Z_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_5_cZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_7\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_15\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16\ : std_logic;
signal \b2v_inst200.count_0_17\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\ : std_logic;
signal \b2v_inst11.count_off_1_3_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_3\ : std_logic;
signal \b2v_inst11.count_offZ0Z_4\ : std_logic;
signal \b2v_inst11.count_off_1_3\ : std_logic;
signal \b2v_inst11.count_offZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\ : std_logic;
signal \b2v_inst11.count_offZ0Z_3\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\ : std_logic;
signal \b2v_inst11.count_off_0_4\ : std_logic;
signal \b2v_inst11.count_off_0_14\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_14\ : std_logic;
signal \b2v_inst11.count_off_1_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_2\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\ : std_logic;
signal \b2v_inst11.count_offZ0Z_2\ : std_logic;
signal \b2v_inst11.count_offZ0Z_5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_1\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_0\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_2\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_1_cascade_\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_3\ : std_logic;
signal \b2v_inst11.un34_clk_100khz_12\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\ : std_logic;
signal \b2v_inst11.count_off_0_5\ : std_logic;
signal \b2v_inst11.count_offZ0Z_6\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\ : std_logic;
signal \b2v_inst11.count_off_1_9\ : std_logic;
signal \b2v_inst11.count_offZ0Z_9\ : std_logic;
signal \b2v_inst11.count_off_1_9_cascade_\ : std_logic;
signal \b2v_inst11.un3_count_off_1_axb_9\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\ : std_logic;
signal \b2v_inst11.count_off_1_6\ : std_logic;
signal \b2v_inst11.count_offZ0Z_7\ : std_logic;
signal \b2v_inst11.count_off_enZ0\ : std_logic;
signal \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\ : std_logic;
signal \b2v_inst11.N_125\ : std_logic;
signal \b2v_inst11.count_off_1_7\ : std_logic;
signal \b2v_inst11.g0_3_0\ : std_logic;
signal \b2v_inst11.g2_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena_8_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_rst_7\ : std_logic;
signal \b2v_inst11.dutycycle_0_3\ : std_logic;
signal \b2v_inst11.dutycycle_rst_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_eena_8\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_0_ccf1\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_43_and_i_0_c\ : std_logic;
signal \b2v_inst11.N_307_cascade_\ : std_logic;
signal \b2v_inst11.N_234_N\ : std_logic;
signal \b2v_inst11.N_308\ : std_logic;
signal \b2v_inst11.N_234_N_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI9R6T4Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.func_state_RNI9R6T4Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_11\ : std_logic;
signal \b2v_inst11.N_159\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\ : std_logic;
signal \b2v_inst11.N_155_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_en_11_cascade_\ : std_logic;
signal \b2v_inst11.N_305\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_6\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst11.i2_mux_cascade_\ : std_logic;
signal \b2v_inst11.N_301\ : std_logic;
signal \b2v_inst11.N_382_cascade_\ : std_logic;
signal \b2v_inst11.g0_2_0_cascade_\ : std_logic;
signal \b2v_inst11.N_430\ : std_logic;
signal \b2v_inst11.func_state_RNIRF2E4Z0Z_0\ : std_logic;
signal \VCCST_EN_i_0_i\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_2_i_o3_sx\ : std_logic;
signal \b2v_inst11.func_state\ : std_logic;
signal \b2v_inst11.func_state_RNI_0Z0Z_0\ : std_logic;
signal \b2v_inst5.N_2897_i_cascade_\ : std_logic;
signal \b2v_inst5.curr_state_0_0\ : std_logic;
signal \b2v_inst5.m4_0_cascade_\ : std_logic;
signal \b2v_inst11.g2_0_1_cascade_\ : std_logic;
signal \dutycycle_RNISSAOS1_0_5_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_1\ : std_logic;
signal \b2v_inst11.N_73_mux_i_i_o7_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIUNGA5Z0Z_5\ : std_logic;
signal \b2v_inst11.N_73_mux_i_i_0\ : std_logic;
signal \b2v_inst11.N_73_mux_i_i_a7_1_cascade_\ : std_logic;
signal g0_0_0 : std_logic;
signal \N_5_0\ : std_logic;
signal b2v_inst11_un1_dutycycle_172_m3_amcf1 : std_logic;
signal \N_73_mux_i_i_a7_4_0_1_cascade_\ : std_logic;
signal \N_73_mux_i_i_a7_4_0_cascade_\ : std_logic;
signal \b2v_inst11.N_73_mux_i_i_1\ : std_logic;
signal \b2v_inst11.N_73_mux_i_i_2\ : std_logic;
signal \N_15\ : std_logic;
signal \b2v_inst11.N_73_mux_i_i_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_0_5\ : std_logic;
signal \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx\ : std_logic;
signal \RSMRSTn_fast_RNIGMH81_cascade_\ : std_logic;
signal \N_7_2\ : std_logic;
signal \N_10_0\ : std_logic;
signal \b2v_inst20.tmp_1_rep1_RNI07FZ0Z73\ : std_logic;
signal \b2v_inst20.counter_1_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst20.counterZ0Z_7\ : std_logic;
signal \b2v_inst20.counterZ0Z_5\ : std_logic;
signal \b2v_inst20.counterZ0Z_6\ : std_logic;
signal \b2v_inst20.counterZ0Z_1\ : std_logic;
signal \b2v_inst20.un4_counter_1_and\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3_fast\ : std_logic;
signal \HDA_SDO_ATP_c\ : std_logic;
signal \b2v_inst200.N_205\ : std_logic;
signal \b2v_inst200.N_205_cascade_\ : std_logic;
signal \G_2734_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_2\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst200.HDA_SDO_ATP_0\ : std_logic;
signal \G_2734\ : std_logic;
signal \b2v_inst200.curr_state_0_2\ : std_logic;
signal \b2v_inst200.countZ0Z_6\ : std_logic;
signal \b2v_inst200.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_8\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\ : std_logic;
signal \b2v_inst200.count_3_6\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0\ : std_logic;
signal \b2v_inst200.count_3_8\ : std_logic;
signal \b2v_inst200.count_1_0\ : std_logic;
signal \b2v_inst200.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst200.count_3_0\ : std_logic;
signal \b2v_inst200.countZ0Z_12\ : std_logic;
signal \b2v_inst200.count_3_13\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\ : std_logic;
signal \b2v_inst200.countZ0Z_13\ : std_logic;
signal \b2v_inst200.countZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_0\ : std_logic;
signal \b2v_inst200.countZ0Z_7\ : std_logic;
signal \b2v_inst200.countZ0Z_5\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_10_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_3\ : std_logic;
signal \b2v_inst200.countZ0Z_15\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\ : std_logic;
signal \b2v_inst200.count_3_15\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\ : std_logic;
signal \b2v_inst200.count_3_14\ : std_logic;
signal \b2v_inst200.countZ0Z_14\ : std_logic;
signal \b2v_inst200.count_0_16\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29\ : std_logic;
signal \b2v_inst200.count_3_11\ : std_logic;
signal \b2v_inst200.countZ0Z_11\ : std_logic;
signal \b2v_inst200.countZ0Z_17\ : std_logic;
signal \b2v_inst200.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_16\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_9\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_12\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_13_cascade_\ : std_logic;
signal \b2v_inst200.un25_clk_100khz_14\ : std_logic;
signal \b2v_inst200.count_RNIC03N_6Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0\ : std_logic;
signal \b2v_inst200.count_3_10\ : std_logic;
signal \b2v_inst200.count_RNI_0_0_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_10\ : std_logic;
signal \b2v_inst16.count_rst_1\ : std_logic;
signal \b2v_inst16.count_4_12\ : std_logic;
signal \b2v_inst16.count_en\ : std_logic;
signal \b2v_inst16.N_2987_i\ : std_logic;
signal \b2v_inst11.N_366\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_2_c\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3_c\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4_c\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5_c\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6_c\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i_0_8\ : std_logic;
signal \VDDQ_OK_c\ : std_logic;
signal \VCCST_EN_i_0_o3_0\ : std_logic;
signal \b2v_inst16.N_208_0\ : std_logic;
signal \b2v_inst11.N_354\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_a2_1_3\ : std_logic;
signal \b2v_inst11.un2_count_clk_17_0_a2_1_2_cascade_\ : std_logic;
signal \b2v_inst11.N_363\ : std_logic;
signal \b2v_inst11.N_360\ : std_logic;
signal \b2v_inst11.N_363_cascade_\ : std_logic;
signal \b2v_inst11.N_365\ : std_logic;
signal \b2v_inst11.N_365_cascade_\ : std_logic;
signal \b2v_inst11.N_293\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_30_1_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_7Z0Z_1\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_2\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_4_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_10_cZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\ : std_logic;
signal \b2v_inst11.dutycycle_RNIP7P13Z0Z_4\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNIP7P13Z0Z_4_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_4\ : std_logic;
signal \b2v_inst11.N_158_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_0_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQZ0Z6\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_6\ : std_logic;
signal \b2v_inst11.func_state_RNI_5Z0Z_1\ : std_logic;
signal \b2v_inst11.N_186_cascade_\ : std_logic;
signal \b2v_inst11.N_426_0\ : std_logic;
signal \b2v_inst11_g0_i_m2_i_a6_1_1_cascade_\ : std_logic;
signal \SLP_S3n_ibuf_RNI9HQHZ0Z3\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_9Z0Z_1\ : std_logic;
signal \b2v_inst11.N_165_0\ : std_logic;
signal \b2v_inst11.g0_i_m2_i_0_1_cascade_\ : std_logic;
signal \N_15_i_0_a4_1_0\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_0\ : std_logic;
signal \b2v_inst11.N_19_i\ : std_logic;
signal \b2v_inst11.N_5572_0\ : std_logic;
signal \b2v_inst11.N_172\ : std_logic;
signal \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_0\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_0\ : std_logic;
signal \b2v_inst11.dutycycle_eena_cascade_\ : std_logic;
signal \b2v_inst11.N_117_f0_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena_0_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_1\ : std_logic;
signal \b2v_inst11.dutycycle_eena_0\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_1\ : std_logic;
signal \b2v_inst5.curr_state_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst5_RSMRSTn_latmux\ : std_logic;
signal \b2v_inst5_RSMRSTn_fast\ : std_logic;
signal \RSMRSTn_0\ : std_logic;
signal \b2v_inst5.N_2897_i\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst5.curr_state_RNIZ0Z_1\ : std_logic;
signal \b2v_inst5.N_51_cascade_\ : std_logic;
signal \b2v_inst11.count_0_9\ : std_logic;
signal \b2v_inst11.count_0_10\ : std_logic;
signal \b2v_inst11.count_0_11\ : std_logic;
signal \b2v_inst11.count_0_2\ : std_logic;
signal \b2v_inst200.N_56_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst200.count_RNI_0_0\ : std_logic;
signal \GPIO_FPGA_SoC_1_c\ : std_logic;
signal \N_411_cascade_\ : std_logic;
signal \b2v_inst200.m6_i_0\ : std_logic;
signal \b2v_inst200.m6_i_0_cascade_\ : std_logic;
signal \b2v_inst200.curr_state_3_0\ : std_logic;
signal \b2v_inst200.N_58_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \N_412\ : std_logic;
signal \N_412_cascade_\ : std_logic;
signal \b2v_inst200.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst200.curr_state_3_1\ : std_logic;
signal \b2v_inst36.count_2_6\ : std_logic;
signal \b2v_inst36.count_2_4\ : std_logic;
signal \b2v_inst36.count_2_9\ : std_logic;
signal \b2v_inst36.count_2_12\ : std_logic;
signal \b2v_inst36.curr_state_RNI8TT2Z0Z_0_cascade_\ : std_logic;
signal \DSW_PWROK_c\ : std_logic;
signal \b2v_inst36.DSW_PWROK_0\ : std_logic;
signal \b2v_inst36.curr_state_0_0\ : std_logic;
signal \b2v_inst36.curr_state_7_0_cascade_\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.N_2939_i_cascade_\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_7_l_fx\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i_0_8\ : std_logic;
signal \b2v_inst11.N_382\ : std_logic;
signal \b2v_inst11.N_302\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_9\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_axb_4_l_fx\ : std_logic;
signal \b2v_inst11.g0_13_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_9_cascade_\ : std_logic;
signal \b2v_inst200.count_RNIC03N_6Z0Z_0\ : std_logic;
signal \N_411\ : std_logic;
signal \b2v_inst200.m11_0_a3_0\ : std_logic;
signal \b2v_inst5.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_4_cascade_\ : std_logic;
signal \b2v_inst5.count_1_8\ : std_logic;
signal \b2v_inst5.count_rst_10\ : std_logic;
signal \b2v_inst5.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst5.count_1_4\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_7_cascade_\ : std_logic;
signal \b2v_inst11.N_8_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\ : std_logic;
signal \b2v_inst11.dutycycle_en_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_14\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_3\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.N_153_N_cascade_\ : std_logic;
signal \b2v_inst11.N_156_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_9_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\ : std_logic;
signal \b2v_inst11.dutycycle_en_10\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_13\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst11.N_326_N\ : std_logic;
signal \b2v_inst11.N_140_N\ : std_logic;
signal \b2v_inst11.N_425\ : std_logic;
signal \b2v_inst11.N_154_N_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_en_4_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_e_1_8\ : std_logic;
signal \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\ : std_logic;
signal \b2v_inst11.dutycycle_en_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_10\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_8\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49\ : std_logic;
signal \b2v_inst11.dutycycle_RNI1KT13Z0Z_8\ : std_logic;
signal \GPIO_FPGA_SoC_4_c\ : std_logic;
signal \N_161\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\ : std_logic;
signal \SLP_S3n_c\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIZ0\ : std_logic;
signal \b2v_inst11.func_state_RNI_2Z0Z_1\ : std_logic;
signal \SLP_S4n_c\ : std_logic;
signal \b2v_inst11.g1_0_0_cascade_\ : std_logic;
signal \b2v_inst11.N_295\ : std_logic;
signal \b2v_inst11.g1\ : std_logic;
signal \b2v_inst11.g1_cascade_\ : std_logic;
signal \b2v_inst11.g1_0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_2\ : std_logic;
signal \RSMRSTn_fast_RNIGMH81\ : std_logic;
signal \func_state_RNI6BE8E_0_1\ : std_logic;
signal b2v_inst11_dutycycle_1_0_iv_0_o3_out : std_logic;
signal \func_state_RNI_4_0\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \b2v_inst11.count_1_2\ : std_logic;
signal \b2v_inst11.un1_count_cry_1\ : std_logic;
signal \b2v_inst11.un1_count_cry_2\ : std_logic;
signal \b2v_inst11.un1_count_cry_3\ : std_logic;
signal \b2v_inst11.un1_count_cry_4\ : std_logic;
signal \b2v_inst11.un1_count_cry_5\ : std_logic;
signal \b2v_inst11.count_1_7\ : std_logic;
signal \b2v_inst11.un1_count_cry_6\ : std_logic;
signal \b2v_inst11.un1_count_cry_7\ : std_logic;
signal \b2v_inst11.un1_count_cry_8\ : std_logic;
signal \b2v_inst11.count_1_9\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \b2v_inst11.count_1_10\ : std_logic;
signal \b2v_inst11.un1_count_cry_9\ : std_logic;
signal \b2v_inst11.count_1_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_10\ : std_logic;
signal \b2v_inst11.un1_count_cry_11\ : std_logic;
signal \b2v_inst11.un1_count_cry_12\ : std_logic;
signal \b2v_inst11.un1_count_cry_13\ : std_logic;
signal \b2v_inst11.un1_count_cry_14\ : std_logic;
signal \b2v_inst11.count_1_5\ : std_logic;
signal \b2v_inst11.count_0_5\ : std_logic;
signal \b2v_inst11.count_1_14\ : std_logic;
signal \b2v_inst11.count_0_14\ : std_logic;
signal \b2v_inst11.count_1_6\ : std_logic;
signal \b2v_inst11.count_0_6\ : std_logic;
signal \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\ : std_logic;
signal \b2v_inst11.count_0_15\ : std_logic;
signal \b2v_inst11.pwm_out_en_cascade_\ : std_logic;
signal \PWRBTN_LED_c\ : std_logic;
signal \b2v_inst11.pwm_out_1_sqmuxa_0\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3_rep1\ : std_logic;
signal \b2v_inst20_un4_counter_7_THRU_CO\ : std_logic;
signal \b2v_inst36.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_9\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_10_cascade_\ : std_logic;
signal \b2v_inst36.count_2_0\ : std_logic;
signal \b2v_inst36.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst36.count_rst_13\ : std_logic;
signal \b2v_inst36.count_rst_13_cascade_\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_1_cascade_\ : std_logic;
signal \b2v_inst36.count_2_1\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_8\ : std_logic;
signal \b2v_inst36.count_rst_14\ : std_logic;
signal \b2v_inst36.count_rst_3_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst36.count_2_11\ : std_logic;
signal \b2v_inst36.count_rst_12_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_2_cascade_\ : std_logic;
signal \b2v_inst36.count_2_2\ : std_logic;
signal \b2v_inst36.curr_state_7_1\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst36.curr_state_0_1\ : std_logic;
signal \b2v_inst36.N_2939_i\ : std_logic;
signal \V33DSW_OK_c\ : std_logic;
signal \b2v_inst36.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst36.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst36.N_2942_i_cascade_\ : std_logic;
signal \b2v_inst200.countZ0Z_9\ : std_logic;
signal \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\ : std_logic;
signal \b2v_inst200.count_3_9\ : std_logic;
signal \b2v_inst200.count_en_g\ : std_logic;
signal \b2v_inst36.count_2_14\ : std_logic;
signal \b2v_inst5.count_1_11\ : std_logic;
signal \b2v_inst5.count_1_12\ : std_logic;
signal \b2v_inst5.count_1_14\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i_0_8\ : std_logic;
signal \b2v_inst5.curr_stateZ0Z_1\ : std_logic;
signal \N_413\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_11\ : std_logic;
signal \b2v_inst11.i7_mux_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_11_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_3Z0Z_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_8_cascade_\ : std_logic;
signal \b2v_inst11.N_15_mux\ : std_logic;
signal \b2v_inst11.i6_mux_i_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_11\ : std_logic;
signal \b2v_inst11.dutycycle_RNI9R6T4Z0Z_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_12\ : std_logic;
signal \b2v_inst11.N_224_iZ0\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_15\ : std_logic;
signal \func_state_RNIVS8U1_3_1\ : std_logic;
signal \b2v_inst11.dutycycle_en_12\ : std_logic;
signal \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_3_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_1_i_i_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_1\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_1_i_0_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_3_cascade_\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_5\ : std_logic;
signal \b2v_inst11.m6_0_1\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_0_1\ : std_logic;
signal \N_18\ : std_logic;
signal \b2v_inst11.g2_0_0\ : std_logic;
signal b2v_inst11_un1_dutycycle_164_0 : std_logic;
signal \b2v_inst5.N_6\ : std_logic;
signal \b2v_inst11_un1_dutycycle_164_0_cascade_\ : std_logic;
signal \b2v_inst5.N_13\ : std_logic;
signal \b2v_inst11.N_3060_i\ : std_logic;
signal \b2v_inst11.un1_dutycycle_96_0_a3_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_7\ : std_logic;
signal \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_5\ : std_logic;
signal \N_73_mux_i_i_o3_1_1\ : std_logic;
signal \b2v_inst11.dutycycleZ1Z_3\ : std_logic;
signal \b2v_inst11.g3_0_1\ : std_logic;
signal \b2v_inst11.N_3038_i\ : std_logic;
signal g3_0_4 : std_logic;
signal \b2v_inst11.count_1_12\ : std_logic;
signal \b2v_inst11.count_0_12\ : std_logic;
signal \b2v_inst11.count_1_3\ : std_logic;
signal \b2v_inst11.count_0_3\ : std_logic;
signal \b2v_inst11.count_1_13\ : std_logic;
signal \b2v_inst11.count_0_13\ : std_logic;
signal \b2v_inst11.count_1_4\ : std_logic;
signal \b2v_inst11.count_0_4\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlt6\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_4_cascade_\ : std_logic;
signal \b2v_inst11.un79_clk_100khzlto15_7\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_13_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_1_1_cascade_\ : std_logic;
signal \b2v_inst11.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst11.count_0_1\ : std_logic;
signal \b2v_inst11.count_0_0\ : std_logic;
signal b2v_inst11_dutycycle_set_1 : std_logic;
signal \G_146\ : std_logic;
signal \N_15_i_0_a4_1\ : std_logic;
signal \N_73_mux_i_i_a7_0_0\ : std_logic;
signal \b2v_inst11.count_1_8\ : std_logic;
signal \b2v_inst11.count_0_8\ : std_logic;
signal \b2v_inst11.g0_2_1\ : std_logic;
signal \b2v_inst11.pwm_outZ0\ : std_logic;
signal \b2v_inst11.pwm_out_1_sqmuxa\ : std_logic;
signal \b2v_inst11.curr_state_3_0_cascade_\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i\ : std_logic;
signal \b2v_inst11.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \b2v_inst11.count_1_0\ : std_logic;
signal \b2v_inst36.un2_count_1_axb_1\ : std_logic;
signal \b2v_inst36.countZ0Z_0\ : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst36.countZ0Z_4\ : std_logic;
signal \b2v_inst36.count_rst_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst36.countZ0Z_6\ : std_logic;
signal \b2v_inst36.count_rst_8\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_8\ : std_logic;
signal \b2v_inst36.countZ0Z_9\ : std_logic;
signal \b2v_inst36.count_rst_5\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst36.countZ0Z_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst36.countZ0Z_12\ : std_logic;
signal \b2v_inst36.count_rst_2\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst36.countZ0Z_14\ : std_logic;
signal \b2v_inst36.count_rst_0\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst36.count_rst_6\ : std_logic;
signal \b2v_inst36.countZ0Z_8\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst36.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst36.count_2_8\ : std_logic;
signal \b2v_inst36.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_10\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst36.countZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst36.count_2_10\ : std_logic;
signal \b2v_inst36.countZ0Z_13\ : std_logic;
signal \b2v_inst36.count_rst_1\ : std_logic;
signal \b2v_inst36.count_2_13\ : std_logic;
signal \b2v_inst36.count_2_15\ : std_logic;
signal \b2v_inst36.count_rst\ : std_logic;
signal \b2v_inst36.countZ0Z_15\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_4\ : std_logic;
signal \b2v_inst5.count_1_2\ : std_logic;
signal \b2v_inst5.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst5.count_1_3\ : std_logic;
signal \b2v_inst5.count_RNIZ0Z_1\ : std_logic;
signal \b2v_inst5.count_1_1\ : std_logic;
signal \b2v_inst5.count_rst_14_cascade_\ : std_logic;
signal \b2v_inst5.count_rst_1_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_13_cascade_\ : std_logic;
signal \b2v_inst5.count_rst_1\ : std_logic;
signal \b2v_inst5.count_1_13\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_5\ : std_logic;
signal \b2v_inst5.count_rst_6\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_8\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i_0_8\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i_0_8\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_3\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_axb_0\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_5Z0Z_1\ : std_logic;
signal \b2v_inst11.mult1_un138_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_0\ : std_logic;
signal \b2v_inst11.mult1_un131_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_1\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_2\ : std_logic;
signal \b2v_inst11.mult1_un124_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_2\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_4Z0Z_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_3\ : std_logic;
signal \b2v_inst11.mult1_un117_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_3\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_4\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_9\ : std_logic;
signal \b2v_inst11.mult1_un103_sum\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_9\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_4\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_6\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_7\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_6\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_11\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_12\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_9\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_9\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_0Z0Z_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_10\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_11\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_11\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_8\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_2Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_12\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_12\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_13\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_15\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15\ : std_logic;
signal \b2v_inst11.dutycycle_RNIZ0Z_14\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_11\ : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \b2v_inst11.CO2\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_7\ : std_logic;
signal \dutycycle_RNISSAOS1_0_5\ : std_logic;
signal \b2v_inst11.dutycycle_RNI_1Z0Z_1\ : std_logic;
signal \b2v_inst11.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst11.count_RNIZ0Z_13\ : std_logic;
signal \b2v_inst11.curr_state_4_0\ : std_logic;
signal \b2v_inst11.CO2_THRU_CO\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_s_6\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_l_fx_6\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_5\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_l_fx_3\ : std_logic;
signal \b2v_inst11.mult1_un47_sum\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_s_4_sf\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\ : std_logic;
signal \b2v_inst11.un1_dutycycle_53_i_29\ : std_logic;
signal \dutycycle_RNIU8G3G_0_2\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_axb_7\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_i_0_8\ : std_logic;
signal \b2v_inst5.N_51\ : std_logic;
signal \b2v_inst5.curr_state_0_1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \b2v_inst36.countZ0Z_2\ : std_logic;
signal \b2v_inst36.un12_clk_100khz_11\ : std_logic;
signal \b2v_inst36.count_rst_11_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_3\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst36.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst36.count_2_3\ : std_logic;
signal \b2v_inst36.count_rst_9_cascade_\ : std_logic;
signal \b2v_inst36.countZ0Z_5\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst36.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst36.count_2_5\ : std_logic;
signal \b2v_inst36.countZ0Z_7\ : std_logic;
signal \b2v_inst36.N_2942_i\ : std_logic;
signal \b2v_inst36.N_1_i\ : std_logic;
signal \b2v_inst36.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst36.count_2_7\ : std_logic;
signal \b2v_inst36.count_en\ : std_logic;
signal \b2v_inst36.count_0_sqmuxa\ : std_logic;
signal \b2v_inst6.count_0_14\ : std_logic;
signal \b2v_inst6.countZ0Z_14_cascade_\ : std_logic;
signal \b2v_inst6.count_0_6\ : std_logic;
signal \b2v_inst5.countZ0Z_1\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_2\ : std_logic;
signal \b2v_inst5.count_rst_12\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst5.countZ0Z_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_4\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst5.countZ0Z_8\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst5.count_rst_3\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst5.countZ0Z_12\ : std_logic;
signal \b2v_inst5.count_rst_2\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_13\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst5.countZ0Z_14\ : std_logic;
signal \b2v_inst5.count_rst_0\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst5.countZ0Z_15\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst5.count_rst\ : std_logic;
signal \b2v_inst5.count_1_15\ : std_logic;
signal \b2v_inst5.count_rst_5_cascade_\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_9\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_9_cascade_\ : std_logic;
signal \b2v_inst5.count_1_9\ : std_logic;
signal \b2v_inst5.count_rst_5\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_6\ : std_logic;
signal \b2v_inst5.count_rst_4_cascade_\ : std_logic;
signal \b2v_inst5.countZ0Z_10\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_9_THRU_CO\ : std_logic;
signal \b2v_inst5.countZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst5.count_1_10\ : std_logic;
signal \b2v_inst5.un2_count_1_cry_0\ : std_logic;
signal \b2v_inst5.N_1_i\ : std_logic;
signal \b2v_inst5.count_1_0\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_5\ : std_logic;
signal \b2v_inst5.count_1_6\ : std_logic;
signal \b2v_inst5.count_rst_8\ : std_logic;
signal \b2v_inst5.countZ0Z_6\ : std_logic;
signal \b2v_inst5.count_rst_9\ : std_logic;
signal \b2v_inst5.countZ0Z_6_cascade_\ : std_logic;
signal \b2v_inst5.count_1_5\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_3\ : std_logic;
signal \b2v_inst5.un2_count_1_axb_7\ : std_logic;
signal \b2v_inst5.count_0_sqmuxa\ : std_logic;
signal \b2v_inst5.count_1_7\ : std_logic;
signal \b2v_inst5.count_rst_7\ : std_logic;
signal \b2v_inst5.countZ0Z_11\ : std_logic;
signal \b2v_inst5.curr_state_RNIFLPH1Z0Z_1\ : std_logic;
signal \b2v_inst5.un12_clk_100khz_2\ : std_logic;
signal \b2v_inst11.mult1_un152_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_s_8\ : std_logic;
signal \b2v_inst11.countZ0Z_0\ : std_logic;
signal \b2v_inst11.un1_count_cry_0_i\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \b2v_inst11.countZ0Z_1\ : std_logic;
signal \b2v_inst11.N_5530_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_0\ : std_logic;
signal \b2v_inst11.countZ0Z_2\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_2\ : std_logic;
signal \b2v_inst11.N_5531_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_1\ : std_logic;
signal \b2v_inst11.countZ0Z_3\ : std_logic;
signal \b2v_inst11.mult1_un145_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5532_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_2\ : std_logic;
signal \b2v_inst11.countZ0Z_4\ : std_logic;
signal \b2v_inst11.mult1_un138_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5533_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_3\ : std_logic;
signal \b2v_inst11.countZ0Z_5\ : std_logic;
signal \b2v_inst11.mult1_un131_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5534_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un124_sum_i_8\ : std_logic;
signal \b2v_inst11.countZ0Z_6\ : std_logic;
signal \b2v_inst11.N_5535_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_5\ : std_logic;
signal \b2v_inst11.countZ0Z_7\ : std_logic;
signal \b2v_inst11.mult1_un117_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5536_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_6\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_7\ : std_logic;
signal \b2v_inst11.countZ0Z_8\ : std_logic;
signal \b2v_inst11.mult1_un110_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5537_i\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \b2v_inst11.countZ0Z_9\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_i_8\ : std_logic;
signal \b2v_inst11.N_5538_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_8\ : std_logic;
signal \b2v_inst11.countZ0Z_10\ : std_logic;
signal \b2v_inst11.N_5539_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_9\ : std_logic;
signal \b2v_inst11.countZ0Z_11\ : std_logic;
signal \b2v_inst11.N_5540_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_10\ : std_logic;
signal \b2v_inst11.countZ0Z_12\ : std_logic;
signal \b2v_inst11.N_5541_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_11\ : std_logic;
signal \b2v_inst11.countZ0Z_13\ : std_logic;
signal \b2v_inst11.N_5542_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_12\ : std_logic;
signal \b2v_inst11.countZ0Z_14\ : std_logic;
signal \b2v_inst11.N_5543_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_13\ : std_logic;
signal \b2v_inst11.countZ0Z_15\ : std_logic;
signal \b2v_inst11.N_5544_i\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_14\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i_8\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_1\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_7\ : std_logic;
signal \b2v_inst11.dutycycle\ : std_logic;
signal \b2v_inst11.mult1_un54_sum\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \V33S_OK_c\ : std_logic;
signal \V5S_OK_c\ : std_logic;
signal \VCCIN_EN_c\ : std_logic;
signal \b2v_inst6.N_276_0_cascade_\ : std_logic;
signal \VR_READY_VCCINAUX_c\ : std_logic;
signal \VR_READY_VCCIN_c\ : std_logic;
signal \b2v_inst6.N_192_cascade_\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_ok_0\ : std_logic;
signal \b2v_inst6.curr_state_RNIUL1J2Z0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.N_276_0\ : std_logic;
signal \N_15_i_0_a4_1_N_3L3_1\ : std_logic;
signal \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\ : std_logic;
signal \N_222\ : std_logic;
signal \b2v_inst11.dutycycleZ0Z_0\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_0\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_2_s\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_1\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_s_7\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un159_sum_cry_5_s\ : std_logic;
signal \G_2836\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_axb_6\ : std_logic;
signal \b2v_inst11.mult1_un166_sum_cry_5\ : std_logic;
signal \b2v_inst11.un85_clk_100khz_0\ : std_logic;
signal \bfn_12_1_0_\ : std_logic;
signal \b2v_inst6.countZ0Z_2\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_1\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4\ : std_logic;
signal \b2v_inst6.countZ0Z_6\ : std_logic;
signal \b2v_inst6.count_rst_8\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_5\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8\ : std_logic;
signal \bfn_12_2_0_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_11\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_12\ : std_logic;
signal \b2v_inst6.countZ0Z_14\ : std_logic;
signal \b2v_inst6.count_rst_0\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_13\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_14\ : std_logic;
signal \b2v_inst6.count_0_13\ : std_logic;
signal \b2v_inst6.count_rst_1\ : std_logic;
signal \b2v_inst6.countZ0Z_13\ : std_logic;
signal \b2v_inst6.count_0_5\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_5_cascade_\ : std_logic;
signal \b2v_inst6.count_rst_9\ : std_logic;
signal \b2v_inst6.count_rst_5\ : std_logic;
signal \b2v_inst6.countZ0Z_9_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_5\ : std_logic;
signal \b2v_inst6.countZ0Z_9\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \b2v_inst6.count_0_9\ : std_logic;
signal \b2v_inst6.countZ0Z_10\ : std_logic;
signal \b2v_inst6.countZ0Z_10_cascade_\ : std_logic;
signal \b2v_inst6.count_0_12\ : std_logic;
signal \b2v_inst6.count_rst_2\ : std_logic;
signal \b2v_inst6.countZ0Z_12\ : std_logic;
signal \b2v_inst6.count_rst_10_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_4\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_4_cascade_\ : std_logic;
signal \b2v_inst6.count_0_4\ : std_logic;
signal \b2v_inst6.count_rst_4\ : std_logic;
signal \b2v_inst6.count_0_10\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \b2v_inst6.count_0_7\ : std_logic;
signal \b2v_inst6.count_rst_7_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_7\ : std_logic;
signal \b2v_inst6.count_rst\ : std_logic;
signal \b2v_inst6.count_0_15\ : std_logic;
signal \b2v_inst6.count_rst_12\ : std_logic;
signal \b2v_inst6.count_0_2\ : std_logic;
signal \b2v_inst6.count_rst_6\ : std_logic;
signal \b2v_inst6.countZ0Z_8\ : std_logic;
signal \b2v_inst6.countZ0Z_8_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \b2v_inst6.count_0_8\ : std_logic;
signal \b2v_inst6.count_rst_11_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \b2v_inst6.countZ0Z_3_cascade_\ : std_logic;
signal \b2v_inst6.count_0_3\ : std_logic;
signal \b2v_inst6.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \b2v_inst6.N_394_cascade_\ : std_logic;
signal \b2v_inst6.count_0_11\ : std_logic;
signal \b2v_inst6.count_rst_3_cascade_\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_1\ : std_logic;
signal \b2v_inst6.un2_count_1_axb_1_cascade_\ : std_logic;
signal \V1P8A_OK_c\ : std_logic;
signal \V33A_OK_c\ : std_logic;
signal \V5A_OK_c\ : std_logic;
signal \VCCST_CPU_OK_c\ : std_logic;
signal \N_1661\ : std_logic;
signal \b2v_inst6.count_0_1\ : std_logic;
signal \b2v_inst6.count_RNI_0_1\ : std_logic;
signal \b2v_inst6.countZ0Z_15\ : std_logic;
signal \b2v_inst6.countZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.countZ0Z_11\ : std_logic;
signal \b2v_inst6.count_1_i_a3_8_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_9_0\ : std_logic;
signal \b2v_inst6.count_1_i_a3_7_0_cascade_\ : std_logic;
signal \b2v_inst6.count_1_i_a3_10_0\ : std_logic;
signal \b2v_inst6.N_389\ : std_logic;
signal \b2v_inst6.N_389_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i_8\ : std_logic;
signal \b2v_inst6.count_en\ : std_logic;
signal \b2v_inst6.count_RNIM2CM2Z0Z_0\ : std_logic;
signal \b2v_inst6.count_en_cascade_\ : std_logic;
signal \b2v_inst6.count_0_0\ : std_logic;
signal \b2v_inst6.countZ0Z_0\ : std_logic;
signal \b2v_inst11.mult1_un96_sum\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un103_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un96_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum\ : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un89_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum\ : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un82_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_2\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_3_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_3\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_4_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_4\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_5_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_5\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_cry_6_s\ : std_logic;
signal \b2v_inst11.mult1_un61_sum_i_0_8\ : std_logic;
signal \b2v_inst11.mult1_un75_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_6\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_axb_8\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_cry_7\ : std_logic;
signal \b2v_inst11.mult1_un68_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_s_8\ : std_logic;
signal \b2v_inst11.mult1_un54_sum_i_8\ : std_logic;
signal \b2v_inst6.N_192\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \b2v_inst6.count_0_sqmuxa\ : std_logic;
signal \b2v_inst6.curr_state_1_0\ : std_logic;
signal \SYNTHESIZED_WIRE_1keep_3\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_0\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_RNIUL1J2Z0Z_0\ : std_logic;
signal \b2v_inst6.curr_state_7_0\ : std_logic;
signal \b2v_inst6.N_2937_i\ : std_logic;
signal \b2v_inst6.curr_stateZ0Z_1\ : std_logic;
signal \b2v_inst6.N_394\ : std_logic;
signal \b2v_inst6.m6_i_a3\ : std_logic;
signal \b2v_inst6.N_241\ : std_logic;
signal \b2v_inst6.m6_i_a3_cascade_\ : std_logic;
signal \b2v_inst6.curr_state_1_1\ : std_logic;
signal \FPGA_OSC_0_c_g\ : std_logic;
signal \N_606_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \FPGA_OSC_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;

begin
    \FPGA_OSC_wire\ <= FPGA_OSC;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \V5A_OK_wire\ <= V5A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V5S_ENn <= \V5S_ENn_wire\;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    \SLP_S3n_wire\ <= SLP_S3n;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    VCCST_EN <= \VCCST_EN_wire\;
    \VPP_OK_wire\ <= VPP_OK;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    VPP_EN <= \VPP_EN_wire\;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    V33S_ENn <= \V33S_ENn_wire\;
    RSMRSTn <= \RSMRSTn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    DSW_PWROK <= \DSW_PWROK_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    VDDQ_EN <= \VDDQ_EN_wire\;
    V5A_EN <= \V5A_EN_wire\;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    V33A_ENn <= \V33A_ENn_wire\;
    \V5S_OK_wire\ <= V5S_OK;
    \V33A_OK_wire\ <= V33A_OK;

    \FPGA_OSC_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__37127\,
            GLOBALBUFFEROUTPUT => \FPGA_OSC_0_c_g\
        );

    \FPGA_OSC_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37129\,
            DIN => \N__37128\,
            DOUT => \N__37127\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \FPGA_OSC_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37129\,
            PADOUT => \N__37128\,
            PADIN => \N__37127\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V1P8A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37118\,
            DIN => \N__37117\,
            DOUT => \N__37116\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \V1P8A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37118\,
            PADOUT => \N__37117\,
            PADIN => \N__37116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V1P8A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37109\,
            DIN => \N__37108\,
            DOUT => \N__37107\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \V5A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37109\,
            PADOUT => \N__37108\,
            PADIN => \N__37107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCH_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37100\,
            DIN => \N__37099\,
            DOUT => \N__37098\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \PCH_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37100\,
            PADOUT => \N__37099\,
            PADIN => \N__37098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18636\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCIN_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37091\,
            DIN => \N__37090\,
            DOUT => \N__37089\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \VCCIN_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37091\,
            PADOUT => \N__37090\,
            PADIN => \N__37089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33S_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37082\,
            DIN => \N__37081\,
            DOUT => \N__37080\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \V33S_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37082\,
            PADOUT => \N__37081\,
            PADIN => \N__37080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33S_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5S_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37073\,
            DIN => \N__37072\,
            DOUT => \N__37071\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \V5S_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37073\,
            PADOUT => \N__37072\,
            PADIN => \N__37071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_S4n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37064\,
            DIN => \N__37063\,
            DOUT => \N__37062\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \SLP_S4n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37064\,
            PADOUT => \N__37063\,
            PADIN => \N__37062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SLP_S4n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VR_READY_VCCINAUX_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37055\,
            DIN => \N__37054\,
            DOUT => \N__37053\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \VR_READY_VCCINAUX_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37055\,
            PADOUT => \N__37054\,
            PADIN => \N__37053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VR_READY_VCCINAUX_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SLP_S3n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37046\,
            DIN => \N__37045\,
            DOUT => \N__37044\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \SLP_S3n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37046\,
            PADOUT => \N__37045\,
            PADIN => \N__37044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SLP_S3n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_PWRGD_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37037\,
            DIN => \N__37036\,
            DOUT => \N__37035\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \VCCST_PWRGD_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37037\,
            PADOUT => \N__37036\,
            PADIN => \N__37035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18640\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HDA_SDO_ATP_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37028\,
            DIN => \N__37027\,
            DOUT => \N__37026\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \HDA_SDO_ATP_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37028\,
            PADOUT => \N__37027\,
            PADIN => \N__37026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20227\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37019\,
            DIN => \N__37018\,
            DOUT => \N__37017\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \VCCST_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__37019\,
            PADOUT => \N__37018\,
            PADIN => \N__37017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19873\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VPP_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37010\,
            DIN => \N__37009\,
            DOUT => \N__37008\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \VPP_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37010\,
            PADOUT => \N__37009\,
            PADIN => \N__37008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VPP_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO_FPGA_SoC_1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__37001\,
            DIN => \N__37000\,
            DOUT => \N__36999\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \GPIO_FPGA_SoC_1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__37001\,
            PADOUT => \N__37000\,
            PADIN => \N__36999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \GPIO_FPGA_SoC_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCST_CPU_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36992\,
            DIN => \N__36991\,
            DOUT => \N__36990\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \VCCST_CPU_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36992\,
            PADOUT => \N__36991\,
            PADIN => \N__36990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VCCST_CPU_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \GPIO_FPGA_SoC_4_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36983\,
            DIN => \N__36982\,
            DOUT => \N__36981\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \GPIO_FPGA_SoC_4_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36983\,
            PADOUT => \N__36982\,
            PADIN => \N__36981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \GPIO_FPGA_SoC_4_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VPP_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36974\,
            DIN => \N__36973\,
            DOUT => \N__36972\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \VPP_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36974\,
            PADOUT => \N__36973\,
            PADIN => \N__36972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PWRBTN_LED_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36965\,
            DIN => \N__36964\,
            DOUT => \N__36963\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \PWRBTN_LED_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36965\,
            PADOUT => \N__36964\,
            PADIN => \N__36963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24946\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33S_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36956\,
            DIN => \N__36955\,
            DOUT => \N__36954\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \V33S_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36956\,
            PADOUT => \N__36955\,
            PADIN => \N__36954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33792\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RSMRSTn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36947\,
            DIN => \N__36946\,
            DOUT => \N__36945\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \RSMRSTn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36947\,
            PADOUT => \N__36946\,
            PADIN => \N__36945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23911\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V1P8A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36938\,
            DIN => \N__36937\,
            DOUT => \N__36936\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \V1P8A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36938\,
            PADOUT => \N__36937\,
            PADIN => \N__36936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VDDQ_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36929\,
            DIN => \N__36928\,
            DOUT => \N__36927\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \VDDQ_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36929\,
            PADOUT => \N__36928\,
            PADIN => \N__36927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VDDQ_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DSW_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36920\,
            DIN => \N__36919\,
            DOUT => \N__36918\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \DSW_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36920\,
            PADOUT => \N__36919\,
            PADIN => \N__36918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22351\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SYS_PWROK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36911\,
            DIN => \N__36910\,
            DOUT => \N__36909\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \SYS_PWROK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36911\,
            PADOUT => \N__36910\,
            PADIN => \N__36909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18635\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33DSW_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36902\,
            DIN => \N__36901\,
            DOUT => \N__36900\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \V33DSW_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36902\,
            PADOUT => \N__36901\,
            PADIN => \N__36900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33DSW_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VR_READY_VCCIN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36893\,
            DIN => \N__36892\,
            DOUT => \N__36891\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \VR_READY_VCCIN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36893\,
            PADOUT => \N__36892\,
            PADIN => \N__36891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \VR_READY_VCCIN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VDDQ_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36884\,
            DIN => \N__36883\,
            DOUT => \N__36882\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \VDDQ_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36884\,
            PADOUT => \N__36883\,
            PADIN => \N__36882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16966\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5A_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36875\,
            DIN => \N__36874\,
            DOUT => \N__36873\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \V5A_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36875\,
            PADOUT => \N__36874\,
            PADIN => \N__36873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__30442\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VCCINAUX_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36866\,
            DIN => \N__36865\,
            DOUT => \N__36864\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \VCCINAUX_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36866\,
            PADOUT => \N__36865\,
            PADIN => \N__36864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33403\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33A_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36857\,
            DIN => \N__36856\,
            DOUT => \N__36855\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \V33A_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__36857\,
            PADOUT => \N__36856\,
            PADIN => \N__36855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V5S_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36848\,
            DIN => \N__36847\,
            DOUT => \N__36846\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \V5S_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36848\,
            PADOUT => \N__36847\,
            PADIN => \N__36846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V5S_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \V33A_OK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__36839\,
            DIN => \N__36838\,
            DOUT => \N__36837\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \V33A_OK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__36839\,
            PADOUT => \N__36838\,
            PADIN => \N__36837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \V33A_OK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__8612\ : InMux
    port map (
            O => \N__36820\,
            I => \N__36814\
        );

    \I__8611\ : InMux
    port map (
            O => \N__36819\,
            I => \N__36807\
        );

    \I__8610\ : InMux
    port map (
            O => \N__36818\,
            I => \N__36807\
        );

    \I__8609\ : InMux
    port map (
            O => \N__36817\,
            I => \N__36807\
        );

    \I__8608\ : LocalMux
    port map (
            O => \N__36814\,
            I => \b2v_inst6.N_2937_i\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__36807\,
            I => \b2v_inst6.N_2937_i\
        );

    \I__8606\ : InMux
    port map (
            O => \N__36802\,
            I => \N__36793\
        );

    \I__8605\ : InMux
    port map (
            O => \N__36801\,
            I => \N__36793\
        );

    \I__8604\ : InMux
    port map (
            O => \N__36800\,
            I => \N__36793\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__36793\,
            I => \b2v_inst6.curr_stateZ0Z_1\
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__36790\,
            I => \N__36784\
        );

    \I__8601\ : CascadeMux
    port map (
            O => \N__36789\,
            I => \N__36778\
        );

    \I__8600\ : CascadeMux
    port map (
            O => \N__36788\,
            I => \N__36775\
        );

    \I__8599\ : InMux
    port map (
            O => \N__36787\,
            I => \N__36765\
        );

    \I__8598\ : InMux
    port map (
            O => \N__36784\,
            I => \N__36765\
        );

    \I__8597\ : InMux
    port map (
            O => \N__36783\,
            I => \N__36762\
        );

    \I__8596\ : InMux
    port map (
            O => \N__36782\,
            I => \N__36753\
        );

    \I__8595\ : InMux
    port map (
            O => \N__36781\,
            I => \N__36753\
        );

    \I__8594\ : InMux
    port map (
            O => \N__36778\,
            I => \N__36742\
        );

    \I__8593\ : InMux
    port map (
            O => \N__36775\,
            I => \N__36742\
        );

    \I__8592\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36742\
        );

    \I__8591\ : InMux
    port map (
            O => \N__36773\,
            I => \N__36742\
        );

    \I__8590\ : InMux
    port map (
            O => \N__36772\,
            I => \N__36742\
        );

    \I__8589\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36737\
        );

    \I__8588\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36737\
        );

    \I__8587\ : LocalMux
    port map (
            O => \N__36765\,
            I => \N__36732\
        );

    \I__8586\ : LocalMux
    port map (
            O => \N__36762\,
            I => \N__36732\
        );

    \I__8585\ : InMux
    port map (
            O => \N__36761\,
            I => \N__36727\
        );

    \I__8584\ : InMux
    port map (
            O => \N__36760\,
            I => \N__36727\
        );

    \I__8583\ : InMux
    port map (
            O => \N__36759\,
            I => \N__36722\
        );

    \I__8582\ : InMux
    port map (
            O => \N__36758\,
            I => \N__36722\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__36753\,
            I => \N__36713\
        );

    \I__8580\ : LocalMux
    port map (
            O => \N__36742\,
            I => \N__36713\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__36737\,
            I => \N__36713\
        );

    \I__8578\ : Span12Mux_s8_v
    port map (
            O => \N__36732\,
            I => \N__36713\
        );

    \I__8577\ : LocalMux
    port map (
            O => \N__36727\,
            I => \b2v_inst6.N_394\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__36722\,
            I => \b2v_inst6.N_394\
        );

    \I__8575\ : Odrv12
    port map (
            O => \N__36713\,
            I => \b2v_inst6.N_394\
        );

    \I__8574\ : InMux
    port map (
            O => \N__36706\,
            I => \N__36703\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__36703\,
            I => \b2v_inst6.m6_i_a3\
        );

    \I__8572\ : CascadeMux
    port map (
            O => \N__36700\,
            I => \N__36696\
        );

    \I__8571\ : InMux
    port map (
            O => \N__36699\,
            I => \N__36693\
        );

    \I__8570\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36689\
        );

    \I__8569\ : LocalMux
    port map (
            O => \N__36693\,
            I => \N__36686\
        );

    \I__8568\ : InMux
    port map (
            O => \N__36692\,
            I => \N__36683\
        );

    \I__8567\ : LocalMux
    port map (
            O => \N__36689\,
            I => \N__36678\
        );

    \I__8566\ : Span4Mux_v
    port map (
            O => \N__36686\,
            I => \N__36678\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__36683\,
            I => \b2v_inst6.N_241\
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__36678\,
            I => \b2v_inst6.N_241\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__36673\,
            I => \b2v_inst6.m6_i_a3_cascade_\
        );

    \I__8562\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36667\
        );

    \I__8561\ : LocalMux
    port map (
            O => \N__36667\,
            I => \b2v_inst6.curr_state_1_1\
        );

    \I__8560\ : ClkMux
    port map (
            O => \N__36664\,
            I => \N__36415\
        );

    \I__8559\ : ClkMux
    port map (
            O => \N__36663\,
            I => \N__36415\
        );

    \I__8558\ : ClkMux
    port map (
            O => \N__36662\,
            I => \N__36415\
        );

    \I__8557\ : ClkMux
    port map (
            O => \N__36661\,
            I => \N__36415\
        );

    \I__8556\ : ClkMux
    port map (
            O => \N__36660\,
            I => \N__36415\
        );

    \I__8555\ : ClkMux
    port map (
            O => \N__36659\,
            I => \N__36415\
        );

    \I__8554\ : ClkMux
    port map (
            O => \N__36658\,
            I => \N__36415\
        );

    \I__8553\ : ClkMux
    port map (
            O => \N__36657\,
            I => \N__36415\
        );

    \I__8552\ : ClkMux
    port map (
            O => \N__36656\,
            I => \N__36415\
        );

    \I__8551\ : ClkMux
    port map (
            O => \N__36655\,
            I => \N__36415\
        );

    \I__8550\ : ClkMux
    port map (
            O => \N__36654\,
            I => \N__36415\
        );

    \I__8549\ : ClkMux
    port map (
            O => \N__36653\,
            I => \N__36415\
        );

    \I__8548\ : ClkMux
    port map (
            O => \N__36652\,
            I => \N__36415\
        );

    \I__8547\ : ClkMux
    port map (
            O => \N__36651\,
            I => \N__36415\
        );

    \I__8546\ : ClkMux
    port map (
            O => \N__36650\,
            I => \N__36415\
        );

    \I__8545\ : ClkMux
    port map (
            O => \N__36649\,
            I => \N__36415\
        );

    \I__8544\ : ClkMux
    port map (
            O => \N__36648\,
            I => \N__36415\
        );

    \I__8543\ : ClkMux
    port map (
            O => \N__36647\,
            I => \N__36415\
        );

    \I__8542\ : ClkMux
    port map (
            O => \N__36646\,
            I => \N__36415\
        );

    \I__8541\ : ClkMux
    port map (
            O => \N__36645\,
            I => \N__36415\
        );

    \I__8540\ : ClkMux
    port map (
            O => \N__36644\,
            I => \N__36415\
        );

    \I__8539\ : ClkMux
    port map (
            O => \N__36643\,
            I => \N__36415\
        );

    \I__8538\ : ClkMux
    port map (
            O => \N__36642\,
            I => \N__36415\
        );

    \I__8537\ : ClkMux
    port map (
            O => \N__36641\,
            I => \N__36415\
        );

    \I__8536\ : ClkMux
    port map (
            O => \N__36640\,
            I => \N__36415\
        );

    \I__8535\ : ClkMux
    port map (
            O => \N__36639\,
            I => \N__36415\
        );

    \I__8534\ : ClkMux
    port map (
            O => \N__36638\,
            I => \N__36415\
        );

    \I__8533\ : ClkMux
    port map (
            O => \N__36637\,
            I => \N__36415\
        );

    \I__8532\ : ClkMux
    port map (
            O => \N__36636\,
            I => \N__36415\
        );

    \I__8531\ : ClkMux
    port map (
            O => \N__36635\,
            I => \N__36415\
        );

    \I__8530\ : ClkMux
    port map (
            O => \N__36634\,
            I => \N__36415\
        );

    \I__8529\ : ClkMux
    port map (
            O => \N__36633\,
            I => \N__36415\
        );

    \I__8528\ : ClkMux
    port map (
            O => \N__36632\,
            I => \N__36415\
        );

    \I__8527\ : ClkMux
    port map (
            O => \N__36631\,
            I => \N__36415\
        );

    \I__8526\ : ClkMux
    port map (
            O => \N__36630\,
            I => \N__36415\
        );

    \I__8525\ : ClkMux
    port map (
            O => \N__36629\,
            I => \N__36415\
        );

    \I__8524\ : ClkMux
    port map (
            O => \N__36628\,
            I => \N__36415\
        );

    \I__8523\ : ClkMux
    port map (
            O => \N__36627\,
            I => \N__36415\
        );

    \I__8522\ : ClkMux
    port map (
            O => \N__36626\,
            I => \N__36415\
        );

    \I__8521\ : ClkMux
    port map (
            O => \N__36625\,
            I => \N__36415\
        );

    \I__8520\ : ClkMux
    port map (
            O => \N__36624\,
            I => \N__36415\
        );

    \I__8519\ : ClkMux
    port map (
            O => \N__36623\,
            I => \N__36415\
        );

    \I__8518\ : ClkMux
    port map (
            O => \N__36622\,
            I => \N__36415\
        );

    \I__8517\ : ClkMux
    port map (
            O => \N__36621\,
            I => \N__36415\
        );

    \I__8516\ : ClkMux
    port map (
            O => \N__36620\,
            I => \N__36415\
        );

    \I__8515\ : ClkMux
    port map (
            O => \N__36619\,
            I => \N__36415\
        );

    \I__8514\ : ClkMux
    port map (
            O => \N__36618\,
            I => \N__36415\
        );

    \I__8513\ : ClkMux
    port map (
            O => \N__36617\,
            I => \N__36415\
        );

    \I__8512\ : ClkMux
    port map (
            O => \N__36616\,
            I => \N__36415\
        );

    \I__8511\ : ClkMux
    port map (
            O => \N__36615\,
            I => \N__36415\
        );

    \I__8510\ : ClkMux
    port map (
            O => \N__36614\,
            I => \N__36415\
        );

    \I__8509\ : ClkMux
    port map (
            O => \N__36613\,
            I => \N__36415\
        );

    \I__8508\ : ClkMux
    port map (
            O => \N__36612\,
            I => \N__36415\
        );

    \I__8507\ : ClkMux
    port map (
            O => \N__36611\,
            I => \N__36415\
        );

    \I__8506\ : ClkMux
    port map (
            O => \N__36610\,
            I => \N__36415\
        );

    \I__8505\ : ClkMux
    port map (
            O => \N__36609\,
            I => \N__36415\
        );

    \I__8504\ : ClkMux
    port map (
            O => \N__36608\,
            I => \N__36415\
        );

    \I__8503\ : ClkMux
    port map (
            O => \N__36607\,
            I => \N__36415\
        );

    \I__8502\ : ClkMux
    port map (
            O => \N__36606\,
            I => \N__36415\
        );

    \I__8501\ : ClkMux
    port map (
            O => \N__36605\,
            I => \N__36415\
        );

    \I__8500\ : ClkMux
    port map (
            O => \N__36604\,
            I => \N__36415\
        );

    \I__8499\ : ClkMux
    port map (
            O => \N__36603\,
            I => \N__36415\
        );

    \I__8498\ : ClkMux
    port map (
            O => \N__36602\,
            I => \N__36415\
        );

    \I__8497\ : ClkMux
    port map (
            O => \N__36601\,
            I => \N__36415\
        );

    \I__8496\ : ClkMux
    port map (
            O => \N__36600\,
            I => \N__36415\
        );

    \I__8495\ : ClkMux
    port map (
            O => \N__36599\,
            I => \N__36415\
        );

    \I__8494\ : ClkMux
    port map (
            O => \N__36598\,
            I => \N__36415\
        );

    \I__8493\ : ClkMux
    port map (
            O => \N__36597\,
            I => \N__36415\
        );

    \I__8492\ : ClkMux
    port map (
            O => \N__36596\,
            I => \N__36415\
        );

    \I__8491\ : ClkMux
    port map (
            O => \N__36595\,
            I => \N__36415\
        );

    \I__8490\ : ClkMux
    port map (
            O => \N__36594\,
            I => \N__36415\
        );

    \I__8489\ : ClkMux
    port map (
            O => \N__36593\,
            I => \N__36415\
        );

    \I__8488\ : ClkMux
    port map (
            O => \N__36592\,
            I => \N__36415\
        );

    \I__8487\ : ClkMux
    port map (
            O => \N__36591\,
            I => \N__36415\
        );

    \I__8486\ : ClkMux
    port map (
            O => \N__36590\,
            I => \N__36415\
        );

    \I__8485\ : ClkMux
    port map (
            O => \N__36589\,
            I => \N__36415\
        );

    \I__8484\ : ClkMux
    port map (
            O => \N__36588\,
            I => \N__36415\
        );

    \I__8483\ : ClkMux
    port map (
            O => \N__36587\,
            I => \N__36415\
        );

    \I__8482\ : ClkMux
    port map (
            O => \N__36586\,
            I => \N__36415\
        );

    \I__8481\ : ClkMux
    port map (
            O => \N__36585\,
            I => \N__36415\
        );

    \I__8480\ : ClkMux
    port map (
            O => \N__36584\,
            I => \N__36415\
        );

    \I__8479\ : ClkMux
    port map (
            O => \N__36583\,
            I => \N__36415\
        );

    \I__8478\ : ClkMux
    port map (
            O => \N__36582\,
            I => \N__36415\
        );

    \I__8477\ : GlobalMux
    port map (
            O => \N__36415\,
            I => \N__36412\
        );

    \I__8476\ : gio2CtrlBuf
    port map (
            O => \N__36412\,
            I => \FPGA_OSC_0_c_g\
        );

    \I__8475\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36397\
        );

    \I__8474\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36394\
        );

    \I__8473\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36391\
        );

    \I__8472\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36384\
        );

    \I__8471\ : InMux
    port map (
            O => \N__36405\,
            I => \N__36384\
        );

    \I__8470\ : InMux
    port map (
            O => \N__36404\,
            I => \N__36384\
        );

    \I__8469\ : InMux
    port map (
            O => \N__36403\,
            I => \N__36381\
        );

    \I__8468\ : InMux
    port map (
            O => \N__36402\,
            I => \N__36376\
        );

    \I__8467\ : InMux
    port map (
            O => \N__36401\,
            I => \N__36376\
        );

    \I__8466\ : InMux
    port map (
            O => \N__36400\,
            I => \N__36373\
        );

    \I__8465\ : LocalMux
    port map (
            O => \N__36397\,
            I => \N__36370\
        );

    \I__8464\ : LocalMux
    port map (
            O => \N__36394\,
            I => \N__36352\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__36391\,
            I => \N__36349\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__36384\,
            I => \N__36346\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__36381\,
            I => \N__36343\
        );

    \I__8460\ : LocalMux
    port map (
            O => \N__36376\,
            I => \N__36340\
        );

    \I__8459\ : LocalMux
    port map (
            O => \N__36373\,
            I => \N__36337\
        );

    \I__8458\ : Glb2LocalMux
    port map (
            O => \N__36370\,
            I => \N__36292\
        );

    \I__8457\ : CEMux
    port map (
            O => \N__36369\,
            I => \N__36292\
        );

    \I__8456\ : CEMux
    port map (
            O => \N__36368\,
            I => \N__36292\
        );

    \I__8455\ : CEMux
    port map (
            O => \N__36367\,
            I => \N__36292\
        );

    \I__8454\ : CEMux
    port map (
            O => \N__36366\,
            I => \N__36292\
        );

    \I__8453\ : CEMux
    port map (
            O => \N__36365\,
            I => \N__36292\
        );

    \I__8452\ : CEMux
    port map (
            O => \N__36364\,
            I => \N__36292\
        );

    \I__8451\ : CEMux
    port map (
            O => \N__36363\,
            I => \N__36292\
        );

    \I__8450\ : CEMux
    port map (
            O => \N__36362\,
            I => \N__36292\
        );

    \I__8449\ : CEMux
    port map (
            O => \N__36361\,
            I => \N__36292\
        );

    \I__8448\ : CEMux
    port map (
            O => \N__36360\,
            I => \N__36292\
        );

    \I__8447\ : CEMux
    port map (
            O => \N__36359\,
            I => \N__36292\
        );

    \I__8446\ : CEMux
    port map (
            O => \N__36358\,
            I => \N__36292\
        );

    \I__8445\ : CEMux
    port map (
            O => \N__36357\,
            I => \N__36292\
        );

    \I__8444\ : CEMux
    port map (
            O => \N__36356\,
            I => \N__36292\
        );

    \I__8443\ : CEMux
    port map (
            O => \N__36355\,
            I => \N__36292\
        );

    \I__8442\ : Glb2LocalMux
    port map (
            O => \N__36352\,
            I => \N__36292\
        );

    \I__8441\ : Glb2LocalMux
    port map (
            O => \N__36349\,
            I => \N__36292\
        );

    \I__8440\ : Glb2LocalMux
    port map (
            O => \N__36346\,
            I => \N__36292\
        );

    \I__8439\ : Glb2LocalMux
    port map (
            O => \N__36343\,
            I => \N__36292\
        );

    \I__8438\ : Glb2LocalMux
    port map (
            O => \N__36340\,
            I => \N__36292\
        );

    \I__8437\ : Glb2LocalMux
    port map (
            O => \N__36337\,
            I => \N__36292\
        );

    \I__8436\ : GlobalMux
    port map (
            O => \N__36292\,
            I => \N__36289\
        );

    \I__8435\ : gio2CtrlBuf
    port map (
            O => \N__36289\,
            I => \N_606_g\
        );

    \I__8434\ : InMux
    port map (
            O => \N__36286\,
            I => \b2v_inst11.mult1_un68_sum_cry_5\
        );

    \I__8433\ : InMux
    port map (
            O => \N__36283\,
            I => \N__36280\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__36280\,
            I => \N__36277\
        );

    \I__8431\ : Odrv4
    port map (
            O => \N__36277\,
            I => \b2v_inst11.mult1_un61_sum_cry_6_s\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__36274\,
            I => \N__36270\
        );

    \I__8429\ : CascadeMux
    port map (
            O => \N__36273\,
            I => \N__36266\
        );

    \I__8428\ : InMux
    port map (
            O => \N__36270\,
            I => \N__36259\
        );

    \I__8427\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36259\
        );

    \I__8426\ : InMux
    port map (
            O => \N__36266\,
            I => \N__36259\
        );

    \I__8425\ : LocalMux
    port map (
            O => \N__36259\,
            I => \b2v_inst11.mult1_un61_sum_i_0_8\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__36256\,
            I => \N__36253\
        );

    \I__8423\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36250\
        );

    \I__8422\ : LocalMux
    port map (
            O => \N__36250\,
            I => \b2v_inst11.mult1_un75_sum_axb_8\
        );

    \I__8421\ : InMux
    port map (
            O => \N__36247\,
            I => \b2v_inst11.mult1_un68_sum_cry_6\
        );

    \I__8420\ : CascadeMux
    port map (
            O => \N__36244\,
            I => \N__36241\
        );

    \I__8419\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36238\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__36238\,
            I => \b2v_inst11.mult1_un68_sum_axb_8\
        );

    \I__8417\ : InMux
    port map (
            O => \N__36235\,
            I => \b2v_inst11.mult1_un68_sum_cry_7\
        );

    \I__8416\ : InMux
    port map (
            O => \N__36232\,
            I => \N__36227\
        );

    \I__8415\ : CascadeMux
    port map (
            O => \N__36231\,
            I => \N__36223\
        );

    \I__8414\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36219\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__36227\,
            I => \N__36216\
        );

    \I__8412\ : InMux
    port map (
            O => \N__36226\,
            I => \N__36211\
        );

    \I__8411\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36211\
        );

    \I__8410\ : InMux
    port map (
            O => \N__36222\,
            I => \N__36208\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36205\
        );

    \I__8408\ : Odrv12
    port map (
            O => \N__36216\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__8407\ : LocalMux
    port map (
            O => \N__36211\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__36208\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__36205\,
            I => \b2v_inst11.mult1_un68_sum_s_8\
        );

    \I__8404\ : CascadeMux
    port map (
            O => \N__36196\,
            I => \N__36191\
        );

    \I__8403\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36188\
        );

    \I__8402\ : InMux
    port map (
            O => \N__36194\,
            I => \N__36182\
        );

    \I__8401\ : InMux
    port map (
            O => \N__36191\,
            I => \N__36182\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__36188\,
            I => \N__36179\
        );

    \I__8399\ : InMux
    port map (
            O => \N__36187\,
            I => \N__36176\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__36182\,
            I => \N__36171\
        );

    \I__8397\ : Span4Mux_s0_h
    port map (
            O => \N__36179\,
            I => \N__36171\
        );

    \I__8396\ : LocalMux
    port map (
            O => \N__36176\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__36171\,
            I => \b2v_inst11.mult1_un54_sum_s_8\
        );

    \I__8394\ : CascadeMux
    port map (
            O => \N__36166\,
            I => \N__36162\
        );

    \I__8393\ : CascadeMux
    port map (
            O => \N__36165\,
            I => \N__36158\
        );

    \I__8392\ : InMux
    port map (
            O => \N__36162\,
            I => \N__36151\
        );

    \I__8391\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36151\
        );

    \I__8390\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36151\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__36151\,
            I => \b2v_inst11.mult1_un54_sum_i_8\
        );

    \I__8388\ : InMux
    port map (
            O => \N__36148\,
            I => \N__36141\
        );

    \I__8387\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36141\
        );

    \I__8386\ : InMux
    port map (
            O => \N__36146\,
            I => \N__36138\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__36141\,
            I => \b2v_inst6.N_192\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__36138\,
            I => \b2v_inst6.N_192\
        );

    \I__8383\ : CascadeMux
    port map (
            O => \N__36133\,
            I => \b2v_inst6.curr_stateZ0Z_0_cascade_\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__36130\,
            I => \N__36125\
        );

    \I__8381\ : SRMux
    port map (
            O => \N__36129\,
            I => \N__36121\
        );

    \I__8380\ : SRMux
    port map (
            O => \N__36128\,
            I => \N__36115\
        );

    \I__8379\ : InMux
    port map (
            O => \N__36125\,
            I => \N__36107\
        );

    \I__8378\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36107\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__36121\,
            I => \N__36104\
        );

    \I__8376\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36099\
        );

    \I__8375\ : SRMux
    port map (
            O => \N__36119\,
            I => \N__36099\
        );

    \I__8374\ : SRMux
    port map (
            O => \N__36118\,
            I => \N__36096\
        );

    \I__8373\ : LocalMux
    port map (
            O => \N__36115\,
            I => \N__36093\
        );

    \I__8372\ : SRMux
    port map (
            O => \N__36114\,
            I => \N__36090\
        );

    \I__8371\ : InMux
    port map (
            O => \N__36113\,
            I => \N__36077\
        );

    \I__8370\ : InMux
    port map (
            O => \N__36112\,
            I => \N__36077\
        );

    \I__8369\ : LocalMux
    port map (
            O => \N__36107\,
            I => \N__36067\
        );

    \I__8368\ : Span4Mux_s1_v
    port map (
            O => \N__36104\,
            I => \N__36067\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__36099\,
            I => \N__36067\
        );

    \I__8366\ : LocalMux
    port map (
            O => \N__36096\,
            I => \N__36067\
        );

    \I__8365\ : Span4Mux_v
    port map (
            O => \N__36093\,
            I => \N__36062\
        );

    \I__8364\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36062\
        );

    \I__8363\ : InMux
    port map (
            O => \N__36089\,
            I => \N__36057\
        );

    \I__8362\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36057\
        );

    \I__8361\ : InMux
    port map (
            O => \N__36087\,
            I => \N__36050\
        );

    \I__8360\ : InMux
    port map (
            O => \N__36086\,
            I => \N__36050\
        );

    \I__8359\ : InMux
    port map (
            O => \N__36085\,
            I => \N__36050\
        );

    \I__8358\ : InMux
    port map (
            O => \N__36084\,
            I => \N__36043\
        );

    \I__8357\ : InMux
    port map (
            O => \N__36083\,
            I => \N__36043\
        );

    \I__8356\ : InMux
    port map (
            O => \N__36082\,
            I => \N__36043\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__36077\,
            I => \N__36040\
        );

    \I__8354\ : CascadeMux
    port map (
            O => \N__36076\,
            I => \N__36033\
        );

    \I__8353\ : Span4Mux_v
    port map (
            O => \N__36067\,
            I => \N__36018\
        );

    \I__8352\ : Span4Mux_v
    port map (
            O => \N__36062\,
            I => \N__36018\
        );

    \I__8351\ : LocalMux
    port map (
            O => \N__36057\,
            I => \N__36009\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__36050\,
            I => \N__36009\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__36043\,
            I => \N__36009\
        );

    \I__8348\ : Sp12to4
    port map (
            O => \N__36040\,
            I => \N__36009\
        );

    \I__8347\ : InMux
    port map (
            O => \N__36039\,
            I => \N__36004\
        );

    \I__8346\ : InMux
    port map (
            O => \N__36038\,
            I => \N__36004\
        );

    \I__8345\ : InMux
    port map (
            O => \N__36037\,
            I => \N__36001\
        );

    \I__8344\ : SRMux
    port map (
            O => \N__36036\,
            I => \N__35996\
        );

    \I__8343\ : InMux
    port map (
            O => \N__36033\,
            I => \N__35996\
        );

    \I__8342\ : InMux
    port map (
            O => \N__36032\,
            I => \N__35991\
        );

    \I__8341\ : InMux
    port map (
            O => \N__36031\,
            I => \N__35991\
        );

    \I__8340\ : InMux
    port map (
            O => \N__36030\,
            I => \N__35984\
        );

    \I__8339\ : InMux
    port map (
            O => \N__36029\,
            I => \N__35984\
        );

    \I__8338\ : InMux
    port map (
            O => \N__36028\,
            I => \N__35984\
        );

    \I__8337\ : InMux
    port map (
            O => \N__36027\,
            I => \N__35975\
        );

    \I__8336\ : InMux
    port map (
            O => \N__36026\,
            I => \N__35975\
        );

    \I__8335\ : InMux
    port map (
            O => \N__36025\,
            I => \N__35975\
        );

    \I__8334\ : InMux
    port map (
            O => \N__36024\,
            I => \N__35975\
        );

    \I__8333\ : InMux
    port map (
            O => \N__36023\,
            I => \N__35972\
        );

    \I__8332\ : Span4Mux_v
    port map (
            O => \N__36018\,
            I => \N__35969\
        );

    \I__8331\ : Span12Mux_s10_v
    port map (
            O => \N__36009\,
            I => \N__35966\
        );

    \I__8330\ : LocalMux
    port map (
            O => \N__36004\,
            I => \N__35951\
        );

    \I__8329\ : LocalMux
    port map (
            O => \N__36001\,
            I => \N__35951\
        );

    \I__8328\ : LocalMux
    port map (
            O => \N__35996\,
            I => \N__35951\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__35991\,
            I => \N__35951\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__35984\,
            I => \N__35951\
        );

    \I__8325\ : LocalMux
    port map (
            O => \N__35975\,
            I => \N__35951\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__35972\,
            I => \N__35951\
        );

    \I__8323\ : Odrv4
    port map (
            O => \N__35969\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8322\ : Odrv12
    port map (
            O => \N__35966\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8321\ : Odrv12
    port map (
            O => \N__35951\,
            I => \b2v_inst6.count_0_sqmuxa\
        );

    \I__8320\ : InMux
    port map (
            O => \N__35944\,
            I => \N__35941\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__35941\,
            I => \b2v_inst6.curr_state_1_0\
        );

    \I__8318\ : CascadeMux
    port map (
            O => \N__35938\,
            I => \N__35935\
        );

    \I__8317\ : InMux
    port map (
            O => \N__35935\,
            I => \N__35926\
        );

    \I__8316\ : CascadeMux
    port map (
            O => \N__35934\,
            I => \N__35919\
        );

    \I__8315\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35910\
        );

    \I__8314\ : InMux
    port map (
            O => \N__35932\,
            I => \N__35910\
        );

    \I__8313\ : InMux
    port map (
            O => \N__35931\,
            I => \N__35905\
        );

    \I__8312\ : InMux
    port map (
            O => \N__35930\,
            I => \N__35905\
        );

    \I__8311\ : CascadeMux
    port map (
            O => \N__35929\,
            I => \N__35893\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__35926\,
            I => \N__35888\
        );

    \I__8309\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35880\
        );

    \I__8308\ : InMux
    port map (
            O => \N__35924\,
            I => \N__35880\
        );

    \I__8307\ : InMux
    port map (
            O => \N__35923\,
            I => \N__35871\
        );

    \I__8306\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35871\
        );

    \I__8305\ : InMux
    port map (
            O => \N__35919\,
            I => \N__35871\
        );

    \I__8304\ : InMux
    port map (
            O => \N__35918\,
            I => \N__35871\
        );

    \I__8303\ : InMux
    port map (
            O => \N__35917\,
            I => \N__35867\
        );

    \I__8302\ : InMux
    port map (
            O => \N__35916\,
            I => \N__35862\
        );

    \I__8301\ : InMux
    port map (
            O => \N__35915\,
            I => \N__35862\
        );

    \I__8300\ : LocalMux
    port map (
            O => \N__35910\,
            I => \N__35854\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__35905\,
            I => \N__35854\
        );

    \I__8298\ : InMux
    port map (
            O => \N__35904\,
            I => \N__35847\
        );

    \I__8297\ : InMux
    port map (
            O => \N__35903\,
            I => \N__35847\
        );

    \I__8296\ : InMux
    port map (
            O => \N__35902\,
            I => \N__35847\
        );

    \I__8295\ : InMux
    port map (
            O => \N__35901\,
            I => \N__35844\
        );

    \I__8294\ : InMux
    port map (
            O => \N__35900\,
            I => \N__35837\
        );

    \I__8293\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35837\
        );

    \I__8292\ : InMux
    port map (
            O => \N__35898\,
            I => \N__35837\
        );

    \I__8291\ : InMux
    port map (
            O => \N__35897\,
            I => \N__35834\
        );

    \I__8290\ : InMux
    port map (
            O => \N__35896\,
            I => \N__35831\
        );

    \I__8289\ : InMux
    port map (
            O => \N__35893\,
            I => \N__35828\
        );

    \I__8288\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35821\
        );

    \I__8287\ : InMux
    port map (
            O => \N__35891\,
            I => \N__35821\
        );

    \I__8286\ : Span4Mux_v
    port map (
            O => \N__35888\,
            I => \N__35816\
        );

    \I__8285\ : InMux
    port map (
            O => \N__35887\,
            I => \N__35807\
        );

    \I__8284\ : InMux
    port map (
            O => \N__35886\,
            I => \N__35802\
        );

    \I__8283\ : InMux
    port map (
            O => \N__35885\,
            I => \N__35802\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__35880\,
            I => \N__35797\
        );

    \I__8281\ : LocalMux
    port map (
            O => \N__35871\,
            I => \N__35797\
        );

    \I__8280\ : InMux
    port map (
            O => \N__35870\,
            I => \N__35794\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__35867\,
            I => \N__35789\
        );

    \I__8278\ : LocalMux
    port map (
            O => \N__35862\,
            I => \N__35789\
        );

    \I__8277\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35782\
        );

    \I__8276\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35782\
        );

    \I__8275\ : InMux
    port map (
            O => \N__35859\,
            I => \N__35782\
        );

    \I__8274\ : Span12Mux_s9_h
    port map (
            O => \N__35854\,
            I => \N__35779\
        );

    \I__8273\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35776\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__35844\,
            I => \N__35769\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__35837\,
            I => \N__35769\
        );

    \I__8270\ : LocalMux
    port map (
            O => \N__35834\,
            I => \N__35764\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__35831\,
            I => \N__35764\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__35828\,
            I => \N__35761\
        );

    \I__8267\ : InMux
    port map (
            O => \N__35827\,
            I => \N__35758\
        );

    \I__8266\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35755\
        );

    \I__8265\ : LocalMux
    port map (
            O => \N__35821\,
            I => \N__35752\
        );

    \I__8264\ : InMux
    port map (
            O => \N__35820\,
            I => \N__35749\
        );

    \I__8263\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35746\
        );

    \I__8262\ : Span4Mux_v
    port map (
            O => \N__35816\,
            I => \N__35741\
        );

    \I__8261\ : InMux
    port map (
            O => \N__35815\,
            I => \N__35736\
        );

    \I__8260\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35736\
        );

    \I__8259\ : InMux
    port map (
            O => \N__35813\,
            I => \N__35731\
        );

    \I__8258\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35731\
        );

    \I__8257\ : InMux
    port map (
            O => \N__35811\,
            I => \N__35726\
        );

    \I__8256\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35726\
        );

    \I__8255\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35715\
        );

    \I__8254\ : LocalMux
    port map (
            O => \N__35802\,
            I => \N__35715\
        );

    \I__8253\ : Span4Mux_v
    port map (
            O => \N__35797\,
            I => \N__35715\
        );

    \I__8252\ : LocalMux
    port map (
            O => \N__35794\,
            I => \N__35715\
        );

    \I__8251\ : Span4Mux_s1_v
    port map (
            O => \N__35789\,
            I => \N__35715\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__35782\,
            I => \N__35710\
        );

    \I__8249\ : Span12Mux_v
    port map (
            O => \N__35779\,
            I => \N__35710\
        );

    \I__8248\ : Span12Mux_s4_h
    port map (
            O => \N__35776\,
            I => \N__35707\
        );

    \I__8247\ : InMux
    port map (
            O => \N__35775\,
            I => \N__35702\
        );

    \I__8246\ : InMux
    port map (
            O => \N__35774\,
            I => \N__35702\
        );

    \I__8245\ : Span12Mux_s7_h
    port map (
            O => \N__35769\,
            I => \N__35699\
        );

    \I__8244\ : Span4Mux_v
    port map (
            O => \N__35764\,
            I => \N__35684\
        );

    \I__8243\ : Span4Mux_h
    port map (
            O => \N__35761\,
            I => \N__35684\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__35758\,
            I => \N__35684\
        );

    \I__8241\ : LocalMux
    port map (
            O => \N__35755\,
            I => \N__35684\
        );

    \I__8240\ : Span4Mux_h
    port map (
            O => \N__35752\,
            I => \N__35684\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__35749\,
            I => \N__35684\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__35746\,
            I => \N__35684\
        );

    \I__8237\ : InMux
    port map (
            O => \N__35745\,
            I => \N__35679\
        );

    \I__8236\ : InMux
    port map (
            O => \N__35744\,
            I => \N__35679\
        );

    \I__8235\ : Odrv4
    port map (
            O => \N__35741\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8234\ : LocalMux
    port map (
            O => \N__35736\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__35731\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8232\ : LocalMux
    port map (
            O => \N__35726\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__35715\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8230\ : Odrv12
    port map (
            O => \N__35710\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8229\ : Odrv12
    port map (
            O => \N__35707\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__35702\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8227\ : Odrv12
    port map (
            O => \N__35699\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8226\ : Odrv4
    port map (
            O => \N__35684\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__35679\,
            I => \SYNTHESIZED_WIRE_1keep_3\
        );

    \I__8224\ : InMux
    port map (
            O => \N__35656\,
            I => \N__35647\
        );

    \I__8223\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35647\
        );

    \I__8222\ : InMux
    port map (
            O => \N__35654\,
            I => \N__35640\
        );

    \I__8221\ : InMux
    port map (
            O => \N__35653\,
            I => \N__35640\
        );

    \I__8220\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35640\
        );

    \I__8219\ : LocalMux
    port map (
            O => \N__35647\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__35640\,
            I => \b2v_inst6.curr_stateZ0Z_0\
        );

    \I__8217\ : CascadeMux
    port map (
            O => \N__35635\,
            I => \b2v_inst6.curr_stateZ0Z_1_cascade_\
        );

    \I__8216\ : InMux
    port map (
            O => \N__35632\,
            I => \N__35627\
        );

    \I__8215\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35622\
        );

    \I__8214\ : InMux
    port map (
            O => \N__35630\,
            I => \N__35622\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__35627\,
            I => \b2v_inst6.curr_state_RNIUL1J2Z0Z_0\
        );

    \I__8212\ : LocalMux
    port map (
            O => \N__35622\,
            I => \b2v_inst6.curr_state_RNIUL1J2Z0Z_0\
        );

    \I__8211\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35614\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__35614\,
            I => \b2v_inst6.curr_state_7_0\
        );

    \I__8209\ : InMux
    port map (
            O => \N__35611\,
            I => \b2v_inst11.mult1_un75_sum_cry_5\
        );

    \I__8208\ : CascadeMux
    port map (
            O => \N__35608\,
            I => \N__35604\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__35607\,
            I => \N__35600\
        );

    \I__8206\ : InMux
    port map (
            O => \N__35604\,
            I => \N__35593\
        );

    \I__8205\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35593\
        );

    \I__8204\ : InMux
    port map (
            O => \N__35600\,
            I => \N__35593\
        );

    \I__8203\ : LocalMux
    port map (
            O => \N__35593\,
            I => \b2v_inst11.mult1_un68_sum_i_0_8\
        );

    \I__8202\ : CascadeMux
    port map (
            O => \N__35590\,
            I => \N__35587\
        );

    \I__8201\ : InMux
    port map (
            O => \N__35587\,
            I => \N__35584\
        );

    \I__8200\ : LocalMux
    port map (
            O => \N__35584\,
            I => \b2v_inst11.mult1_un82_sum_axb_8\
        );

    \I__8199\ : InMux
    port map (
            O => \N__35581\,
            I => \b2v_inst11.mult1_un75_sum_cry_6\
        );

    \I__8198\ : InMux
    port map (
            O => \N__35578\,
            I => \b2v_inst11.mult1_un75_sum_cry_7\
        );

    \I__8197\ : InMux
    port map (
            O => \N__35575\,
            I => \N__35571\
        );

    \I__8196\ : CascadeMux
    port map (
            O => \N__35574\,
            I => \N__35567\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__35571\,
            I => \N__35563\
        );

    \I__8194\ : InMux
    port map (
            O => \N__35570\,
            I => \N__35558\
        );

    \I__8193\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35558\
        );

    \I__8192\ : InMux
    port map (
            O => \N__35566\,
            I => \N__35555\
        );

    \I__8191\ : Odrv12
    port map (
            O => \N__35563\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__35558\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__35555\,
            I => \b2v_inst11.mult1_un75_sum_s_8\
        );

    \I__8188\ : CascadeMux
    port map (
            O => \N__35548\,
            I => \b2v_inst11.mult1_un75_sum_s_8_cascade_\
        );

    \I__8187\ : CascadeMux
    port map (
            O => \N__35545\,
            I => \N__35541\
        );

    \I__8186\ : CascadeMux
    port map (
            O => \N__35544\,
            I => \N__35537\
        );

    \I__8185\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35530\
        );

    \I__8184\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35530\
        );

    \I__8183\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35530\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__35530\,
            I => \b2v_inst11.mult1_un75_sum_i_0_8\
        );

    \I__8181\ : InMux
    port map (
            O => \N__35527\,
            I => \N__35523\
        );

    \I__8180\ : InMux
    port map (
            O => \N__35526\,
            I => \N__35520\
        );

    \I__8179\ : LocalMux
    port map (
            O => \N__35523\,
            I => \N__35517\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__35520\,
            I => \N__35514\
        );

    \I__8177\ : Span4Mux_v
    port map (
            O => \N__35517\,
            I => \N__35511\
        );

    \I__8176\ : Span4Mux_s2_h
    port map (
            O => \N__35514\,
            I => \N__35508\
        );

    \I__8175\ : Odrv4
    port map (
            O => \N__35511\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__8174\ : Odrv4
    port map (
            O => \N__35508\,
            I => \b2v_inst11.mult1_un68_sum\
        );

    \I__8173\ : InMux
    port map (
            O => \N__35503\,
            I => \N__35500\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__35500\,
            I => \b2v_inst11.mult1_un61_sum_i\
        );

    \I__8171\ : CascadeMux
    port map (
            O => \N__35497\,
            I => \N__35494\
        );

    \I__8170\ : InMux
    port map (
            O => \N__35494\,
            I => \N__35491\
        );

    \I__8169\ : LocalMux
    port map (
            O => \N__35491\,
            I => \b2v_inst11.mult1_un68_sum_cry_3_s\
        );

    \I__8168\ : InMux
    port map (
            O => \N__35488\,
            I => \b2v_inst11.mult1_un68_sum_cry_2\
        );

    \I__8167\ : CascadeMux
    port map (
            O => \N__35485\,
            I => \N__35482\
        );

    \I__8166\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35479\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__35479\,
            I => \b2v_inst11.mult1_un61_sum_cry_3_s\
        );

    \I__8164\ : InMux
    port map (
            O => \N__35476\,
            I => \N__35473\
        );

    \I__8163\ : LocalMux
    port map (
            O => \N__35473\,
            I => \b2v_inst11.mult1_un68_sum_cry_4_s\
        );

    \I__8162\ : InMux
    port map (
            O => \N__35470\,
            I => \b2v_inst11.mult1_un68_sum_cry_3\
        );

    \I__8161\ : InMux
    port map (
            O => \N__35467\,
            I => \N__35464\
        );

    \I__8160\ : LocalMux
    port map (
            O => \N__35464\,
            I => \b2v_inst11.mult1_un61_sum_cry_4_s\
        );

    \I__8159\ : CascadeMux
    port map (
            O => \N__35461\,
            I => \N__35458\
        );

    \I__8158\ : InMux
    port map (
            O => \N__35458\,
            I => \N__35455\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__35455\,
            I => \b2v_inst11.mult1_un68_sum_cry_5_s\
        );

    \I__8156\ : InMux
    port map (
            O => \N__35452\,
            I => \b2v_inst11.mult1_un68_sum_cry_4\
        );

    \I__8155\ : CascadeMux
    port map (
            O => \N__35449\,
            I => \N__35444\
        );

    \I__8154\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35440\
        );

    \I__8153\ : InMux
    port map (
            O => \N__35447\,
            I => \N__35435\
        );

    \I__8152\ : InMux
    port map (
            O => \N__35444\,
            I => \N__35435\
        );

    \I__8151\ : InMux
    port map (
            O => \N__35443\,
            I => \N__35432\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__35440\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__8149\ : LocalMux
    port map (
            O => \N__35435\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__8148\ : LocalMux
    port map (
            O => \N__35432\,
            I => \b2v_inst11.mult1_un61_sum_s_8\
        );

    \I__8147\ : CascadeMux
    port map (
            O => \N__35425\,
            I => \N__35422\
        );

    \I__8146\ : InMux
    port map (
            O => \N__35422\,
            I => \N__35419\
        );

    \I__8145\ : LocalMux
    port map (
            O => \N__35419\,
            I => \b2v_inst11.mult1_un61_sum_cry_5_s\
        );

    \I__8144\ : InMux
    port map (
            O => \N__35416\,
            I => \N__35413\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__35413\,
            I => \b2v_inst11.mult1_un68_sum_cry_6_s\
        );

    \I__8142\ : InMux
    port map (
            O => \N__35410\,
            I => \N__35407\
        );

    \I__8141\ : LocalMux
    port map (
            O => \N__35407\,
            I => \N__35404\
        );

    \I__8140\ : Odrv4
    port map (
            O => \N__35404\,
            I => \b2v_inst11.mult1_un82_sum_cry_6_s\
        );

    \I__8139\ : InMux
    port map (
            O => \N__35401\,
            I => \b2v_inst11.mult1_un82_sum_cry_5\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__35398\,
            I => \N__35395\
        );

    \I__8137\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35392\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__35392\,
            I => \b2v_inst11.mult1_un89_sum_axb_8\
        );

    \I__8135\ : InMux
    port map (
            O => \N__35389\,
            I => \b2v_inst11.mult1_un82_sum_cry_6\
        );

    \I__8134\ : InMux
    port map (
            O => \N__35386\,
            I => \b2v_inst11.mult1_un82_sum_cry_7\
        );

    \I__8133\ : CascadeMux
    port map (
            O => \N__35383\,
            I => \N__35378\
        );

    \I__8132\ : InMux
    port map (
            O => \N__35382\,
            I => \N__35374\
        );

    \I__8131\ : InMux
    port map (
            O => \N__35381\,
            I => \N__35369\
        );

    \I__8130\ : InMux
    port map (
            O => \N__35378\,
            I => \N__35369\
        );

    \I__8129\ : InMux
    port map (
            O => \N__35377\,
            I => \N__35366\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__35374\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__35369\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__35366\,
            I => \b2v_inst11.mult1_un82_sum_s_8\
        );

    \I__8125\ : CascadeMux
    port map (
            O => \N__35359\,
            I => \b2v_inst11.mult1_un82_sum_s_8_cascade_\
        );

    \I__8124\ : CascadeMux
    port map (
            O => \N__35356\,
            I => \N__35352\
        );

    \I__8123\ : CascadeMux
    port map (
            O => \N__35355\,
            I => \N__35348\
        );

    \I__8122\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35341\
        );

    \I__8121\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35341\
        );

    \I__8120\ : InMux
    port map (
            O => \N__35348\,
            I => \N__35341\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__35341\,
            I => \b2v_inst11.mult1_un82_sum_i_0_8\
        );

    \I__8118\ : InMux
    port map (
            O => \N__35338\,
            I => \N__35334\
        );

    \I__8117\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35331\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__35334\,
            I => \N__35328\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__35331\,
            I => \N__35323\
        );

    \I__8114\ : Span4Mux_v
    port map (
            O => \N__35328\,
            I => \N__35323\
        );

    \I__8113\ : Odrv4
    port map (
            O => \N__35323\,
            I => \b2v_inst11.mult1_un75_sum\
        );

    \I__8112\ : InMux
    port map (
            O => \N__35320\,
            I => \N__35317\
        );

    \I__8111\ : LocalMux
    port map (
            O => \N__35317\,
            I => \b2v_inst11.mult1_un68_sum_i\
        );

    \I__8110\ : CascadeMux
    port map (
            O => \N__35314\,
            I => \N__35311\
        );

    \I__8109\ : InMux
    port map (
            O => \N__35311\,
            I => \N__35308\
        );

    \I__8108\ : LocalMux
    port map (
            O => \N__35308\,
            I => \b2v_inst11.mult1_un75_sum_cry_3_s\
        );

    \I__8107\ : InMux
    port map (
            O => \N__35305\,
            I => \b2v_inst11.mult1_un75_sum_cry_2\
        );

    \I__8106\ : InMux
    port map (
            O => \N__35302\,
            I => \N__35299\
        );

    \I__8105\ : LocalMux
    port map (
            O => \N__35299\,
            I => \b2v_inst11.mult1_un75_sum_cry_4_s\
        );

    \I__8104\ : InMux
    port map (
            O => \N__35296\,
            I => \b2v_inst11.mult1_un75_sum_cry_3\
        );

    \I__8103\ : CascadeMux
    port map (
            O => \N__35293\,
            I => \N__35290\
        );

    \I__8102\ : InMux
    port map (
            O => \N__35290\,
            I => \N__35287\
        );

    \I__8101\ : LocalMux
    port map (
            O => \N__35287\,
            I => \b2v_inst11.mult1_un75_sum_cry_5_s\
        );

    \I__8100\ : InMux
    port map (
            O => \N__35284\,
            I => \b2v_inst11.mult1_un75_sum_cry_4\
        );

    \I__8099\ : InMux
    port map (
            O => \N__35281\,
            I => \N__35278\
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__35278\,
            I => \b2v_inst11.mult1_un75_sum_cry_6_s\
        );

    \I__8097\ : InMux
    port map (
            O => \N__35275\,
            I => \N__35272\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__35272\,
            I => \b2v_inst11.mult1_un89_sum_cry_5_s\
        );

    \I__8095\ : InMux
    port map (
            O => \N__35269\,
            I => \N__35266\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__35266\,
            I => \N__35263\
        );

    \I__8093\ : Span4Mux_h
    port map (
            O => \N__35263\,
            I => \N__35260\
        );

    \I__8092\ : Odrv4
    port map (
            O => \N__35260\,
            I => \b2v_inst11.mult1_un96_sum_cry_6_s\
        );

    \I__8091\ : InMux
    port map (
            O => \N__35257\,
            I => \b2v_inst11.mult1_un96_sum_cry_5\
        );

    \I__8090\ : InMux
    port map (
            O => \N__35254\,
            I => \N__35251\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__35251\,
            I => \b2v_inst11.mult1_un89_sum_cry_6_s\
        );

    \I__8088\ : CascadeMux
    port map (
            O => \N__35248\,
            I => \N__35245\
        );

    \I__8087\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35242\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__35242\,
            I => \N__35239\
        );

    \I__8085\ : Span4Mux_h
    port map (
            O => \N__35239\,
            I => \N__35236\
        );

    \I__8084\ : Odrv4
    port map (
            O => \N__35236\,
            I => \b2v_inst11.mult1_un103_sum_axb_8\
        );

    \I__8083\ : InMux
    port map (
            O => \N__35233\,
            I => \b2v_inst11.mult1_un96_sum_cry_6\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__35230\,
            I => \N__35227\
        );

    \I__8081\ : InMux
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__35224\,
            I => \b2v_inst11.mult1_un96_sum_axb_8\
        );

    \I__8079\ : InMux
    port map (
            O => \N__35221\,
            I => \b2v_inst11.mult1_un96_sum_cry_7\
        );

    \I__8078\ : CascadeMux
    port map (
            O => \N__35218\,
            I => \N__35214\
        );

    \I__8077\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35208\
        );

    \I__8076\ : InMux
    port map (
            O => \N__35214\,
            I => \N__35208\
        );

    \I__8075\ : InMux
    port map (
            O => \N__35213\,
            I => \N__35205\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__35208\,
            I => \N__35198\
        );

    \I__8073\ : LocalMux
    port map (
            O => \N__35205\,
            I => \N__35198\
        );

    \I__8072\ : InMux
    port map (
            O => \N__35204\,
            I => \N__35195\
        );

    \I__8071\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35192\
        );

    \I__8070\ : Span4Mux_h
    port map (
            O => \N__35198\,
            I => \N__35189\
        );

    \I__8069\ : LocalMux
    port map (
            O => \N__35195\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__8068\ : LocalMux
    port map (
            O => \N__35192\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__8067\ : Odrv4
    port map (
            O => \N__35189\,
            I => \b2v_inst11.mult1_un96_sum_s_8\
        );

    \I__8066\ : CascadeMux
    port map (
            O => \N__35182\,
            I => \N__35177\
        );

    \I__8065\ : InMux
    port map (
            O => \N__35181\,
            I => \N__35172\
        );

    \I__8064\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35169\
        );

    \I__8063\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35162\
        );

    \I__8062\ : InMux
    port map (
            O => \N__35176\,
            I => \N__35162\
        );

    \I__8061\ : InMux
    port map (
            O => \N__35175\,
            I => \N__35162\
        );

    \I__8060\ : LocalMux
    port map (
            O => \N__35172\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__35169\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__35162\,
            I => \b2v_inst11.mult1_un89_sum_s_8\
        );

    \I__8057\ : CascadeMux
    port map (
            O => \N__35155\,
            I => \N__35151\
        );

    \I__8056\ : CascadeMux
    port map (
            O => \N__35154\,
            I => \N__35147\
        );

    \I__8055\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35140\
        );

    \I__8054\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35140\
        );

    \I__8053\ : InMux
    port map (
            O => \N__35147\,
            I => \N__35140\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__35140\,
            I => \b2v_inst11.mult1_un89_sum_i_0_8\
        );

    \I__8051\ : InMux
    port map (
            O => \N__35137\,
            I => \N__35133\
        );

    \I__8050\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35130\
        );

    \I__8049\ : LocalMux
    port map (
            O => \N__35133\,
            I => \N__35127\
        );

    \I__8048\ : LocalMux
    port map (
            O => \N__35130\,
            I => \N__35124\
        );

    \I__8047\ : Span4Mux_s3_h
    port map (
            O => \N__35127\,
            I => \N__35121\
        );

    \I__8046\ : Odrv4
    port map (
            O => \N__35124\,
            I => \b2v_inst11.mult1_un82_sum\
        );

    \I__8045\ : Odrv4
    port map (
            O => \N__35121\,
            I => \b2v_inst11.mult1_un82_sum\
        );

    \I__8044\ : InMux
    port map (
            O => \N__35116\,
            I => \N__35113\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__35113\,
            I => \b2v_inst11.mult1_un75_sum_i\
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__35110\,
            I => \N__35107\
        );

    \I__8041\ : InMux
    port map (
            O => \N__35107\,
            I => \N__35104\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__35104\,
            I => \b2v_inst11.mult1_un82_sum_cry_3_s\
        );

    \I__8039\ : InMux
    port map (
            O => \N__35101\,
            I => \b2v_inst11.mult1_un82_sum_cry_2\
        );

    \I__8038\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35095\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__35095\,
            I => \b2v_inst11.mult1_un82_sum_cry_4_s\
        );

    \I__8036\ : InMux
    port map (
            O => \N__35092\,
            I => \b2v_inst11.mult1_un82_sum_cry_3\
        );

    \I__8035\ : CascadeMux
    port map (
            O => \N__35089\,
            I => \N__35086\
        );

    \I__8034\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35083\
        );

    \I__8033\ : LocalMux
    port map (
            O => \N__35083\,
            I => \b2v_inst11.mult1_un82_sum_cry_5_s\
        );

    \I__8032\ : InMux
    port map (
            O => \N__35080\,
            I => \b2v_inst11.mult1_un82_sum_cry_4\
        );

    \I__8031\ : InMux
    port map (
            O => \N__35077\,
            I => \N__35074\
        );

    \I__8030\ : LocalMux
    port map (
            O => \N__35074\,
            I => \N__35071\
        );

    \I__8029\ : Span4Mux_h
    port map (
            O => \N__35071\,
            I => \N__35068\
        );

    \I__8028\ : Odrv4
    port map (
            O => \N__35068\,
            I => \b2v_inst11.mult1_un96_sum_i\
        );

    \I__8027\ : InMux
    port map (
            O => \N__35065\,
            I => \N__35062\
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__35062\,
            I => \b2v_inst11.mult1_un68_sum_i_8\
        );

    \I__8025\ : CEMux
    port map (
            O => \N__35059\,
            I => \N__35054\
        );

    \I__8024\ : CEMux
    port map (
            O => \N__35058\,
            I => \N__35050\
        );

    \I__8023\ : CascadeMux
    port map (
            O => \N__35057\,
            I => \N__35047\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__35054\,
            I => \N__35035\
        );

    \I__8021\ : CEMux
    port map (
            O => \N__35053\,
            I => \N__35032\
        );

    \I__8020\ : LocalMux
    port map (
            O => \N__35050\,
            I => \N__35029\
        );

    \I__8019\ : InMux
    port map (
            O => \N__35047\,
            I => \N__35024\
        );

    \I__8018\ : CEMux
    port map (
            O => \N__35046\,
            I => \N__35024\
        );

    \I__8017\ : InMux
    port map (
            O => \N__35045\,
            I => \N__35011\
        );

    \I__8016\ : CEMux
    port map (
            O => \N__35044\,
            I => \N__35011\
        );

    \I__8015\ : InMux
    port map (
            O => \N__35043\,
            I => \N__35008\
        );

    \I__8014\ : InMux
    port map (
            O => \N__35042\,
            I => \N__35003\
        );

    \I__8013\ : InMux
    port map (
            O => \N__35041\,
            I => \N__35003\
        );

    \I__8012\ : InMux
    port map (
            O => \N__35040\,
            I => \N__34996\
        );

    \I__8011\ : InMux
    port map (
            O => \N__35039\,
            I => \N__34996\
        );

    \I__8010\ : InMux
    port map (
            O => \N__35038\,
            I => \N__34996\
        );

    \I__8009\ : Span4Mux_s2_v
    port map (
            O => \N__35035\,
            I => \N__34990\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__35032\,
            I => \N__34990\
        );

    \I__8007\ : Span4Mux_s3_v
    port map (
            O => \N__35029\,
            I => \N__34987\
        );

    \I__8006\ : LocalMux
    port map (
            O => \N__35024\,
            I => \N__34984\
        );

    \I__8005\ : InMux
    port map (
            O => \N__35023\,
            I => \N__34981\
        );

    \I__8004\ : InMux
    port map (
            O => \N__35022\,
            I => \N__34978\
        );

    \I__8003\ : InMux
    port map (
            O => \N__35021\,
            I => \N__34971\
        );

    \I__8002\ : InMux
    port map (
            O => \N__35020\,
            I => \N__34971\
        );

    \I__8001\ : InMux
    port map (
            O => \N__35019\,
            I => \N__34971\
        );

    \I__8000\ : CEMux
    port map (
            O => \N__35018\,
            I => \N__34964\
        );

    \I__7999\ : InMux
    port map (
            O => \N__35017\,
            I => \N__34964\
        );

    \I__7998\ : InMux
    port map (
            O => \N__35016\,
            I => \N__34964\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__35011\,
            I => \N__34955\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__35008\,
            I => \N__34955\
        );

    \I__7995\ : LocalMux
    port map (
            O => \N__35003\,
            I => \N__34955\
        );

    \I__7994\ : LocalMux
    port map (
            O => \N__34996\,
            I => \N__34955\
        );

    \I__7993\ : CascadeMux
    port map (
            O => \N__34995\,
            I => \N__34952\
        );

    \I__7992\ : Span4Mux_v
    port map (
            O => \N__34990\,
            I => \N__34949\
        );

    \I__7991\ : Span4Mux_v
    port map (
            O => \N__34987\,
            I => \N__34944\
        );

    \I__7990\ : Span4Mux_s0_h
    port map (
            O => \N__34984\,
            I => \N__34944\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__34981\,
            I => \N__34933\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__34978\,
            I => \N__34933\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__34971\,
            I => \N__34933\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__34964\,
            I => \N__34933\
        );

    \I__7985\ : Sp12to4
    port map (
            O => \N__34955\,
            I => \N__34933\
        );

    \I__7984\ : InMux
    port map (
            O => \N__34952\,
            I => \N__34930\
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__34949\,
            I => \b2v_inst6.count_en\
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__34944\,
            I => \b2v_inst6.count_en\
        );

    \I__7981\ : Odrv12
    port map (
            O => \N__34933\,
            I => \b2v_inst6.count_en\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__34930\,
            I => \b2v_inst6.count_en\
        );

    \I__7979\ : InMux
    port map (
            O => \N__34921\,
            I => \N__34918\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__34918\,
            I => \N__34915\
        );

    \I__7977\ : Span4Mux_v
    port map (
            O => \N__34915\,
            I => \N__34912\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__34912\,
            I => \b2v_inst6.count_RNIM2CM2Z0Z_0\
        );

    \I__7975\ : CascadeMux
    port map (
            O => \N__34909\,
            I => \b2v_inst6.count_en_cascade_\
        );

    \I__7974\ : InMux
    port map (
            O => \N__34906\,
            I => \N__34903\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__34903\,
            I => \b2v_inst6.count_0_0\
        );

    \I__7972\ : InMux
    port map (
            O => \N__34900\,
            I => \N__34896\
        );

    \I__7971\ : CascadeMux
    port map (
            O => \N__34899\,
            I => \N__34893\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__34896\,
            I => \N__34889\
        );

    \I__7969\ : InMux
    port map (
            O => \N__34893\,
            I => \N__34884\
        );

    \I__7968\ : InMux
    port map (
            O => \N__34892\,
            I => \N__34884\
        );

    \I__7967\ : Span12Mux_s3_v
    port map (
            O => \N__34889\,
            I => \N__34879\
        );

    \I__7966\ : LocalMux
    port map (
            O => \N__34884\,
            I => \N__34876\
        );

    \I__7965\ : InMux
    port map (
            O => \N__34883\,
            I => \N__34871\
        );

    \I__7964\ : InMux
    port map (
            O => \N__34882\,
            I => \N__34871\
        );

    \I__7963\ : Odrv12
    port map (
            O => \N__34879\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7962\ : Odrv4
    port map (
            O => \N__34876\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__34871\,
            I => \b2v_inst6.countZ0Z_0\
        );

    \I__7960\ : InMux
    port map (
            O => \N__34864\,
            I => \N__34860\
        );

    \I__7959\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34857\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__34860\,
            I => \N__34854\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__34857\,
            I => \N__34851\
        );

    \I__7956\ : Span4Mux_s2_h
    port map (
            O => \N__34854\,
            I => \N__34848\
        );

    \I__7955\ : Odrv12
    port map (
            O => \N__34851\,
            I => \b2v_inst11.mult1_un96_sum\
        );

    \I__7954\ : Odrv4
    port map (
            O => \N__34848\,
            I => \b2v_inst11.mult1_un96_sum\
        );

    \I__7953\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34840\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__34840\,
            I => \b2v_inst11.mult1_un89_sum_i\
        );

    \I__7951\ : CascadeMux
    port map (
            O => \N__34837\,
            I => \N__34834\
        );

    \I__7950\ : InMux
    port map (
            O => \N__34834\,
            I => \N__34831\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__34831\,
            I => \N__34828\
        );

    \I__7948\ : Span4Mux_h
    port map (
            O => \N__34828\,
            I => \N__34825\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__34825\,
            I => \b2v_inst11.mult1_un96_sum_cry_3_s\
        );

    \I__7946\ : InMux
    port map (
            O => \N__34822\,
            I => \b2v_inst11.mult1_un96_sum_cry_2\
        );

    \I__7945\ : CascadeMux
    port map (
            O => \N__34819\,
            I => \N__34816\
        );

    \I__7944\ : InMux
    port map (
            O => \N__34816\,
            I => \N__34813\
        );

    \I__7943\ : LocalMux
    port map (
            O => \N__34813\,
            I => \b2v_inst11.mult1_un89_sum_cry_3_s\
        );

    \I__7942\ : InMux
    port map (
            O => \N__34810\,
            I => \N__34807\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__34807\,
            I => \N__34804\
        );

    \I__7940\ : Span4Mux_v
    port map (
            O => \N__34804\,
            I => \N__34801\
        );

    \I__7939\ : Odrv4
    port map (
            O => \N__34801\,
            I => \b2v_inst11.mult1_un96_sum_cry_4_s\
        );

    \I__7938\ : InMux
    port map (
            O => \N__34798\,
            I => \b2v_inst11.mult1_un96_sum_cry_3\
        );

    \I__7937\ : CascadeMux
    port map (
            O => \N__34795\,
            I => \N__34792\
        );

    \I__7936\ : InMux
    port map (
            O => \N__34792\,
            I => \N__34789\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__34789\,
            I => \b2v_inst11.mult1_un89_sum_cry_4_s\
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__34786\,
            I => \N__34783\
        );

    \I__7933\ : InMux
    port map (
            O => \N__34783\,
            I => \N__34780\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__34780\,
            I => \N__34777\
        );

    \I__7931\ : Span4Mux_v
    port map (
            O => \N__34777\,
            I => \N__34774\
        );

    \I__7930\ : Odrv4
    port map (
            O => \N__34774\,
            I => \b2v_inst11.mult1_un96_sum_cry_5_s\
        );

    \I__7929\ : InMux
    port map (
            O => \N__34771\,
            I => \b2v_inst11.mult1_un96_sum_cry_4\
        );

    \I__7928\ : CascadeMux
    port map (
            O => \N__34768\,
            I => \b2v_inst6.un2_count_1_axb_1_cascade_\
        );

    \I__7927\ : InMux
    port map (
            O => \N__34765\,
            I => \N__34762\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34759\
        );

    \I__7925\ : IoSpan4Mux
    port map (
            O => \N__34759\,
            I => \N__34756\
        );

    \I__7924\ : Odrv4
    port map (
            O => \N__34756\,
            I => \V1P8A_OK_c\
        );

    \I__7923\ : InMux
    port map (
            O => \N__34753\,
            I => \N__34750\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__34750\,
            I => \N__34747\
        );

    \I__7921\ : Span4Mux_v
    port map (
            O => \N__34747\,
            I => \N__34744\
        );

    \I__7920\ : Span4Mux_v
    port map (
            O => \N__34744\,
            I => \N__34741\
        );

    \I__7919\ : Odrv4
    port map (
            O => \N__34741\,
            I => \V33A_OK_c\
        );

    \I__7918\ : CascadeMux
    port map (
            O => \N__34738\,
            I => \N__34735\
        );

    \I__7917\ : InMux
    port map (
            O => \N__34735\,
            I => \N__34732\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__34732\,
            I => \V5A_OK_c\
        );

    \I__7915\ : InMux
    port map (
            O => \N__34729\,
            I => \N__34726\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__34726\,
            I => \VCCST_CPU_OK_c\
        );

    \I__7913\ : CascadeMux
    port map (
            O => \N__34723\,
            I => \N__34718\
        );

    \I__7912\ : CascadeMux
    port map (
            O => \N__34722\,
            I => \N__34713\
        );

    \I__7911\ : InMux
    port map (
            O => \N__34721\,
            I => \N__34702\
        );

    \I__7910\ : InMux
    port map (
            O => \N__34718\,
            I => \N__34702\
        );

    \I__7909\ : InMux
    port map (
            O => \N__34717\,
            I => \N__34702\
        );

    \I__7908\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34702\
        );

    \I__7907\ : InMux
    port map (
            O => \N__34713\,
            I => \N__34697\
        );

    \I__7906\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34697\
        );

    \I__7905\ : InMux
    port map (
            O => \N__34711\,
            I => \N__34694\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__34702\,
            I => \N__34689\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__34697\,
            I => \N__34689\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__34694\,
            I => \N__34686\
        );

    \I__7901\ : Span12Mux_s8_v
    port map (
            O => \N__34689\,
            I => \N__34683\
        );

    \I__7900\ : Span4Mux_v
    port map (
            O => \N__34686\,
            I => \N__34680\
        );

    \I__7899\ : Odrv12
    port map (
            O => \N__34683\,
            I => \N_1661\
        );

    \I__7898\ : Odrv4
    port map (
            O => \N__34680\,
            I => \N_1661\
        );

    \I__7897\ : InMux
    port map (
            O => \N__34675\,
            I => \N__34669\
        );

    \I__7896\ : InMux
    port map (
            O => \N__34674\,
            I => \N__34669\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__34669\,
            I => \b2v_inst6.count_0_1\
        );

    \I__7894\ : CascadeMux
    port map (
            O => \N__34666\,
            I => \N__34663\
        );

    \I__7893\ : InMux
    port map (
            O => \N__34663\,
            I => \N__34654\
        );

    \I__7892\ : InMux
    port map (
            O => \N__34662\,
            I => \N__34654\
        );

    \I__7891\ : InMux
    port map (
            O => \N__34661\,
            I => \N__34654\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__34654\,
            I => \b2v_inst6.count_RNI_0_1\
        );

    \I__7889\ : InMux
    port map (
            O => \N__34651\,
            I => \N__34648\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__34648\,
            I => \N__34645\
        );

    \I__7887\ : Span4Mux_s3_v
    port map (
            O => \N__34645\,
            I => \N__34641\
        );

    \I__7886\ : InMux
    port map (
            O => \N__34644\,
            I => \N__34638\
        );

    \I__7885\ : Span4Mux_s0_h
    port map (
            O => \N__34641\,
            I => \N__34633\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__34638\,
            I => \N__34633\
        );

    \I__7883\ : Odrv4
    port map (
            O => \N__34633\,
            I => \b2v_inst6.countZ0Z_15\
        );

    \I__7882\ : CascadeMux
    port map (
            O => \N__34630\,
            I => \b2v_inst6.countZ0Z_1_cascade_\
        );

    \I__7881\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34621\
        );

    \I__7880\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34618\
        );

    \I__7879\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34615\
        );

    \I__7878\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34612\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__34621\,
            I => \N__34607\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34607\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__34615\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__7874\ : LocalMux
    port map (
            O => \N__34612\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__7873\ : Odrv12
    port map (
            O => \N__34607\,
            I => \b2v_inst6.countZ0Z_11\
        );

    \I__7872\ : InMux
    port map (
            O => \N__34600\,
            I => \N__34597\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__34597\,
            I => \N__34594\
        );

    \I__7870\ : Span4Mux_v
    port map (
            O => \N__34594\,
            I => \N__34591\
        );

    \I__7869\ : Odrv4
    port map (
            O => \N__34591\,
            I => \b2v_inst6.count_1_i_a3_8_0\
        );

    \I__7868\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34585\
        );

    \I__7867\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34582\
        );

    \I__7866\ : Odrv12
    port map (
            O => \N__34582\,
            I => \b2v_inst6.count_1_i_a3_9_0\
        );

    \I__7865\ : CascadeMux
    port map (
            O => \N__34579\,
            I => \b2v_inst6.count_1_i_a3_7_0_cascade_\
        );

    \I__7864\ : InMux
    port map (
            O => \N__34576\,
            I => \N__34573\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__34573\,
            I => \N__34570\
        );

    \I__7862\ : Span4Mux_v
    port map (
            O => \N__34570\,
            I => \N__34567\
        );

    \I__7861\ : Odrv4
    port map (
            O => \N__34567\,
            I => \b2v_inst6.count_1_i_a3_10_0\
        );

    \I__7860\ : InMux
    port map (
            O => \N__34564\,
            I => \N__34558\
        );

    \I__7859\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34558\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__34558\,
            I => \b2v_inst6.N_389\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__34555\,
            I => \b2v_inst6.N_389_cascade_\
        );

    \I__7856\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34549\
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__34549\,
            I => \b2v_inst11.mult1_un75_sum_i_8\
        );

    \I__7854\ : InMux
    port map (
            O => \N__34546\,
            I => \N__34543\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__34543\,
            I => \b2v_inst11.mult1_un96_sum_i_8\
        );

    \I__7852\ : CascadeMux
    port map (
            O => \N__34540\,
            I => \b2v_inst6.count_rst_11_cascade_\
        );

    \I__7851\ : CascadeMux
    port map (
            O => \N__34537\,
            I => \N__34532\
        );

    \I__7850\ : InMux
    port map (
            O => \N__34536\,
            I => \N__34529\
        );

    \I__7849\ : InMux
    port map (
            O => \N__34535\,
            I => \N__34526\
        );

    \I__7848\ : InMux
    port map (
            O => \N__34532\,
            I => \N__34523\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__34529\,
            I => \N__34518\
        );

    \I__7846\ : LocalMux
    port map (
            O => \N__34526\,
            I => \N__34518\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__34523\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__7844\ : Odrv12
    port map (
            O => \N__34518\,
            I => \b2v_inst6.countZ0Z_3\
        );

    \I__7843\ : InMux
    port map (
            O => \N__34513\,
            I => \N__34507\
        );

    \I__7842\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34507\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__34507\,
            I => \N__34504\
        );

    \I__7840\ : Odrv12
    port map (
            O => \N__34504\,
            I => \b2v_inst6.un2_count_1_cry_2_THRU_CO\
        );

    \I__7839\ : CascadeMux
    port map (
            O => \N__34501\,
            I => \b2v_inst6.countZ0Z_3_cascade_\
        );

    \I__7838\ : InMux
    port map (
            O => \N__34498\,
            I => \N__34495\
        );

    \I__7837\ : LocalMux
    port map (
            O => \N__34495\,
            I => \b2v_inst6.count_0_3\
        );

    \I__7836\ : CascadeMux
    port map (
            O => \N__34492\,
            I => \N__34489\
        );

    \I__7835\ : InMux
    port map (
            O => \N__34489\,
            I => \N__34485\
        );

    \I__7834\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34482\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__34485\,
            I => \N__34477\
        );

    \I__7832\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34477\
        );

    \I__7831\ : Span4Mux_v
    port map (
            O => \N__34477\,
            I => \N__34474\
        );

    \I__7830\ : Odrv4
    port map (
            O => \N__34474\,
            I => \b2v_inst6.un2_count_1_cry_10_THRU_CO\
        );

    \I__7829\ : CascadeMux
    port map (
            O => \N__34471\,
            I => \b2v_inst6.N_394_cascade_\
        );

    \I__7828\ : InMux
    port map (
            O => \N__34468\,
            I => \N__34465\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__34465\,
            I => \b2v_inst6.count_0_11\
        );

    \I__7826\ : CascadeMux
    port map (
            O => \N__34462\,
            I => \b2v_inst6.count_rst_3_cascade_\
        );

    \I__7825\ : CascadeMux
    port map (
            O => \N__34459\,
            I => \N__34456\
        );

    \I__7824\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34453\
        );

    \I__7823\ : LocalMux
    port map (
            O => \N__34453\,
            I => \N__34450\
        );

    \I__7822\ : Span4Mux_s3_v
    port map (
            O => \N__34450\,
            I => \N__34447\
        );

    \I__7821\ : Odrv4
    port map (
            O => \N__34447\,
            I => \b2v_inst6.un2_count_1_axb_1\
        );

    \I__7820\ : InMux
    port map (
            O => \N__34444\,
            I => \N__34441\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__34441\,
            I => \b2v_inst6.count_0_10\
        );

    \I__7818\ : InMux
    port map (
            O => \N__34438\,
            I => \N__34434\
        );

    \I__7817\ : InMux
    port map (
            O => \N__34437\,
            I => \N__34431\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__34434\,
            I => \N__34426\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__34431\,
            I => \N__34426\
        );

    \I__7814\ : Odrv12
    port map (
            O => \N__34426\,
            I => \b2v_inst6.un2_count_1_cry_6_THRU_CO\
        );

    \I__7813\ : InMux
    port map (
            O => \N__34423\,
            I => \N__34420\
        );

    \I__7812\ : LocalMux
    port map (
            O => \N__34420\,
            I => \N__34417\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__34417\,
            I => \b2v_inst6.count_0_7\
        );

    \I__7810\ : CascadeMux
    port map (
            O => \N__34414\,
            I => \b2v_inst6.count_rst_7_cascade_\
        );

    \I__7809\ : InMux
    port map (
            O => \N__34411\,
            I => \N__34403\
        );

    \I__7808\ : InMux
    port map (
            O => \N__34410\,
            I => \N__34403\
        );

    \I__7807\ : InMux
    port map (
            O => \N__34409\,
            I => \N__34400\
        );

    \I__7806\ : InMux
    port map (
            O => \N__34408\,
            I => \N__34397\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__34403\,
            I => \N__34392\
        );

    \I__7804\ : LocalMux
    port map (
            O => \N__34400\,
            I => \N__34392\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__34397\,
            I => \b2v_inst6.countZ0Z_7\
        );

    \I__7802\ : Odrv12
    port map (
            O => \N__34392\,
            I => \b2v_inst6.countZ0Z_7\
        );

    \I__7801\ : InMux
    port map (
            O => \N__34387\,
            I => \N__34381\
        );

    \I__7800\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34381\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__34381\,
            I => \N__34378\
        );

    \I__7798\ : Odrv4
    port map (
            O => \N__34378\,
            I => \b2v_inst6.count_rst\
        );

    \I__7797\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34372\
        );

    \I__7796\ : LocalMux
    port map (
            O => \N__34372\,
            I => \b2v_inst6.count_0_15\
        );

    \I__7795\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34366\
        );

    \I__7794\ : LocalMux
    port map (
            O => \N__34366\,
            I => \N__34363\
        );

    \I__7793\ : Span4Mux_v
    port map (
            O => \N__34363\,
            I => \N__34359\
        );

    \I__7792\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34356\
        );

    \I__7791\ : Odrv4
    port map (
            O => \N__34359\,
            I => \b2v_inst6.count_rst_12\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__34356\,
            I => \b2v_inst6.count_rst_12\
        );

    \I__7789\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34348\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__34348\,
            I => \N__34345\
        );

    \I__7787\ : Span4Mux_s1_v
    port map (
            O => \N__34345\,
            I => \N__34342\
        );

    \I__7786\ : Odrv4
    port map (
            O => \N__34342\,
            I => \b2v_inst6.count_0_2\
        );

    \I__7785\ : InMux
    port map (
            O => \N__34339\,
            I => \N__34336\
        );

    \I__7784\ : LocalMux
    port map (
            O => \N__34336\,
            I => \b2v_inst6.count_rst_6\
        );

    \I__7783\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34328\
        );

    \I__7782\ : CascadeMux
    port map (
            O => \N__34332\,
            I => \N__34325\
        );

    \I__7781\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34322\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__34328\,
            I => \N__34319\
        );

    \I__7779\ : InMux
    port map (
            O => \N__34325\,
            I => \N__34316\
        );

    \I__7778\ : LocalMux
    port map (
            O => \N__34322\,
            I => \N__34311\
        );

    \I__7777\ : Span4Mux_s1_v
    port map (
            O => \N__34319\,
            I => \N__34311\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__34316\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__7775\ : Odrv4
    port map (
            O => \N__34311\,
            I => \b2v_inst6.countZ0Z_8\
        );

    \I__7774\ : CascadeMux
    port map (
            O => \N__34306\,
            I => \b2v_inst6.countZ0Z_8_cascade_\
        );

    \I__7773\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34299\
        );

    \I__7772\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34296\
        );

    \I__7771\ : LocalMux
    port map (
            O => \N__34299\,
            I => \N__34291\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__34296\,
            I => \N__34291\
        );

    \I__7769\ : Span4Mux_v
    port map (
            O => \N__34291\,
            I => \N__34288\
        );

    \I__7768\ : Odrv4
    port map (
            O => \N__34288\,
            I => \b2v_inst6.un2_count_1_cry_7_THRU_CO\
        );

    \I__7767\ : InMux
    port map (
            O => \N__34285\,
            I => \N__34282\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__34282\,
            I => \b2v_inst6.count_0_8\
        );

    \I__7765\ : InMux
    port map (
            O => \N__34279\,
            I => \N__34276\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__34276\,
            I => \N__34273\
        );

    \I__7763\ : Odrv12
    port map (
            O => \N__34273\,
            I => \b2v_inst6.countZ0Z_10\
        );

    \I__7762\ : CascadeMux
    port map (
            O => \N__34270\,
            I => \b2v_inst6.countZ0Z_10_cascade_\
        );

    \I__7761\ : InMux
    port map (
            O => \N__34267\,
            I => \N__34264\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__34264\,
            I => \b2v_inst6.count_0_12\
        );

    \I__7759\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34255\
        );

    \I__7758\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34255\
        );

    \I__7757\ : LocalMux
    port map (
            O => \N__34255\,
            I => \N__34252\
        );

    \I__7756\ : Odrv4
    port map (
            O => \N__34252\,
            I => \b2v_inst6.count_rst_2\
        );

    \I__7755\ : CascadeMux
    port map (
            O => \N__34249\,
            I => \N__34246\
        );

    \I__7754\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34242\
        );

    \I__7753\ : InMux
    port map (
            O => \N__34245\,
            I => \N__34239\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__34242\,
            I => \N__34236\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__34239\,
            I => \b2v_inst6.countZ0Z_12\
        );

    \I__7750\ : Odrv4
    port map (
            O => \N__34236\,
            I => \b2v_inst6.countZ0Z_12\
        );

    \I__7749\ : CascadeMux
    port map (
            O => \N__34231\,
            I => \b2v_inst6.count_rst_10_cascade_\
        );

    \I__7748\ : CascadeMux
    port map (
            O => \N__34228\,
            I => \N__34224\
        );

    \I__7747\ : InMux
    port map (
            O => \N__34227\,
            I => \N__34220\
        );

    \I__7746\ : InMux
    port map (
            O => \N__34224\,
            I => \N__34217\
        );

    \I__7745\ : InMux
    port map (
            O => \N__34223\,
            I => \N__34214\
        );

    \I__7744\ : LocalMux
    port map (
            O => \N__34220\,
            I => \N__34211\
        );

    \I__7743\ : LocalMux
    port map (
            O => \N__34217\,
            I => \b2v_inst6.countZ0Z_4\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__34214\,
            I => \b2v_inst6.countZ0Z_4\
        );

    \I__7741\ : Odrv12
    port map (
            O => \N__34211\,
            I => \b2v_inst6.countZ0Z_4\
        );

    \I__7740\ : InMux
    port map (
            O => \N__34204\,
            I => \N__34198\
        );

    \I__7739\ : InMux
    port map (
            O => \N__34203\,
            I => \N__34198\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__34198\,
            I => \N__34195\
        );

    \I__7737\ : Odrv12
    port map (
            O => \N__34195\,
            I => \b2v_inst6.un2_count_1_cry_3_THRU_CO\
        );

    \I__7736\ : CascadeMux
    port map (
            O => \N__34192\,
            I => \b2v_inst6.countZ0Z_4_cascade_\
        );

    \I__7735\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34186\
        );

    \I__7734\ : LocalMux
    port map (
            O => \N__34186\,
            I => \b2v_inst6.count_0_4\
        );

    \I__7733\ : InMux
    port map (
            O => \N__34183\,
            I => \N__34177\
        );

    \I__7732\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34177\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__34177\,
            I => \N__34174\
        );

    \I__7730\ : Odrv4
    port map (
            O => \N__34174\,
            I => \b2v_inst6.count_rst_4\
        );

    \I__7729\ : InMux
    port map (
            O => \N__34171\,
            I => \b2v_inst6.un2_count_1_cry_14\
        );

    \I__7728\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34165\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__34165\,
            I => \N__34162\
        );

    \I__7726\ : Odrv4
    port map (
            O => \N__34162\,
            I => \b2v_inst6.count_0_13\
        );

    \I__7725\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34155\
        );

    \I__7724\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34152\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__34155\,
            I => \b2v_inst6.count_rst_1\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__34152\,
            I => \b2v_inst6.count_rst_1\
        );

    \I__7721\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34144\
        );

    \I__7720\ : LocalMux
    port map (
            O => \N__34144\,
            I => \N__34140\
        );

    \I__7719\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34137\
        );

    \I__7718\ : Odrv4
    port map (
            O => \N__34140\,
            I => \b2v_inst6.countZ0Z_13\
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__34137\,
            I => \b2v_inst6.countZ0Z_13\
        );

    \I__7716\ : InMux
    port map (
            O => \N__34132\,
            I => \N__34129\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__34129\,
            I => \b2v_inst6.count_0_5\
        );

    \I__7714\ : InMux
    port map (
            O => \N__34126\,
            I => \N__34120\
        );

    \I__7713\ : InMux
    port map (
            O => \N__34125\,
            I => \N__34120\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__34120\,
            I => \N__34117\
        );

    \I__7711\ : Odrv12
    port map (
            O => \N__34117\,
            I => \b2v_inst6.un2_count_1_cry_4_THRU_CO\
        );

    \I__7710\ : CascadeMux
    port map (
            O => \N__34114\,
            I => \b2v_inst6.countZ0Z_5_cascade_\
        );

    \I__7709\ : InMux
    port map (
            O => \N__34111\,
            I => \N__34108\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__34108\,
            I => \b2v_inst6.count_rst_9\
        );

    \I__7707\ : InMux
    port map (
            O => \N__34105\,
            I => \N__34102\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__34102\,
            I => \b2v_inst6.count_rst_5\
        );

    \I__7705\ : CascadeMux
    port map (
            O => \N__34099\,
            I => \b2v_inst6.countZ0Z_9_cascade_\
        );

    \I__7704\ : InMux
    port map (
            O => \N__34096\,
            I => \N__34091\
        );

    \I__7703\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34086\
        );

    \I__7702\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34086\
        );

    \I__7701\ : LocalMux
    port map (
            O => \N__34091\,
            I => \N__34083\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__34086\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__7699\ : Odrv4
    port map (
            O => \N__34083\,
            I => \b2v_inst6.countZ0Z_5\
        );

    \I__7698\ : CascadeMux
    port map (
            O => \N__34078\,
            I => \N__34075\
        );

    \I__7697\ : InMux
    port map (
            O => \N__34075\,
            I => \N__34068\
        );

    \I__7696\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34068\
        );

    \I__7695\ : InMux
    port map (
            O => \N__34073\,
            I => \N__34065\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__34068\,
            I => \b2v_inst6.countZ0Z_9\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__34065\,
            I => \b2v_inst6.countZ0Z_9\
        );

    \I__7692\ : InMux
    port map (
            O => \N__34060\,
            I => \N__34054\
        );

    \I__7691\ : InMux
    port map (
            O => \N__34059\,
            I => \N__34054\
        );

    \I__7690\ : LocalMux
    port map (
            O => \N__34054\,
            I => \b2v_inst6.un2_count_1_cry_8_THRU_CO\
        );

    \I__7689\ : InMux
    port map (
            O => \N__34051\,
            I => \N__34048\
        );

    \I__7688\ : LocalMux
    port map (
            O => \N__34048\,
            I => \b2v_inst6.count_0_9\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__34045\,
            I => \N__34041\
        );

    \I__7686\ : InMux
    port map (
            O => \N__34044\,
            I => \N__34038\
        );

    \I__7685\ : InMux
    port map (
            O => \N__34041\,
            I => \N__34035\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__34038\,
            I => \b2v_inst6.countZ0Z_6\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__34035\,
            I => \b2v_inst6.countZ0Z_6\
        );

    \I__7682\ : InMux
    port map (
            O => \N__34030\,
            I => \N__34024\
        );

    \I__7681\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34024\
        );

    \I__7680\ : LocalMux
    port map (
            O => \N__34024\,
            I => \b2v_inst6.count_rst_8\
        );

    \I__7679\ : InMux
    port map (
            O => \N__34021\,
            I => \b2v_inst6.un2_count_1_cry_5\
        );

    \I__7678\ : InMux
    port map (
            O => \N__34018\,
            I => \b2v_inst6.un2_count_1_cry_6\
        );

    \I__7677\ : InMux
    port map (
            O => \N__34015\,
            I => \b2v_inst6.un2_count_1_cry_7\
        );

    \I__7676\ : InMux
    port map (
            O => \N__34012\,
            I => \bfn_12_2_0_\
        );

    \I__7675\ : InMux
    port map (
            O => \N__34009\,
            I => \b2v_inst6.un2_count_1_cry_9\
        );

    \I__7674\ : InMux
    port map (
            O => \N__34006\,
            I => \b2v_inst6.un2_count_1_cry_10\
        );

    \I__7673\ : InMux
    port map (
            O => \N__34003\,
            I => \b2v_inst6.un2_count_1_cry_11\
        );

    \I__7672\ : InMux
    port map (
            O => \N__34000\,
            I => \b2v_inst6.un2_count_1_cry_12\
        );

    \I__7671\ : InMux
    port map (
            O => \N__33997\,
            I => \N__33994\
        );

    \I__7670\ : LocalMux
    port map (
            O => \N__33994\,
            I => \b2v_inst6.countZ0Z_14\
        );

    \I__7669\ : InMux
    port map (
            O => \N__33991\,
            I => \N__33985\
        );

    \I__7668\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33985\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__33985\,
            I => \b2v_inst6.count_rst_0\
        );

    \I__7666\ : InMux
    port map (
            O => \N__33982\,
            I => \b2v_inst6.un2_count_1_cry_13\
        );

    \I__7665\ : InMux
    port map (
            O => \N__33979\,
            I => \N__33976\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__33973\,
            I => \b2v_inst11.mult1_un159_sum_cry_4_s\
        );

    \I__7662\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33967\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33967\,
            I => \N__33962\
        );

    \I__7660\ : CascadeMux
    port map (
            O => \N__33966\,
            I => \N__33959\
        );

    \I__7659\ : CascadeMux
    port map (
            O => \N__33965\,
            I => \N__33956\
        );

    \I__7658\ : Span4Mux_v
    port map (
            O => \N__33962\,
            I => \N__33951\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33948\
        );

    \I__7656\ : InMux
    port map (
            O => \N__33956\,
            I => \N__33943\
        );

    \I__7655\ : InMux
    port map (
            O => \N__33955\,
            I => \N__33943\
        );

    \I__7654\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33940\
        );

    \I__7653\ : Span4Mux_v
    port map (
            O => \N__33951\,
            I => \N__33931\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__33948\,
            I => \N__33931\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__33943\,
            I => \N__33931\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__33940\,
            I => \N__33931\
        );

    \I__7649\ : Odrv4
    port map (
            O => \N__33931\,
            I => \b2v_inst11.mult1_un159_sum_s_7\
        );

    \I__7648\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33925\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33922\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__33922\,
            I => \b2v_inst11.mult1_un159_sum_cry_5_s\
        );

    \I__7645\ : CascadeMux
    port map (
            O => \N__33919\,
            I => \N__33915\
        );

    \I__7644\ : CascadeMux
    port map (
            O => \N__33918\,
            I => \N__33911\
        );

    \I__7643\ : InMux
    port map (
            O => \N__33915\,
            I => \N__33904\
        );

    \I__7642\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33904\
        );

    \I__7641\ : InMux
    port map (
            O => \N__33911\,
            I => \N__33904\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__33904\,
            I => \G_2836\
        );

    \I__7639\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33898\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__33898\,
            I => \N__33895\
        );

    \I__7637\ : Odrv12
    port map (
            O => \N__33895\,
            I => \b2v_inst11.mult1_un166_sum_axb_6\
        );

    \I__7636\ : InMux
    port map (
            O => \N__33892\,
            I => \b2v_inst11.mult1_un166_sum_cry_5\
        );

    \I__7635\ : CascadeMux
    port map (
            O => \N__33889\,
            I => \N__33886\
        );

    \I__7634\ : InMux
    port map (
            O => \N__33886\,
            I => \N__33883\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__33883\,
            I => \N__33880\
        );

    \I__7632\ : Span4Mux_v
    port map (
            O => \N__33880\,
            I => \N__33877\
        );

    \I__7631\ : Span4Mux_v
    port map (
            O => \N__33877\,
            I => \N__33874\
        );

    \I__7630\ : Odrv4
    port map (
            O => \N__33874\,
            I => \b2v_inst11.un85_clk_100khz_0\
        );

    \I__7629\ : InMux
    port map (
            O => \N__33871\,
            I => \N__33867\
        );

    \I__7628\ : InMux
    port map (
            O => \N__33870\,
            I => \N__33864\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__33867\,
            I => \b2v_inst6.countZ0Z_2\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__33864\,
            I => \b2v_inst6.countZ0Z_2\
        );

    \I__7625\ : InMux
    port map (
            O => \N__33859\,
            I => \b2v_inst6.un2_count_1_cry_1\
        );

    \I__7624\ : InMux
    port map (
            O => \N__33856\,
            I => \b2v_inst6.un2_count_1_cry_2\
        );

    \I__7623\ : InMux
    port map (
            O => \N__33853\,
            I => \b2v_inst6.un2_count_1_cry_3\
        );

    \I__7622\ : InMux
    port map (
            O => \N__33850\,
            I => \b2v_inst6.un2_count_1_cry_4\
        );

    \I__7621\ : CascadeMux
    port map (
            O => \N__33847\,
            I => \b2v_inst6.N_276_0_cascade_\
        );

    \I__7620\ : InMux
    port map (
            O => \N__33844\,
            I => \N__33841\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__33841\,
            I => \N__33838\
        );

    \I__7618\ : Span4Mux_v
    port map (
            O => \N__33838\,
            I => \N__33835\
        );

    \I__7617\ : Odrv4
    port map (
            O => \N__33835\,
            I => \VR_READY_VCCINAUX_c\
        );

    \I__7616\ : InMux
    port map (
            O => \N__33832\,
            I => \N__33829\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__33829\,
            I => \N__33826\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__33826\,
            I => \VR_READY_VCCIN_c\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__33823\,
            I => \b2v_inst6.N_192_cascade_\
        );

    \I__7612\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33814\
        );

    \I__7611\ : InMux
    port map (
            O => \N__33819\,
            I => \N__33814\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__33814\,
            I => \b2v_inst6.delayed_vccin_vccinaux_ok_0\
        );

    \I__7609\ : CascadeMux
    port map (
            O => \N__33811\,
            I => \b2v_inst6.curr_state_RNIUL1J2Z0Z_0_cascade_\
        );

    \I__7608\ : InMux
    port map (
            O => \N__33808\,
            I => \N__33805\
        );

    \I__7607\ : LocalMux
    port map (
            O => \N__33805\,
            I => \b2v_inst6.N_276_0\
        );

    \I__7606\ : CascadeMux
    port map (
            O => \N__33802\,
            I => \N__33798\
        );

    \I__7605\ : IoInMux
    port map (
            O => \N__33801\,
            I => \N__33793\
        );

    \I__7604\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33785\
        );

    \I__7603\ : InMux
    port map (
            O => \N__33797\,
            I => \N__33785\
        );

    \I__7602\ : InMux
    port map (
            O => \N__33796\,
            I => \N__33785\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33777\
        );

    \I__7600\ : IoInMux
    port map (
            O => \N__33792\,
            I => \N__33774\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__33785\,
            I => \N__33771\
        );

    \I__7598\ : InMux
    port map (
            O => \N__33784\,
            I => \N__33768\
        );

    \I__7597\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33765\
        );

    \I__7596\ : InMux
    port map (
            O => \N__33782\,
            I => \N__33762\
        );

    \I__7595\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33759\
        );

    \I__7594\ : CascadeMux
    port map (
            O => \N__33780\,
            I => \N__33756\
        );

    \I__7593\ : IoSpan4Mux
    port map (
            O => \N__33777\,
            I => \N__33749\
        );

    \I__7592\ : LocalMux
    port map (
            O => \N__33774\,
            I => \N__33749\
        );

    \I__7591\ : Span4Mux_v
    port map (
            O => \N__33771\,
            I => \N__33746\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__33768\,
            I => \N__33743\
        );

    \I__7589\ : LocalMux
    port map (
            O => \N__33765\,
            I => \N__33738\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__33762\,
            I => \N__33738\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__33759\,
            I => \N__33735\
        );

    \I__7586\ : InMux
    port map (
            O => \N__33756\,
            I => \N__33730\
        );

    \I__7585\ : InMux
    port map (
            O => \N__33755\,
            I => \N__33730\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__33754\,
            I => \N__33726\
        );

    \I__7583\ : Span4Mux_s3_h
    port map (
            O => \N__33749\,
            I => \N__33720\
        );

    \I__7582\ : Span4Mux_h
    port map (
            O => \N__33746\,
            I => \N__33720\
        );

    \I__7581\ : Span4Mux_v
    port map (
            O => \N__33743\,
            I => \N__33715\
        );

    \I__7580\ : Span4Mux_h
    port map (
            O => \N__33738\,
            I => \N__33715\
        );

    \I__7579\ : Span4Mux_h
    port map (
            O => \N__33735\,
            I => \N__33710\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__33730\,
            I => \N__33710\
        );

    \I__7577\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33705\
        );

    \I__7576\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33705\
        );

    \I__7575\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33702\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__33720\,
            I => \N_15_i_0_a4_1_N_3L3_1\
        );

    \I__7573\ : Odrv4
    port map (
            O => \N__33715\,
            I => \N_15_i_0_a4_1_N_3L3_1\
        );

    \I__7572\ : Odrv4
    port map (
            O => \N__33710\,
            I => \N_15_i_0_a4_1_N_3L3_1\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__33705\,
            I => \N_15_i_0_a4_1_N_3L3_1\
        );

    \I__7570\ : LocalMux
    port map (
            O => \N__33702\,
            I => \N_15_i_0_a4_1_N_3L3_1\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__33691\,
            I => \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\
        );

    \I__7568\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33680\
        );

    \I__7567\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33675\
        );

    \I__7566\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33675\
        );

    \I__7565\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33668\
        );

    \I__7564\ : InMux
    port map (
            O => \N__33684\,
            I => \N__33668\
        );

    \I__7563\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33668\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__33680\,
            I => \N__33665\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__33675\,
            I => \N__33662\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__33668\,
            I => \N__33659\
        );

    \I__7559\ : Span4Mux_s2_v
    port map (
            O => \N__33665\,
            I => \N__33656\
        );

    \I__7558\ : Span4Mux_s2_v
    port map (
            O => \N__33662\,
            I => \N__33653\
        );

    \I__7557\ : Span4Mux_s1_v
    port map (
            O => \N__33659\,
            I => \N__33650\
        );

    \I__7556\ : Span4Mux_h
    port map (
            O => \N__33656\,
            I => \N__33647\
        );

    \I__7555\ : Span4Mux_h
    port map (
            O => \N__33653\,
            I => \N__33644\
        );

    \I__7554\ : Span4Mux_h
    port map (
            O => \N__33650\,
            I => \N__33641\
        );

    \I__7553\ : Odrv4
    port map (
            O => \N__33647\,
            I => \N_222\
        );

    \I__7552\ : Odrv4
    port map (
            O => \N__33644\,
            I => \N_222\
        );

    \I__7551\ : Odrv4
    port map (
            O => \N__33641\,
            I => \N_222\
        );

    \I__7550\ : CascadeMux
    port map (
            O => \N__33634\,
            I => \N__33630\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__33633\,
            I => \N__33625\
        );

    \I__7548\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33622\
        );

    \I__7547\ : InMux
    port map (
            O => \N__33629\,
            I => \N__33618\
        );

    \I__7546\ : InMux
    port map (
            O => \N__33628\,
            I => \N__33614\
        );

    \I__7545\ : InMux
    port map (
            O => \N__33625\,
            I => \N__33610\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__33622\,
            I => \N__33607\
        );

    \I__7543\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33604\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__33618\,
            I => \N__33601\
        );

    \I__7541\ : CascadeMux
    port map (
            O => \N__33617\,
            I => \N__33598\
        );

    \I__7540\ : LocalMux
    port map (
            O => \N__33614\,
            I => \N__33592\
        );

    \I__7539\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33589\
        );

    \I__7538\ : LocalMux
    port map (
            O => \N__33610\,
            I => \N__33583\
        );

    \I__7537\ : Span4Mux_h
    port map (
            O => \N__33607\,
            I => \N__33580\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__33604\,
            I => \N__33577\
        );

    \I__7535\ : Span4Mux_h
    port map (
            O => \N__33601\,
            I => \N__33574\
        );

    \I__7534\ : InMux
    port map (
            O => \N__33598\,
            I => \N__33571\
        );

    \I__7533\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33566\
        );

    \I__7532\ : InMux
    port map (
            O => \N__33596\,
            I => \N__33566\
        );

    \I__7531\ : InMux
    port map (
            O => \N__33595\,
            I => \N__33563\
        );

    \I__7530\ : Span12Mux_s6_h
    port map (
            O => \N__33592\,
            I => \N__33558\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__33589\,
            I => \N__33558\
        );

    \I__7528\ : InMux
    port map (
            O => \N__33588\,
            I => \N__33551\
        );

    \I__7527\ : InMux
    port map (
            O => \N__33587\,
            I => \N__33551\
        );

    \I__7526\ : InMux
    port map (
            O => \N__33586\,
            I => \N__33551\
        );

    \I__7525\ : Span4Mux_h
    port map (
            O => \N__33583\,
            I => \N__33544\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__33580\,
            I => \N__33544\
        );

    \I__7523\ : Span4Mux_h
    port map (
            O => \N__33577\,
            I => \N__33544\
        );

    \I__7522\ : Odrv4
    port map (
            O => \N__33574\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__33571\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7520\ : LocalMux
    port map (
            O => \N__33566\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__33563\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7518\ : Odrv12
    port map (
            O => \N__33558\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__33551\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7516\ : Odrv4
    port map (
            O => \N__33544\,
            I => \b2v_inst11.dutycycleZ0Z_0\
        );

    \I__7515\ : InMux
    port map (
            O => \N__33529\,
            I => \N__33526\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__33526\,
            I => \N__33523\
        );

    \I__7513\ : Odrv12
    port map (
            O => \N__33523\,
            I => \b2v_inst11.mult1_un159_sum_i\
        );

    \I__7512\ : CascadeMux
    port map (
            O => \N__33520\,
            I => \N__33517\
        );

    \I__7511\ : InMux
    port map (
            O => \N__33517\,
            I => \N__33514\
        );

    \I__7510\ : LocalMux
    port map (
            O => \N__33514\,
            I => \N__33511\
        );

    \I__7509\ : Odrv4
    port map (
            O => \N__33511\,
            I => \b2v_inst11.mult1_un159_sum_cry_2_s\
        );

    \I__7508\ : InMux
    port map (
            O => \N__33508\,
            I => \N__33505\
        );

    \I__7507\ : LocalMux
    port map (
            O => \N__33505\,
            I => \N__33502\
        );

    \I__7506\ : Odrv12
    port map (
            O => \N__33502\,
            I => \b2v_inst11.mult1_un159_sum_cry_3_s\
        );

    \I__7505\ : CascadeMux
    port map (
            O => \N__33499\,
            I => \N__33496\
        );

    \I__7504\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__33493\,
            I => \N__33490\
        );

    \I__7502\ : Span4Mux_s1_h
    port map (
            O => \N__33490\,
            I => \N__33487\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__33487\,
            I => \b2v_inst11.mult1_un54_sum_cry_3_s\
        );

    \I__7500\ : InMux
    port map (
            O => \N__33484\,
            I => \b2v_inst11.mult1_un61_sum_cry_3\
        );

    \I__7499\ : InMux
    port map (
            O => \N__33481\,
            I => \N__33478\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__33478\,
            I => \N__33475\
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__33475\,
            I => \b2v_inst11.mult1_un54_sum_cry_4_s\
        );

    \I__7496\ : InMux
    port map (
            O => \N__33472\,
            I => \b2v_inst11.mult1_un61_sum_cry_4\
        );

    \I__7495\ : CascadeMux
    port map (
            O => \N__33469\,
            I => \N__33466\
        );

    \I__7494\ : InMux
    port map (
            O => \N__33466\,
            I => \N__33463\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__33463\,
            I => \N__33460\
        );

    \I__7492\ : Odrv4
    port map (
            O => \N__33460\,
            I => \b2v_inst11.mult1_un54_sum_cry_5_s\
        );

    \I__7491\ : InMux
    port map (
            O => \N__33457\,
            I => \b2v_inst11.mult1_un61_sum_cry_5\
        );

    \I__7490\ : InMux
    port map (
            O => \N__33454\,
            I => \N__33451\
        );

    \I__7489\ : LocalMux
    port map (
            O => \N__33451\,
            I => \N__33448\
        );

    \I__7488\ : Odrv4
    port map (
            O => \N__33448\,
            I => \b2v_inst11.mult1_un54_sum_cry_6_s\
        );

    \I__7487\ : InMux
    port map (
            O => \N__33445\,
            I => \b2v_inst11.mult1_un61_sum_cry_6\
        );

    \I__7486\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \N__33439\
        );

    \I__7485\ : InMux
    port map (
            O => \N__33439\,
            I => \N__33436\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__33436\,
            I => \N__33433\
        );

    \I__7483\ : Odrv4
    port map (
            O => \N__33433\,
            I => \b2v_inst11.mult1_un61_sum_axb_8\
        );

    \I__7482\ : InMux
    port map (
            O => \N__33430\,
            I => \b2v_inst11.mult1_un61_sum_cry_7\
        );

    \I__7481\ : CascadeMux
    port map (
            O => \N__33427\,
            I => \b2v_inst11.mult1_un61_sum_s_8_cascade_\
        );

    \I__7480\ : InMux
    port map (
            O => \N__33424\,
            I => \N__33421\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__33421\,
            I => \N__33418\
        );

    \I__7478\ : IoSpan4Mux
    port map (
            O => \N__33418\,
            I => \N__33415\
        );

    \I__7477\ : Odrv4
    port map (
            O => \N__33415\,
            I => \V33S_OK_c\
        );

    \I__7476\ : InMux
    port map (
            O => \N__33412\,
            I => \N__33409\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__33409\,
            I => \N__33406\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__33406\,
            I => \V5S_OK_c\
        );

    \I__7473\ : IoInMux
    port map (
            O => \N__33403\,
            I => \N__33400\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__33400\,
            I => \N__33396\
        );

    \I__7471\ : IoInMux
    port map (
            O => \N__33399\,
            I => \N__33393\
        );

    \I__7470\ : Span4Mux_s2_h
    port map (
            O => \N__33396\,
            I => \N__33390\
        );

    \I__7469\ : LocalMux
    port map (
            O => \N__33393\,
            I => \N__33387\
        );

    \I__7468\ : Span4Mux_v
    port map (
            O => \N__33390\,
            I => \N__33384\
        );

    \I__7467\ : Span12Mux_s5_h
    port map (
            O => \N__33387\,
            I => \N__33381\
        );

    \I__7466\ : Span4Mux_h
    port map (
            O => \N__33384\,
            I => \N__33378\
        );

    \I__7465\ : Span12Mux_v
    port map (
            O => \N__33381\,
            I => \N__33375\
        );

    \I__7464\ : Span4Mux_h
    port map (
            O => \N__33378\,
            I => \N__33372\
        );

    \I__7463\ : Odrv12
    port map (
            O => \N__33375\,
            I => \VCCIN_EN_c\
        );

    \I__7462\ : Odrv4
    port map (
            O => \N__33372\,
            I => \VCCIN_EN_c\
        );

    \I__7461\ : InMux
    port map (
            O => \N__33367\,
            I => \b2v_inst11.mult1_un89_sum_cry_7\
        );

    \I__7460\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33356\
        );

    \I__7459\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33349\
        );

    \I__7458\ : InMux
    port map (
            O => \N__33362\,
            I => \N__33346\
        );

    \I__7457\ : InMux
    port map (
            O => \N__33361\,
            I => \N__33343\
        );

    \I__7456\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33338\
        );

    \I__7455\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33338\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__33356\,
            I => \N__33335\
        );

    \I__7453\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33332\
        );

    \I__7452\ : CascadeMux
    port map (
            O => \N__33354\,
            I => \N__33329\
        );

    \I__7451\ : CascadeMux
    port map (
            O => \N__33353\,
            I => \N__33326\
        );

    \I__7450\ : InMux
    port map (
            O => \N__33352\,
            I => \N__33323\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__33349\,
            I => \N__33317\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__33346\,
            I => \N__33312\
        );

    \I__7447\ : LocalMux
    port map (
            O => \N__33343\,
            I => \N__33312\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__33338\,
            I => \N__33309\
        );

    \I__7445\ : Span4Mux_s2_h
    port map (
            O => \N__33335\,
            I => \N__33304\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__33332\,
            I => \N__33304\
        );

    \I__7443\ : InMux
    port map (
            O => \N__33329\,
            I => \N__33301\
        );

    \I__7442\ : InMux
    port map (
            O => \N__33326\,
            I => \N__33298\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__33323\,
            I => \N__33295\
        );

    \I__7440\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33290\
        );

    \I__7439\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33290\
        );

    \I__7438\ : InMux
    port map (
            O => \N__33320\,
            I => \N__33287\
        );

    \I__7437\ : Span4Mux_h
    port map (
            O => \N__33317\,
            I => \N__33282\
        );

    \I__7436\ : Span4Mux_h
    port map (
            O => \N__33312\,
            I => \N__33282\
        );

    \I__7435\ : Span4Mux_v
    port map (
            O => \N__33309\,
            I => \N__33277\
        );

    \I__7434\ : Span4Mux_h
    port map (
            O => \N__33304\,
            I => \N__33277\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__33301\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7432\ : LocalMux
    port map (
            O => \N__33298\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7431\ : Odrv12
    port map (
            O => \N__33295\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__33290\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__33287\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__33282\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7427\ : Odrv4
    port map (
            O => \N__33277\,
            I => \b2v_inst11.dutycycle\
        );

    \I__7426\ : InMux
    port map (
            O => \N__33262\,
            I => \N__33258\
        );

    \I__7425\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33255\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__33258\,
            I => \N__33252\
        );

    \I__7423\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33249\
        );

    \I__7422\ : Span4Mux_s2_h
    port map (
            O => \N__33252\,
            I => \N__33246\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__33249\,
            I => \N__33243\
        );

    \I__7420\ : Odrv4
    port map (
            O => \N__33246\,
            I => \b2v_inst11.mult1_un54_sum\
        );

    \I__7419\ : Odrv4
    port map (
            O => \N__33243\,
            I => \b2v_inst11.mult1_un54_sum\
        );

    \I__7418\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__7417\ : LocalMux
    port map (
            O => \N__33235\,
            I => \N__33232\
        );

    \I__7416\ : Odrv12
    port map (
            O => \N__33232\,
            I => \b2v_inst11.mult1_un61_sum_i_8\
        );

    \I__7415\ : InMux
    port map (
            O => \N__33229\,
            I => \N__33225\
        );

    \I__7414\ : InMux
    port map (
            O => \N__33228\,
            I => \N__33222\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__33225\,
            I => \N__33219\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__33222\,
            I => \N__33216\
        );

    \I__7411\ : Span4Mux_s2_h
    port map (
            O => \N__33219\,
            I => \N__33213\
        );

    \I__7410\ : Span4Mux_s2_h
    port map (
            O => \N__33216\,
            I => \N__33210\
        );

    \I__7409\ : Odrv4
    port map (
            O => \N__33213\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__7408\ : Odrv4
    port map (
            O => \N__33210\,
            I => \b2v_inst11.mult1_un61_sum\
        );

    \I__7407\ : InMux
    port map (
            O => \N__33205\,
            I => \N__33202\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__33202\,
            I => \b2v_inst11.mult1_un54_sum_i\
        );

    \I__7405\ : InMux
    port map (
            O => \N__33199\,
            I => \b2v_inst11.mult1_un61_sum_cry_2\
        );

    \I__7404\ : InMux
    port map (
            O => \N__33196\,
            I => \N__33193\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__33193\,
            I => \b2v_inst11.mult1_un89_sum_i_8\
        );

    \I__7402\ : CascadeMux
    port map (
            O => \N__33190\,
            I => \N__33187\
        );

    \I__7401\ : InMux
    port map (
            O => \N__33187\,
            I => \N__33184\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__7399\ : Span4Mux_v
    port map (
            O => \N__33181\,
            I => \N__33178\
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__33178\,
            I => \b2v_inst11.un85_clk_100khz_1\
        );

    \I__7397\ : InMux
    port map (
            O => \N__33175\,
            I => \N__33172\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__33172\,
            I => \b2v_inst11.mult1_un82_sum_i_8\
        );

    \I__7395\ : InMux
    port map (
            O => \N__33169\,
            I => \N__33165\
        );

    \I__7394\ : InMux
    port map (
            O => \N__33168\,
            I => \N__33162\
        );

    \I__7393\ : LocalMux
    port map (
            O => \N__33165\,
            I => \N__33159\
        );

    \I__7392\ : LocalMux
    port map (
            O => \N__33162\,
            I => \N__33156\
        );

    \I__7391\ : Span4Mux_s2_h
    port map (
            O => \N__33159\,
            I => \N__33153\
        );

    \I__7390\ : Odrv4
    port map (
            O => \N__33156\,
            I => \b2v_inst11.mult1_un89_sum\
        );

    \I__7389\ : Odrv4
    port map (
            O => \N__33153\,
            I => \b2v_inst11.mult1_un89_sum\
        );

    \I__7388\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33145\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__33145\,
            I => \b2v_inst11.mult1_un82_sum_i\
        );

    \I__7386\ : InMux
    port map (
            O => \N__33142\,
            I => \b2v_inst11.mult1_un89_sum_cry_2\
        );

    \I__7385\ : InMux
    port map (
            O => \N__33139\,
            I => \b2v_inst11.mult1_un89_sum_cry_3\
        );

    \I__7384\ : InMux
    port map (
            O => \N__33136\,
            I => \b2v_inst11.mult1_un89_sum_cry_4\
        );

    \I__7383\ : InMux
    port map (
            O => \N__33133\,
            I => \b2v_inst11.mult1_un89_sum_cry_5\
        );

    \I__7382\ : InMux
    port map (
            O => \N__33130\,
            I => \b2v_inst11.mult1_un89_sum_cry_6\
        );

    \I__7381\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33124\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__33124\,
            I => \N__33121\
        );

    \I__7379\ : Span4Mux_h
    port map (
            O => \N__33121\,
            I => \N__33116\
        );

    \I__7378\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33113\
        );

    \I__7377\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33110\
        );

    \I__7376\ : Odrv4
    port map (
            O => \N__33116\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__33113\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__33110\,
            I => \b2v_inst11.countZ0Z_12\
        );

    \I__7373\ : CascadeMux
    port map (
            O => \N__33103\,
            I => \N__33100\
        );

    \I__7372\ : InMux
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__7371\ : LocalMux
    port map (
            O => \N__33097\,
            I => \b2v_inst11.N_5541_i\
        );

    \I__7370\ : InMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__7369\ : LocalMux
    port map (
            O => \N__33091\,
            I => \N__33088\
        );

    \I__7368\ : Span4Mux_s3_h
    port map (
            O => \N__33088\,
            I => \N__33083\
        );

    \I__7367\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33080\
        );

    \I__7366\ : InMux
    port map (
            O => \N__33086\,
            I => \N__33077\
        );

    \I__7365\ : Odrv4
    port map (
            O => \N__33083\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__33080\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__7363\ : LocalMux
    port map (
            O => \N__33077\,
            I => \b2v_inst11.countZ0Z_13\
        );

    \I__7362\ : CascadeMux
    port map (
            O => \N__33070\,
            I => \N__33067\
        );

    \I__7361\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33064\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__33064\,
            I => \b2v_inst11.N_5542_i\
        );

    \I__7359\ : InMux
    port map (
            O => \N__33061\,
            I => \N__33058\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__33058\,
            I => \N__33055\
        );

    \I__7357\ : Span4Mux_h
    port map (
            O => \N__33055\,
            I => \N__33052\
        );

    \I__7356\ : Span4Mux_v
    port map (
            O => \N__33052\,
            I => \N__33047\
        );

    \I__7355\ : InMux
    port map (
            O => \N__33051\,
            I => \N__33044\
        );

    \I__7354\ : InMux
    port map (
            O => \N__33050\,
            I => \N__33041\
        );

    \I__7353\ : Odrv4
    port map (
            O => \N__33047\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__7352\ : LocalMux
    port map (
            O => \N__33044\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__33041\,
            I => \b2v_inst11.countZ0Z_14\
        );

    \I__7350\ : CascadeMux
    port map (
            O => \N__33034\,
            I => \N__33031\
        );

    \I__7349\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33028\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__33028\,
            I => \b2v_inst11.N_5543_i\
        );

    \I__7347\ : InMux
    port map (
            O => \N__33025\,
            I => \N__33022\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__33022\,
            I => \N__33019\
        );

    \I__7345\ : Span12Mux_s5_h
    port map (
            O => \N__33019\,
            I => \N__33014\
        );

    \I__7344\ : InMux
    port map (
            O => \N__33018\,
            I => \N__33011\
        );

    \I__7343\ : InMux
    port map (
            O => \N__33017\,
            I => \N__33008\
        );

    \I__7342\ : Odrv12
    port map (
            O => \N__33014\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__7341\ : LocalMux
    port map (
            O => \N__33011\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__7340\ : LocalMux
    port map (
            O => \N__33008\,
            I => \b2v_inst11.countZ0Z_15\
        );

    \I__7339\ : CascadeMux
    port map (
            O => \N__33001\,
            I => \N__32998\
        );

    \I__7338\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32995\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__32995\,
            I => \b2v_inst11.N_5544_i\
        );

    \I__7336\ : InMux
    port map (
            O => \N__32992\,
            I => \bfn_11_10_0_\
        );

    \I__7335\ : CascadeMux
    port map (
            O => \N__32989\,
            I => \N__32984\
        );

    \I__7334\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32978\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32978\
        );

    \I__7332\ : InMux
    port map (
            O => \N__32984\,
            I => \N__32975\
        );

    \I__7331\ : InMux
    port map (
            O => \N__32983\,
            I => \N__32972\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32969\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32966\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__32972\,
            I => \N__32961\
        );

    \I__7327\ : Span4Mux_s2_v
    port map (
            O => \N__32969\,
            I => \N__32961\
        );

    \I__7326\ : Span12Mux_s6_v
    port map (
            O => \N__32966\,
            I => \N__32958\
        );

    \I__7325\ : Span4Mux_v
    port map (
            O => \N__32961\,
            I => \N__32955\
        );

    \I__7324\ : Odrv12
    port map (
            O => \N__32958\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__7323\ : Odrv4
    port map (
            O => \N__32955\,
            I => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__7322\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32947\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__32947\,
            I => \N__32944\
        );

    \I__7320\ : Span4Mux_v
    port map (
            O => \N__32944\,
            I => \N__32941\
        );

    \I__7319\ : Span4Mux_v
    port map (
            O => \N__32941\,
            I => \N__32936\
        );

    \I__7318\ : InMux
    port map (
            O => \N__32940\,
            I => \N__32933\
        );

    \I__7317\ : InMux
    port map (
            O => \N__32939\,
            I => \N__32930\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__32936\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__32933\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__32930\,
            I => \b2v_inst11.countZ0Z_4\
        );

    \I__7313\ : CascadeMux
    port map (
            O => \N__32923\,
            I => \N__32920\
        );

    \I__7312\ : InMux
    port map (
            O => \N__32920\,
            I => \N__32917\
        );

    \I__7311\ : LocalMux
    port map (
            O => \N__32917\,
            I => \b2v_inst11.mult1_un138_sum_i_8\
        );

    \I__7310\ : InMux
    port map (
            O => \N__32914\,
            I => \N__32911\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__32911\,
            I => \b2v_inst11.N_5533_i\
        );

    \I__7308\ : InMux
    port map (
            O => \N__32908\,
            I => \N__32905\
        );

    \I__7307\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32902\
        );

    \I__7306\ : Span4Mux_v
    port map (
            O => \N__32902\,
            I => \N__32898\
        );

    \I__7305\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32895\
        );

    \I__7304\ : Span4Mux_h
    port map (
            O => \N__32898\,
            I => \N__32889\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32889\
        );

    \I__7302\ : InMux
    port map (
            O => \N__32894\,
            I => \N__32886\
        );

    \I__7301\ : Odrv4
    port map (
            O => \N__32889\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__32886\,
            I => \b2v_inst11.countZ0Z_5\
        );

    \I__7299\ : CascadeMux
    port map (
            O => \N__32881\,
            I => \N__32878\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32878\,
            I => \N__32875\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__32875\,
            I => \N__32872\
        );

    \I__7296\ : Span4Mux_v
    port map (
            O => \N__32872\,
            I => \N__32869\
        );

    \I__7295\ : Odrv4
    port map (
            O => \N__32869\,
            I => \b2v_inst11.mult1_un131_sum_i_8\
        );

    \I__7294\ : InMux
    port map (
            O => \N__32866\,
            I => \N__32863\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__32863\,
            I => \b2v_inst11.N_5534_i\
        );

    \I__7292\ : CascadeMux
    port map (
            O => \N__32860\,
            I => \N__32857\
        );

    \I__7291\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32854\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__32854\,
            I => \b2v_inst11.mult1_un124_sum_i_8\
        );

    \I__7289\ : InMux
    port map (
            O => \N__32851\,
            I => \N__32848\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__32848\,
            I => \N__32844\
        );

    \I__7287\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32841\
        );

    \I__7286\ : Span12Mux_v
    port map (
            O => \N__32844\,
            I => \N__32837\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__32841\,
            I => \N__32834\
        );

    \I__7284\ : InMux
    port map (
            O => \N__32840\,
            I => \N__32831\
        );

    \I__7283\ : Odrv12
    port map (
            O => \N__32837\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__7282\ : Odrv4
    port map (
            O => \N__32834\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__32831\,
            I => \b2v_inst11.countZ0Z_6\
        );

    \I__7280\ : InMux
    port map (
            O => \N__32824\,
            I => \N__32821\
        );

    \I__7279\ : LocalMux
    port map (
            O => \N__32821\,
            I => \b2v_inst11.N_5535_i\
        );

    \I__7278\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32815\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__32815\,
            I => \N__32812\
        );

    \I__7276\ : Span4Mux_v
    port map (
            O => \N__32812\,
            I => \N__32808\
        );

    \I__7275\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32805\
        );

    \I__7274\ : Span4Mux_v
    port map (
            O => \N__32808\,
            I => \N__32801\
        );

    \I__7273\ : LocalMux
    port map (
            O => \N__32805\,
            I => \N__32798\
        );

    \I__7272\ : InMux
    port map (
            O => \N__32804\,
            I => \N__32795\
        );

    \I__7271\ : Span4Mux_h
    port map (
            O => \N__32801\,
            I => \N__32788\
        );

    \I__7270\ : Span4Mux_s3_v
    port map (
            O => \N__32798\,
            I => \N__32788\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__32795\,
            I => \N__32788\
        );

    \I__7268\ : Odrv4
    port map (
            O => \N__32788\,
            I => \b2v_inst11.countZ0Z_7\
        );

    \I__7267\ : CascadeMux
    port map (
            O => \N__32785\,
            I => \N__32782\
        );

    \I__7266\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32779\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__32779\,
            I => \b2v_inst11.mult1_un117_sum_i_8\
        );

    \I__7264\ : InMux
    port map (
            O => \N__32776\,
            I => \N__32773\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__32773\,
            I => \b2v_inst11.N_5536_i\
        );

    \I__7262\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32767\
        );

    \I__7261\ : LocalMux
    port map (
            O => \N__32767\,
            I => \N__32763\
        );

    \I__7260\ : InMux
    port map (
            O => \N__32766\,
            I => \N__32760\
        );

    \I__7259\ : Span12Mux_s4_h
    port map (
            O => \N__32763\,
            I => \N__32756\
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__32760\,
            I => \N__32753\
        );

    \I__7257\ : InMux
    port map (
            O => \N__32759\,
            I => \N__32750\
        );

    \I__7256\ : Odrv12
    port map (
            O => \N__32756\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__7255\ : Odrv4
    port map (
            O => \N__32753\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__32750\,
            I => \b2v_inst11.countZ0Z_8\
        );

    \I__7253\ : InMux
    port map (
            O => \N__32743\,
            I => \N__32740\
        );

    \I__7252\ : LocalMux
    port map (
            O => \N__32740\,
            I => \N__32737\
        );

    \I__7251\ : Odrv4
    port map (
            O => \N__32737\,
            I => \b2v_inst11.mult1_un110_sum_i_8\
        );

    \I__7250\ : CascadeMux
    port map (
            O => \N__32734\,
            I => \N__32731\
        );

    \I__7249\ : InMux
    port map (
            O => \N__32731\,
            I => \N__32728\
        );

    \I__7248\ : LocalMux
    port map (
            O => \N__32728\,
            I => \b2v_inst11.N_5537_i\
        );

    \I__7247\ : InMux
    port map (
            O => \N__32725\,
            I => \N__32722\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__32722\,
            I => \N__32719\
        );

    \I__7245\ : Span4Mux_v
    port map (
            O => \N__32719\,
            I => \N__32715\
        );

    \I__7244\ : InMux
    port map (
            O => \N__32718\,
            I => \N__32712\
        );

    \I__7243\ : Span4Mux_h
    port map (
            O => \N__32715\,
            I => \N__32706\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__32712\,
            I => \N__32706\
        );

    \I__7241\ : InMux
    port map (
            O => \N__32711\,
            I => \N__32703\
        );

    \I__7240\ : Span4Mux_v
    port map (
            O => \N__32706\,
            I => \N__32700\
        );

    \I__7239\ : LocalMux
    port map (
            O => \N__32703\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__32700\,
            I => \b2v_inst11.countZ0Z_9\
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__32695\,
            I => \N__32692\
        );

    \I__7236\ : InMux
    port map (
            O => \N__32692\,
            I => \N__32689\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__32689\,
            I => \N__32686\
        );

    \I__7234\ : Span4Mux_s3_h
    port map (
            O => \N__32686\,
            I => \N__32683\
        );

    \I__7233\ : Odrv4
    port map (
            O => \N__32683\,
            I => \b2v_inst11.mult1_un103_sum_i_8\
        );

    \I__7232\ : InMux
    port map (
            O => \N__32680\,
            I => \N__32677\
        );

    \I__7231\ : LocalMux
    port map (
            O => \N__32677\,
            I => \b2v_inst11.N_5538_i\
        );

    \I__7230\ : InMux
    port map (
            O => \N__32674\,
            I => \N__32670\
        );

    \I__7229\ : CascadeMux
    port map (
            O => \N__32673\,
            I => \N__32667\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__32670\,
            I => \N__32664\
        );

    \I__7227\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32661\
        );

    \I__7226\ : Span4Mux_v
    port map (
            O => \N__32664\,
            I => \N__32658\
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32654\
        );

    \I__7224\ : Span4Mux_h
    port map (
            O => \N__32658\,
            I => \N__32651\
        );

    \I__7223\ : InMux
    port map (
            O => \N__32657\,
            I => \N__32648\
        );

    \I__7222\ : Span4Mux_h
    port map (
            O => \N__32654\,
            I => \N__32645\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__32651\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__32648\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__7219\ : Odrv4
    port map (
            O => \N__32645\,
            I => \b2v_inst11.countZ0Z_10\
        );

    \I__7218\ : CascadeMux
    port map (
            O => \N__32638\,
            I => \N__32635\
        );

    \I__7217\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32632\
        );

    \I__7216\ : LocalMux
    port map (
            O => \N__32632\,
            I => \b2v_inst11.N_5539_i\
        );

    \I__7215\ : InMux
    port map (
            O => \N__32629\,
            I => \N__32626\
        );

    \I__7214\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32622\
        );

    \I__7213\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32619\
        );

    \I__7212\ : Span4Mux_v
    port map (
            O => \N__32622\,
            I => \N__32616\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__32619\,
            I => \N__32612\
        );

    \I__7210\ : Span4Mux_h
    port map (
            O => \N__32616\,
            I => \N__32609\
        );

    \I__7209\ : InMux
    port map (
            O => \N__32615\,
            I => \N__32606\
        );

    \I__7208\ : Span4Mux_h
    port map (
            O => \N__32612\,
            I => \N__32603\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__32609\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__32606\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__7205\ : Odrv4
    port map (
            O => \N__32603\,
            I => \b2v_inst11.countZ0Z_11\
        );

    \I__7204\ : CascadeMux
    port map (
            O => \N__32596\,
            I => \N__32593\
        );

    \I__7203\ : InMux
    port map (
            O => \N__32593\,
            I => \N__32590\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__32590\,
            I => \b2v_inst11.N_5540_i\
        );

    \I__7201\ : InMux
    port map (
            O => \N__32587\,
            I => \N__32583\
        );

    \I__7200\ : CascadeMux
    port map (
            O => \N__32586\,
            I => \N__32579\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__32583\,
            I => \N__32575\
        );

    \I__7198\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32570\
        );

    \I__7197\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32570\
        );

    \I__7196\ : InMux
    port map (
            O => \N__32578\,
            I => \N__32567\
        );

    \I__7195\ : Odrv12
    port map (
            O => \N__32575\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__32570\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__32567\,
            I => \b2v_inst11.mult1_un117_sum_s_8\
        );

    \I__7192\ : InMux
    port map (
            O => \N__32560\,
            I => \N__32557\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__32557\,
            I => \N__32553\
        );

    \I__7190\ : CascadeMux
    port map (
            O => \N__32556\,
            I => \N__32549\
        );

    \I__7189\ : Span4Mux_h
    port map (
            O => \N__32553\,
            I => \N__32543\
        );

    \I__7188\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32540\
        );

    \I__7187\ : InMux
    port map (
            O => \N__32549\,
            I => \N__32533\
        );

    \I__7186\ : InMux
    port map (
            O => \N__32548\,
            I => \N__32533\
        );

    \I__7185\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32533\
        );

    \I__7184\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32530\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__32543\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__32540\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__32533\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__32530\,
            I => \b2v_inst11.mult1_un124_sum_s_8\
        );

    \I__7179\ : InMux
    port map (
            O => \N__32521\,
            I => \N__32516\
        );

    \I__7178\ : CascadeMux
    port map (
            O => \N__32520\,
            I => \N__32513\
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__32519\,
            I => \N__32510\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__32516\,
            I => \N__32506\
        );

    \I__7175\ : InMux
    port map (
            O => \N__32513\,
            I => \N__32503\
        );

    \I__7174\ : InMux
    port map (
            O => \N__32510\,
            I => \N__32498\
        );

    \I__7173\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32498\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__32506\,
            I => \N__32494\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__32503\,
            I => \N__32489\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__32498\,
            I => \N__32489\
        );

    \I__7169\ : InMux
    port map (
            O => \N__32497\,
            I => \N__32486\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__32494\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__7167\ : Odrv4
    port map (
            O => \N__32489\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__32486\,
            I => \b2v_inst11.mult1_un145_sum_s_8\
        );

    \I__7165\ : InMux
    port map (
            O => \N__32479\,
            I => \N__32476\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__32476\,
            I => \N__32472\
        );

    \I__7163\ : CascadeMux
    port map (
            O => \N__32475\,
            I => \N__32469\
        );

    \I__7162\ : Span4Mux_v
    port map (
            O => \N__32472\,
            I => \N__32463\
        );

    \I__7161\ : InMux
    port map (
            O => \N__32469\,
            I => \N__32456\
        );

    \I__7160\ : InMux
    port map (
            O => \N__32468\,
            I => \N__32456\
        );

    \I__7159\ : InMux
    port map (
            O => \N__32467\,
            I => \N__32456\
        );

    \I__7158\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32453\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__32463\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__32456\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__32453\,
            I => \b2v_inst11.mult1_un138_sum_s_8\
        );

    \I__7154\ : InMux
    port map (
            O => \N__32446\,
            I => \N__32443\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__32443\,
            I => \N__32440\
        );

    \I__7152\ : Span4Mux_v
    port map (
            O => \N__32440\,
            I => \N__32433\
        );

    \I__7151\ : InMux
    port map (
            O => \N__32439\,
            I => \N__32430\
        );

    \I__7150\ : InMux
    port map (
            O => \N__32438\,
            I => \N__32427\
        );

    \I__7149\ : InMux
    port map (
            O => \N__32437\,
            I => \N__32422\
        );

    \I__7148\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32422\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__32433\,
            I => \N__32417\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__32430\,
            I => \N__32417\
        );

    \I__7145\ : LocalMux
    port map (
            O => \N__32427\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__32422\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__7143\ : Odrv4
    port map (
            O => \N__32417\,
            I => \b2v_inst11.countZ0Z_0\
        );

    \I__7142\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32407\
        );

    \I__7141\ : LocalMux
    port map (
            O => \N__32407\,
            I => \b2v_inst11.un1_count_cry_0_i\
        );

    \I__7140\ : InMux
    port map (
            O => \N__32404\,
            I => \N__32401\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__32401\,
            I => \N__32397\
        );

    \I__7138\ : CascadeMux
    port map (
            O => \N__32400\,
            I => \N__32394\
        );

    \I__7137\ : Span4Mux_v
    port map (
            O => \N__32397\,
            I => \N__32390\
        );

    \I__7136\ : InMux
    port map (
            O => \N__32394\,
            I => \N__32387\
        );

    \I__7135\ : InMux
    port map (
            O => \N__32393\,
            I => \N__32384\
        );

    \I__7134\ : Span4Mux_h
    port map (
            O => \N__32390\,
            I => \N__32379\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__32387\,
            I => \N__32379\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__32384\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__32379\,
            I => \b2v_inst11.countZ0Z_1\
        );

    \I__7130\ : InMux
    port map (
            O => \N__32374\,
            I => \N__32371\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__32371\,
            I => \b2v_inst11.N_5530_i\
        );

    \I__7128\ : InMux
    port map (
            O => \N__32368\,
            I => \N__32365\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__32365\,
            I => \N__32362\
        );

    \I__7126\ : Span4Mux_s1_h
    port map (
            O => \N__32362\,
            I => \N__32358\
        );

    \I__7125\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32354\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__32358\,
            I => \N__32351\
        );

    \I__7123\ : InMux
    port map (
            O => \N__32357\,
            I => \N__32348\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__32354\,
            I => \N__32345\
        );

    \I__7121\ : Span4Mux_h
    port map (
            O => \N__32351\,
            I => \N__32340\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__32348\,
            I => \N__32340\
        );

    \I__7119\ : Span4Mux_h
    port map (
            O => \N__32345\,
            I => \N__32337\
        );

    \I__7118\ : Odrv4
    port map (
            O => \N__32340\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__7117\ : Odrv4
    port map (
            O => \N__32337\,
            I => \b2v_inst11.countZ0Z_2\
        );

    \I__7116\ : CascadeMux
    port map (
            O => \N__32332\,
            I => \N__32329\
        );

    \I__7115\ : InMux
    port map (
            O => \N__32329\,
            I => \N__32326\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__32326\,
            I => \b2v_inst11.un85_clk_100khz_2\
        );

    \I__7113\ : InMux
    port map (
            O => \N__32323\,
            I => \N__32320\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__32320\,
            I => \b2v_inst11.N_5531_i\
        );

    \I__7111\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32314\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__32314\,
            I => \N__32311\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__32311\,
            I => \N__32307\
        );

    \I__7108\ : CascadeMux
    port map (
            O => \N__32310\,
            I => \N__32303\
        );

    \I__7107\ : Span4Mux_v
    port map (
            O => \N__32307\,
            I => \N__32300\
        );

    \I__7106\ : InMux
    port map (
            O => \N__32306\,
            I => \N__32297\
        );

    \I__7105\ : InMux
    port map (
            O => \N__32303\,
            I => \N__32294\
        );

    \I__7104\ : Odrv4
    port map (
            O => \N__32300\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__32297\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__32294\,
            I => \b2v_inst11.countZ0Z_3\
        );

    \I__7101\ : CascadeMux
    port map (
            O => \N__32287\,
            I => \N__32284\
        );

    \I__7100\ : InMux
    port map (
            O => \N__32284\,
            I => \N__32281\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__32281\,
            I => \N__32278\
        );

    \I__7098\ : Odrv4
    port map (
            O => \N__32278\,
            I => \b2v_inst11.mult1_un145_sum_i_8\
        );

    \I__7097\ : InMux
    port map (
            O => \N__32275\,
            I => \N__32272\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__32272\,
            I => \b2v_inst11.N_5532_i\
        );

    \I__7095\ : InMux
    port map (
            O => \N__32269\,
            I => \N__32266\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__32266\,
            I => \N__32263\
        );

    \I__7093\ : Odrv12
    port map (
            O => \N__32263\,
            I => \b2v_inst5.un2_count_1_axb_5\
        );

    \I__7092\ : InMux
    port map (
            O => \N__32260\,
            I => \N__32257\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__32257\,
            I => \b2v_inst5.count_1_6\
        );

    \I__7090\ : InMux
    port map (
            O => \N__32254\,
            I => \N__32248\
        );

    \I__7089\ : InMux
    port map (
            O => \N__32253\,
            I => \N__32248\
        );

    \I__7088\ : LocalMux
    port map (
            O => \N__32248\,
            I => \N__32245\
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__32245\,
            I => \b2v_inst5.count_rst_8\
        );

    \I__7086\ : InMux
    port map (
            O => \N__32242\,
            I => \N__32239\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__32239\,
            I => \N__32236\
        );

    \I__7084\ : Odrv12
    port map (
            O => \N__32236\,
            I => \b2v_inst5.countZ0Z_6\
        );

    \I__7083\ : InMux
    port map (
            O => \N__32233\,
            I => \N__32228\
        );

    \I__7082\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32223\
        );

    \I__7081\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32223\
        );

    \I__7080\ : LocalMux
    port map (
            O => \N__32228\,
            I => \N__32218\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__32223\,
            I => \N__32218\
        );

    \I__7078\ : Odrv4
    port map (
            O => \N__32218\,
            I => \b2v_inst5.count_rst_9\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__32215\,
            I => \b2v_inst5.countZ0Z_6_cascade_\
        );

    \I__7076\ : InMux
    port map (
            O => \N__32212\,
            I => \N__32206\
        );

    \I__7075\ : InMux
    port map (
            O => \N__32211\,
            I => \N__32206\
        );

    \I__7074\ : LocalMux
    port map (
            O => \N__32206\,
            I => \b2v_inst5.count_1_5\
        );

    \I__7073\ : InMux
    port map (
            O => \N__32203\,
            I => \N__32200\
        );

    \I__7072\ : LocalMux
    port map (
            O => \N__32200\,
            I => \N__32197\
        );

    \I__7071\ : Span4Mux_v
    port map (
            O => \N__32197\,
            I => \N__32194\
        );

    \I__7070\ : Odrv4
    port map (
            O => \N__32194\,
            I => \b2v_inst5.un12_clk_100khz_3\
        );

    \I__7069\ : InMux
    port map (
            O => \N__32191\,
            I => \N__32188\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__32188\,
            I => \N__32185\
        );

    \I__7067\ : Odrv4
    port map (
            O => \N__32185\,
            I => \b2v_inst5.un2_count_1_axb_7\
        );

    \I__7066\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32163\
        );

    \I__7065\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32163\
        );

    \I__7064\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32163\
        );

    \I__7063\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32160\
        );

    \I__7062\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32155\
        );

    \I__7061\ : InMux
    port map (
            O => \N__32177\,
            I => \N__32155\
        );

    \I__7060\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32150\
        );

    \I__7059\ : InMux
    port map (
            O => \N__32175\,
            I => \N__32150\
        );

    \I__7058\ : SRMux
    port map (
            O => \N__32174\,
            I => \N__32147\
        );

    \I__7057\ : SRMux
    port map (
            O => \N__32173\,
            I => \N__32144\
        );

    \I__7056\ : SRMux
    port map (
            O => \N__32172\,
            I => \N__32136\
        );

    \I__7055\ : SRMux
    port map (
            O => \N__32171\,
            I => \N__32132\
        );

    \I__7054\ : SRMux
    port map (
            O => \N__32170\,
            I => \N__32129\
        );

    \I__7053\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32120\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__32160\,
            I => \N__32120\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__32155\,
            I => \N__32120\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__32150\,
            I => \N__32120\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__32147\,
            I => \N__32117\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__32144\,
            I => \N__32114\
        );

    \I__7047\ : InMux
    port map (
            O => \N__32143\,
            I => \N__32103\
        );

    \I__7046\ : InMux
    port map (
            O => \N__32142\,
            I => \N__32103\
        );

    \I__7045\ : InMux
    port map (
            O => \N__32141\,
            I => \N__32103\
        );

    \I__7044\ : InMux
    port map (
            O => \N__32140\,
            I => \N__32103\
        );

    \I__7043\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32103\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__32100\
        );

    \I__7041\ : SRMux
    port map (
            O => \N__32135\,
            I => \N__32097\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__32132\,
            I => \N__32082\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__32129\,
            I => \N__32077\
        );

    \I__7038\ : Span4Mux_s3_v
    port map (
            O => \N__32120\,
            I => \N__32077\
        );

    \I__7037\ : Span4Mux_s1_h
    port map (
            O => \N__32117\,
            I => \N__32070\
        );

    \I__7036\ : Span4Mux_h
    port map (
            O => \N__32114\,
            I => \N__32070\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__32103\,
            I => \N__32070\
        );

    \I__7034\ : Span4Mux_v
    port map (
            O => \N__32100\,
            I => \N__32067\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N__32064\
        );

    \I__7032\ : InMux
    port map (
            O => \N__32096\,
            I => \N__32057\
        );

    \I__7031\ : InMux
    port map (
            O => \N__32095\,
            I => \N__32057\
        );

    \I__7030\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32057\
        );

    \I__7029\ : InMux
    port map (
            O => \N__32093\,
            I => \N__32046\
        );

    \I__7028\ : SRMux
    port map (
            O => \N__32092\,
            I => \N__32046\
        );

    \I__7027\ : InMux
    port map (
            O => \N__32091\,
            I => \N__32046\
        );

    \I__7026\ : InMux
    port map (
            O => \N__32090\,
            I => \N__32046\
        );

    \I__7025\ : InMux
    port map (
            O => \N__32089\,
            I => \N__32046\
        );

    \I__7024\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32037\
        );

    \I__7023\ : InMux
    port map (
            O => \N__32087\,
            I => \N__32037\
        );

    \I__7022\ : InMux
    port map (
            O => \N__32086\,
            I => \N__32037\
        );

    \I__7021\ : InMux
    port map (
            O => \N__32085\,
            I => \N__32037\
        );

    \I__7020\ : Span4Mux_v
    port map (
            O => \N__32082\,
            I => \N__32032\
        );

    \I__7019\ : Span4Mux_v
    port map (
            O => \N__32077\,
            I => \N__32032\
        );

    \I__7018\ : Span4Mux_v
    port map (
            O => \N__32070\,
            I => \N__32029\
        );

    \I__7017\ : Span4Mux_v
    port map (
            O => \N__32067\,
            I => \N__32026\
        );

    \I__7016\ : Span4Mux_v
    port map (
            O => \N__32064\,
            I => \N__32023\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__32057\,
            I => \N__32020\
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__32046\,
            I => \N__32015\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__32037\,
            I => \N__32015\
        );

    \I__7012\ : Span4Mux_v
    port map (
            O => \N__32032\,
            I => \N__32010\
        );

    \I__7011\ : Span4Mux_v
    port map (
            O => \N__32029\,
            I => \N__32010\
        );

    \I__7010\ : Span4Mux_h
    port map (
            O => \N__32026\,
            I => \N__32007\
        );

    \I__7009\ : Span4Mux_h
    port map (
            O => \N__32023\,
            I => \N__32002\
        );

    \I__7008\ : Span4Mux_v
    port map (
            O => \N__32020\,
            I => \N__32002\
        );

    \I__7007\ : Span12Mux_v
    port map (
            O => \N__32015\,
            I => \N__31999\
        );

    \I__7006\ : Span4Mux_h
    port map (
            O => \N__32010\,
            I => \N__31996\
        );

    \I__7005\ : Odrv4
    port map (
            O => \N__32007\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7004\ : Odrv4
    port map (
            O => \N__32002\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7003\ : Odrv12
    port map (
            O => \N__31999\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7002\ : Odrv4
    port map (
            O => \N__31996\,
            I => \b2v_inst5.count_0_sqmuxa\
        );

    \I__7001\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31981\
        );

    \I__7000\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31981\
        );

    \I__6999\ : LocalMux
    port map (
            O => \N__31981\,
            I => \b2v_inst5.count_1_7\
        );

    \I__6998\ : InMux
    port map (
            O => \N__31978\,
            I => \N__31969\
        );

    \I__6997\ : InMux
    port map (
            O => \N__31977\,
            I => \N__31969\
        );

    \I__6996\ : InMux
    port map (
            O => \N__31976\,
            I => \N__31969\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__31969\,
            I => \N__31966\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__31966\,
            I => \b2v_inst5.count_rst_7\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__31963\,
            I => \N__31960\
        );

    \I__6992\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31957\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31953\
        );

    \I__6990\ : InMux
    port map (
            O => \N__31956\,
            I => \N__31950\
        );

    \I__6989\ : Span4Mux_v
    port map (
            O => \N__31953\,
            I => \N__31945\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__31950\,
            I => \N__31945\
        );

    \I__6987\ : Odrv4
    port map (
            O => \N__31945\,
            I => \b2v_inst5.countZ0Z_11\
        );

    \I__6986\ : InMux
    port map (
            O => \N__31942\,
            I => \N__31934\
        );

    \I__6985\ : CEMux
    port map (
            O => \N__31941\,
            I => \N__31934\
        );

    \I__6984\ : InMux
    port map (
            O => \N__31940\,
            I => \N__31929\
        );

    \I__6983\ : CEMux
    port map (
            O => \N__31939\,
            I => \N__31929\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__31934\,
            I => \N__31924\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__31929\,
            I => \N__31921\
        );

    \I__6980\ : CEMux
    port map (
            O => \N__31928\,
            I => \N__31918\
        );

    \I__6979\ : CEMux
    port map (
            O => \N__31927\,
            I => \N__31915\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__31924\,
            I => \N__31900\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__31921\,
            I => \N__31900\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__31918\,
            I => \N__31900\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__31915\,
            I => \N__31897\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31914\,
            I => \N__31888\
        );

    \I__6973\ : InMux
    port map (
            O => \N__31913\,
            I => \N__31888\
        );

    \I__6972\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31888\
        );

    \I__6971\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31888\
        );

    \I__6970\ : InMux
    port map (
            O => \N__31910\,
            I => \N__31875\
        );

    \I__6969\ : CEMux
    port map (
            O => \N__31909\,
            I => \N__31875\
        );

    \I__6968\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31865\
        );

    \I__6967\ : CEMux
    port map (
            O => \N__31907\,
            I => \N__31865\
        );

    \I__6966\ : Span4Mux_s3_v
    port map (
            O => \N__31900\,
            I => \N__31858\
        );

    \I__6965\ : Span4Mux_s1_h
    port map (
            O => \N__31897\,
            I => \N__31858\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31858\
        );

    \I__6963\ : InMux
    port map (
            O => \N__31887\,
            I => \N__31849\
        );

    \I__6962\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31849\
        );

    \I__6961\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31849\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31849\
        );

    \I__6959\ : CEMux
    port map (
            O => \N__31883\,
            I => \N__31840\
        );

    \I__6958\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31840\
        );

    \I__6957\ : InMux
    port map (
            O => \N__31881\,
            I => \N__31840\
        );

    \I__6956\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31840\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__31875\,
            I => \N__31837\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31874\,
            I => \N__31828\
        );

    \I__6953\ : InMux
    port map (
            O => \N__31873\,
            I => \N__31828\
        );

    \I__6952\ : InMux
    port map (
            O => \N__31872\,
            I => \N__31828\
        );

    \I__6951\ : InMux
    port map (
            O => \N__31871\,
            I => \N__31823\
        );

    \I__6950\ : InMux
    port map (
            O => \N__31870\,
            I => \N__31823\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__31865\,
            I => \N__31820\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__31858\,
            I => \N__31813\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__31849\,
            I => \N__31813\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31813\
        );

    \I__6945\ : Span4Mux_h
    port map (
            O => \N__31837\,
            I => \N__31810\
        );

    \I__6944\ : InMux
    port map (
            O => \N__31836\,
            I => \N__31805\
        );

    \I__6943\ : InMux
    port map (
            O => \N__31835\,
            I => \N__31805\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__31828\,
            I => \N__31800\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__31823\,
            I => \N__31800\
        );

    \I__6940\ : Span4Mux_v
    port map (
            O => \N__31820\,
            I => \N__31795\
        );

    \I__6939\ : Span4Mux_v
    port map (
            O => \N__31813\,
            I => \N__31795\
        );

    \I__6938\ : Span4Mux_v
    port map (
            O => \N__31810\,
            I => \N__31792\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__31805\,
            I => \N__31789\
        );

    \I__6936\ : Sp12to4
    port map (
            O => \N__31800\,
            I => \N__31786\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__31795\,
            I => \N__31783\
        );

    \I__6934\ : Span4Mux_v
    port map (
            O => \N__31792\,
            I => \N__31780\
        );

    \I__6933\ : Span4Mux_v
    port map (
            O => \N__31789\,
            I => \N__31777\
        );

    \I__6932\ : Span12Mux_v
    port map (
            O => \N__31786\,
            I => \N__31774\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__31783\,
            I => \N__31771\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__31780\,
            I => \b2v_inst5.curr_state_RNIFLPH1Z0Z_1\
        );

    \I__6929\ : Odrv4
    port map (
            O => \N__31777\,
            I => \b2v_inst5.curr_state_RNIFLPH1Z0Z_1\
        );

    \I__6928\ : Odrv12
    port map (
            O => \N__31774\,
            I => \b2v_inst5.curr_state_RNIFLPH1Z0Z_1\
        );

    \I__6927\ : Odrv4
    port map (
            O => \N__31771\,
            I => \b2v_inst5.curr_state_RNIFLPH1Z0Z_1\
        );

    \I__6926\ : CascadeMux
    port map (
            O => \N__31762\,
            I => \N__31759\
        );

    \I__6925\ : InMux
    port map (
            O => \N__31759\,
            I => \N__31756\
        );

    \I__6924\ : LocalMux
    port map (
            O => \N__31756\,
            I => \N__31753\
        );

    \I__6923\ : Span4Mux_v
    port map (
            O => \N__31753\,
            I => \N__31750\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__31750\,
            I => \b2v_inst5.un12_clk_100khz_2\
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__31747\,
            I => \N__31743\
        );

    \I__6920\ : CascadeMux
    port map (
            O => \N__31746\,
            I => \N__31740\
        );

    \I__6919\ : InMux
    port map (
            O => \N__31743\,
            I => \N__31736\
        );

    \I__6918\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31731\
        );

    \I__6917\ : InMux
    port map (
            O => \N__31739\,
            I => \N__31731\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__31736\,
            I => \N__31727\
        );

    \I__6915\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31724\
        );

    \I__6914\ : InMux
    port map (
            O => \N__31730\,
            I => \N__31721\
        );

    \I__6913\ : Span4Mux_s2_v
    port map (
            O => \N__31727\,
            I => \N__31716\
        );

    \I__6912\ : Span4Mux_s2_v
    port map (
            O => \N__31724\,
            I => \N__31716\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__31721\,
            I => \N__31713\
        );

    \I__6910\ : Span4Mux_v
    port map (
            O => \N__31716\,
            I => \N__31710\
        );

    \I__6909\ : Span4Mux_v
    port map (
            O => \N__31713\,
            I => \N__31707\
        );

    \I__6908\ : Span4Mux_v
    port map (
            O => \N__31710\,
            I => \N__31703\
        );

    \I__6907\ : Sp12to4
    port map (
            O => \N__31707\,
            I => \N__31700\
        );

    \I__6906\ : InMux
    port map (
            O => \N__31706\,
            I => \N__31697\
        );

    \I__6905\ : Odrv4
    port map (
            O => \N__31703\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__6904\ : Odrv12
    port map (
            O => \N__31700\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__31697\,
            I => \b2v_inst11.mult1_un152_sum_s_8\
        );

    \I__6902\ : InMux
    port map (
            O => \N__31690\,
            I => \N__31686\
        );

    \I__6901\ : CascadeMux
    port map (
            O => \N__31689\,
            I => \N__31682\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__31686\,
            I => \N__31678\
        );

    \I__6899\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31673\
        );

    \I__6898\ : InMux
    port map (
            O => \N__31682\,
            I => \N__31673\
        );

    \I__6897\ : InMux
    port map (
            O => \N__31681\,
            I => \N__31670\
        );

    \I__6896\ : Odrv4
    port map (
            O => \N__31678\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__31673\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__31670\,
            I => \b2v_inst11.mult1_un110_sum_s_8\
        );

    \I__6893\ : CascadeMux
    port map (
            O => \N__31663\,
            I => \b2v_inst5.count_rst_5_cascade_\
        );

    \I__6892\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31656\
        );

    \I__6891\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31653\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__31656\,
            I => \b2v_inst5.un2_count_1_axb_9\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__31653\,
            I => \b2v_inst5.un2_count_1_axb_9\
        );

    \I__6888\ : CascadeMux
    port map (
            O => \N__31648\,
            I => \N__31644\
        );

    \I__6887\ : InMux
    port map (
            O => \N__31647\,
            I => \N__31639\
        );

    \I__6886\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31639\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__31639\,
            I => \b2v_inst5.un2_count_1_cry_8_THRU_CO\
        );

    \I__6884\ : CascadeMux
    port map (
            O => \N__31636\,
            I => \b2v_inst5.un2_count_1_axb_9_cascade_\
        );

    \I__6883\ : InMux
    port map (
            O => \N__31633\,
            I => \N__31627\
        );

    \I__6882\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31627\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__31627\,
            I => \b2v_inst5.count_1_9\
        );

    \I__6880\ : CascadeMux
    port map (
            O => \N__31624\,
            I => \N__31621\
        );

    \I__6879\ : InMux
    port map (
            O => \N__31621\,
            I => \N__31618\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__31618\,
            I => \b2v_inst5.count_rst_5\
        );

    \I__6877\ : InMux
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__6875\ : Span4Mux_h
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__6874\ : Odrv4
    port map (
            O => \N__31606\,
            I => \b2v_inst5.un12_clk_100khz_6\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__31603\,
            I => \b2v_inst5.count_rst_4_cascade_\
        );

    \I__6872\ : CascadeMux
    port map (
            O => \N__31600\,
            I => \N__31596\
        );

    \I__6871\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31592\
        );

    \I__6870\ : InMux
    port map (
            O => \N__31596\,
            I => \N__31587\
        );

    \I__6869\ : InMux
    port map (
            O => \N__31595\,
            I => \N__31587\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__31592\,
            I => \b2v_inst5.countZ0Z_10\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__31587\,
            I => \b2v_inst5.countZ0Z_10\
        );

    \I__6866\ : InMux
    port map (
            O => \N__31582\,
            I => \N__31576\
        );

    \I__6865\ : InMux
    port map (
            O => \N__31581\,
            I => \N__31576\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__31576\,
            I => \b2v_inst5.un2_count_1_cry_9_THRU_CO\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__31573\,
            I => \b2v_inst5.countZ0Z_10_cascade_\
        );

    \I__6862\ : InMux
    port map (
            O => \N__31570\,
            I => \N__31567\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__31567\,
            I => \b2v_inst5.count_1_10\
        );

    \I__6860\ : CascadeMux
    port map (
            O => \N__31564\,
            I => \N__31561\
        );

    \I__6859\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31557\
        );

    \I__6858\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31552\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__31557\,
            I => \N__31549\
        );

    \I__6856\ : InMux
    port map (
            O => \N__31556\,
            I => \N__31543\
        );

    \I__6855\ : InMux
    port map (
            O => \N__31555\,
            I => \N__31543\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__31552\,
            I => \N__31540\
        );

    \I__6853\ : Span4Mux_s3_h
    port map (
            O => \N__31549\,
            I => \N__31537\
        );

    \I__6852\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31534\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__31543\,
            I => \b2v_inst5.un2_count_1_cry_0\
        );

    \I__6850\ : Odrv12
    port map (
            O => \N__31540\,
            I => \b2v_inst5.un2_count_1_cry_0\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__31537\,
            I => \b2v_inst5.un2_count_1_cry_0\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__31534\,
            I => \b2v_inst5.un2_count_1_cry_0\
        );

    \I__6847\ : InMux
    port map (
            O => \N__31525\,
            I => \N__31514\
        );

    \I__6846\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31511\
        );

    \I__6845\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31502\
        );

    \I__6844\ : InMux
    port map (
            O => \N__31522\,
            I => \N__31502\
        );

    \I__6843\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31502\
        );

    \I__6842\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31502\
        );

    \I__6841\ : InMux
    port map (
            O => \N__31519\,
            I => \N__31495\
        );

    \I__6840\ : InMux
    port map (
            O => \N__31518\,
            I => \N__31495\
        );

    \I__6839\ : InMux
    port map (
            O => \N__31517\,
            I => \N__31495\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__31514\,
            I => \N__31488\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__31511\,
            I => \N__31481\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__31502\,
            I => \N__31481\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__31495\,
            I => \N__31481\
        );

    \I__6834\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31478\
        );

    \I__6833\ : InMux
    port map (
            O => \N__31493\,
            I => \N__31471\
        );

    \I__6832\ : InMux
    port map (
            O => \N__31492\,
            I => \N__31471\
        );

    \I__6831\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31471\
        );

    \I__6830\ : Span4Mux_s3_h
    port map (
            O => \N__31488\,
            I => \N__31466\
        );

    \I__6829\ : Span4Mux_s3_h
    port map (
            O => \N__31481\,
            I => \N__31466\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__31478\,
            I => \b2v_inst5.N_1_i\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__31471\,
            I => \b2v_inst5.N_1_i\
        );

    \I__6826\ : Odrv4
    port map (
            O => \N__31466\,
            I => \b2v_inst5.N_1_i\
        );

    \I__6825\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31456\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__31456\,
            I => \N__31453\
        );

    \I__6823\ : Odrv4
    port map (
            O => \N__31453\,
            I => \b2v_inst5.count_1_0\
        );

    \I__6822\ : InMux
    port map (
            O => \N__31450\,
            I => \bfn_11_4_0_\
        );

    \I__6821\ : InMux
    port map (
            O => \N__31447\,
            I => \b2v_inst5.un2_count_1_cry_9\
        );

    \I__6820\ : InMux
    port map (
            O => \N__31444\,
            I => \N__31440\
        );

    \I__6819\ : InMux
    port map (
            O => \N__31443\,
            I => \N__31437\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__31440\,
            I => \N__31432\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__31437\,
            I => \N__31432\
        );

    \I__6816\ : Odrv12
    port map (
            O => \N__31432\,
            I => \b2v_inst5.count_rst_3\
        );

    \I__6815\ : InMux
    port map (
            O => \N__31429\,
            I => \b2v_inst5.un2_count_1_cry_10\
        );

    \I__6814\ : InMux
    port map (
            O => \N__31426\,
            I => \N__31422\
        );

    \I__6813\ : InMux
    port map (
            O => \N__31425\,
            I => \N__31419\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__31422\,
            I => \N__31416\
        );

    \I__6811\ : LocalMux
    port map (
            O => \N__31419\,
            I => \b2v_inst5.countZ0Z_12\
        );

    \I__6810\ : Odrv4
    port map (
            O => \N__31416\,
            I => \b2v_inst5.countZ0Z_12\
        );

    \I__6809\ : InMux
    port map (
            O => \N__31411\,
            I => \N__31407\
        );

    \I__6808\ : InMux
    port map (
            O => \N__31410\,
            I => \N__31404\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__31407\,
            I => \N__31401\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__31404\,
            I => \N__31398\
        );

    \I__6805\ : Odrv12
    port map (
            O => \N__31401\,
            I => \b2v_inst5.count_rst_2\
        );

    \I__6804\ : Odrv4
    port map (
            O => \N__31398\,
            I => \b2v_inst5.count_rst_2\
        );

    \I__6803\ : InMux
    port map (
            O => \N__31393\,
            I => \b2v_inst5.un2_count_1_cry_11\
        );

    \I__6802\ : InMux
    port map (
            O => \N__31390\,
            I => \N__31387\
        );

    \I__6801\ : LocalMux
    port map (
            O => \N__31387\,
            I => \N__31383\
        );

    \I__6800\ : InMux
    port map (
            O => \N__31386\,
            I => \N__31380\
        );

    \I__6799\ : Span4Mux_s2_h
    port map (
            O => \N__31383\,
            I => \N__31377\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__31380\,
            I => \b2v_inst5.un2_count_1_axb_13\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__31377\,
            I => \b2v_inst5.un2_count_1_axb_13\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__31372\,
            I => \N__31368\
        );

    \I__6795\ : InMux
    port map (
            O => \N__31371\,
            I => \N__31365\
        );

    \I__6794\ : InMux
    port map (
            O => \N__31368\,
            I => \N__31362\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__31365\,
            I => \N__31357\
        );

    \I__6792\ : LocalMux
    port map (
            O => \N__31362\,
            I => \N__31357\
        );

    \I__6791\ : Span4Mux_v
    port map (
            O => \N__31357\,
            I => \N__31354\
        );

    \I__6790\ : Span4Mux_h
    port map (
            O => \N__31354\,
            I => \N__31351\
        );

    \I__6789\ : Odrv4
    port map (
            O => \N__31351\,
            I => \b2v_inst5.un2_count_1_cry_12_THRU_CO\
        );

    \I__6788\ : InMux
    port map (
            O => \N__31348\,
            I => \b2v_inst5.un2_count_1_cry_12\
        );

    \I__6787\ : CascadeMux
    port map (
            O => \N__31345\,
            I => \N__31342\
        );

    \I__6786\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31338\
        );

    \I__6785\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31335\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__31338\,
            I => \N__31332\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__31335\,
            I => \N__31329\
        );

    \I__6782\ : Odrv4
    port map (
            O => \N__31332\,
            I => \b2v_inst5.countZ0Z_14\
        );

    \I__6781\ : Odrv4
    port map (
            O => \N__31329\,
            I => \b2v_inst5.countZ0Z_14\
        );

    \I__6780\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31320\
        );

    \I__6779\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31317\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__31320\,
            I => \N__31312\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__31317\,
            I => \N__31312\
        );

    \I__6776\ : Span4Mux_h
    port map (
            O => \N__31312\,
            I => \N__31309\
        );

    \I__6775\ : Odrv4
    port map (
            O => \N__31309\,
            I => \b2v_inst5.count_rst_0\
        );

    \I__6774\ : InMux
    port map (
            O => \N__31306\,
            I => \b2v_inst5.un2_count_1_cry_13\
        );

    \I__6773\ : InMux
    port map (
            O => \N__31303\,
            I => \N__31300\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__31300\,
            I => \N__31296\
        );

    \I__6771\ : InMux
    port map (
            O => \N__31299\,
            I => \N__31293\
        );

    \I__6770\ : Odrv12
    port map (
            O => \N__31296\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__6769\ : LocalMux
    port map (
            O => \N__31293\,
            I => \b2v_inst5.countZ0Z_15\
        );

    \I__6768\ : InMux
    port map (
            O => \N__31288\,
            I => \b2v_inst5.un2_count_1_cry_14\
        );

    \I__6767\ : InMux
    port map (
            O => \N__31285\,
            I => \N__31282\
        );

    \I__6766\ : LocalMux
    port map (
            O => \N__31282\,
            I => \N__31279\
        );

    \I__6765\ : Span4Mux_h
    port map (
            O => \N__31279\,
            I => \N__31275\
        );

    \I__6764\ : InMux
    port map (
            O => \N__31278\,
            I => \N__31272\
        );

    \I__6763\ : Odrv4
    port map (
            O => \N__31275\,
            I => \b2v_inst5.count_rst\
        );

    \I__6762\ : LocalMux
    port map (
            O => \N__31272\,
            I => \b2v_inst5.count_rst\
        );

    \I__6761\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31261\
        );

    \I__6759\ : Span4Mux_h
    port map (
            O => \N__31261\,
            I => \N__31258\
        );

    \I__6758\ : Odrv4
    port map (
            O => \N__31258\,
            I => \b2v_inst5.count_1_15\
        );

    \I__6757\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31252\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__31252\,
            I => \N__31247\
        );

    \I__6755\ : InMux
    port map (
            O => \N__31251\,
            I => \N__31244\
        );

    \I__6754\ : InMux
    port map (
            O => \N__31250\,
            I => \N__31241\
        );

    \I__6753\ : Span4Mux_s2_h
    port map (
            O => \N__31247\,
            I => \N__31238\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__31244\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__6751\ : LocalMux
    port map (
            O => \N__31241\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__6750\ : Odrv4
    port map (
            O => \N__31238\,
            I => \b2v_inst5.countZ0Z_1\
        );

    \I__6749\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31228\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__31228\,
            I => \N__31225\
        );

    \I__6747\ : Span4Mux_s3_v
    port map (
            O => \N__31225\,
            I => \N__31222\
        );

    \I__6746\ : Odrv4
    port map (
            O => \N__31222\,
            I => \b2v_inst5.un2_count_1_axb_2\
        );

    \I__6745\ : CascadeMux
    port map (
            O => \N__31219\,
            I => \N__31216\
        );

    \I__6744\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31207\
        );

    \I__6743\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31207\
        );

    \I__6742\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31207\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__31207\,
            I => \N__31204\
        );

    \I__6740\ : Span4Mux_h
    port map (
            O => \N__31204\,
            I => \N__31201\
        );

    \I__6739\ : Odrv4
    port map (
            O => \N__31201\,
            I => \b2v_inst5.count_rst_12\
        );

    \I__6738\ : InMux
    port map (
            O => \N__31198\,
            I => \b2v_inst5.un2_count_1_cry_1\
        );

    \I__6737\ : InMux
    port map (
            O => \N__31195\,
            I => \N__31192\
        );

    \I__6736\ : LocalMux
    port map (
            O => \N__31192\,
            I => \N__31188\
        );

    \I__6735\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31185\
        );

    \I__6734\ : Span4Mux_s2_h
    port map (
            O => \N__31188\,
            I => \N__31182\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__31185\,
            I => \b2v_inst5.countZ0Z_3\
        );

    \I__6732\ : Odrv4
    port map (
            O => \N__31182\,
            I => \b2v_inst5.countZ0Z_3\
        );

    \I__6731\ : CascadeMux
    port map (
            O => \N__31177\,
            I => \N__31173\
        );

    \I__6730\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31168\
        );

    \I__6729\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31168\
        );

    \I__6728\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31165\
        );

    \I__6727\ : Span4Mux_h
    port map (
            O => \N__31165\,
            I => \N__31162\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__31162\,
            I => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\
        );

    \I__6725\ : InMux
    port map (
            O => \N__31159\,
            I => \b2v_inst5.un2_count_1_cry_2\
        );

    \I__6724\ : InMux
    port map (
            O => \N__31156\,
            I => \N__31153\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__31153\,
            I => \N__31149\
        );

    \I__6722\ : CascadeMux
    port map (
            O => \N__31152\,
            I => \N__31146\
        );

    \I__6721\ : Span4Mux_h
    port map (
            O => \N__31149\,
            I => \N__31143\
        );

    \I__6720\ : InMux
    port map (
            O => \N__31146\,
            I => \N__31140\
        );

    \I__6719\ : Span4Mux_v
    port map (
            O => \N__31143\,
            I => \N__31137\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__31140\,
            I => \b2v_inst5.un2_count_1_axb_4\
        );

    \I__6717\ : Odrv4
    port map (
            O => \N__31137\,
            I => \b2v_inst5.un2_count_1_axb_4\
        );

    \I__6716\ : InMux
    port map (
            O => \N__31132\,
            I => \N__31126\
        );

    \I__6715\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31126\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__31126\,
            I => \N__31123\
        );

    \I__6713\ : Span4Mux_v
    port map (
            O => \N__31123\,
            I => \N__31120\
        );

    \I__6712\ : Span4Mux_h
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__6711\ : Odrv4
    port map (
            O => \N__31117\,
            I => \b2v_inst5.un2_count_1_cry_3_THRU_CO\
        );

    \I__6710\ : InMux
    port map (
            O => \N__31114\,
            I => \b2v_inst5.un2_count_1_cry_3\
        );

    \I__6709\ : InMux
    port map (
            O => \N__31111\,
            I => \b2v_inst5.un2_count_1_cry_4\
        );

    \I__6708\ : InMux
    port map (
            O => \N__31108\,
            I => \b2v_inst5.un2_count_1_cry_5\
        );

    \I__6707\ : InMux
    port map (
            O => \N__31105\,
            I => \b2v_inst5.un2_count_1_cry_6\
        );

    \I__6706\ : CascadeMux
    port map (
            O => \N__31102\,
            I => \N__31098\
        );

    \I__6705\ : InMux
    port map (
            O => \N__31101\,
            I => \N__31095\
        );

    \I__6704\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31092\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31089\
        );

    \I__6702\ : LocalMux
    port map (
            O => \N__31092\,
            I => \N__31086\
        );

    \I__6701\ : Span4Mux_s3_v
    port map (
            O => \N__31089\,
            I => \N__31082\
        );

    \I__6700\ : Span4Mux_v
    port map (
            O => \N__31086\,
            I => \N__31079\
        );

    \I__6699\ : InMux
    port map (
            O => \N__31085\,
            I => \N__31076\
        );

    \I__6698\ : Span4Mux_h
    port map (
            O => \N__31082\,
            I => \N__31073\
        );

    \I__6697\ : Odrv4
    port map (
            O => \N__31079\,
            I => \b2v_inst5.countZ0Z_8\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__31076\,
            I => \b2v_inst5.countZ0Z_8\
        );

    \I__6695\ : Odrv4
    port map (
            O => \N__31073\,
            I => \b2v_inst5.countZ0Z_8\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__31066\,
            I => \N__31063\
        );

    \I__6693\ : InMux
    port map (
            O => \N__31063\,
            I => \N__31060\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__31060\,
            I => \N__31056\
        );

    \I__6691\ : InMux
    port map (
            O => \N__31059\,
            I => \N__31053\
        );

    \I__6690\ : Span4Mux_v
    port map (
            O => \N__31056\,
            I => \N__31048\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__31053\,
            I => \N__31048\
        );

    \I__6688\ : Span4Mux_h
    port map (
            O => \N__31048\,
            I => \N__31045\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__31045\,
            I => \b2v_inst5.un2_count_1_cry_7_THRU_CO\
        );

    \I__6686\ : InMux
    port map (
            O => \N__31042\,
            I => \b2v_inst5.un2_count_1_cry_7\
        );

    \I__6685\ : InMux
    port map (
            O => \N__31039\,
            I => \N__31033\
        );

    \I__6684\ : InMux
    port map (
            O => \N__31038\,
            I => \N__31033\
        );

    \I__6683\ : LocalMux
    port map (
            O => \N__31033\,
            I => \N__31030\
        );

    \I__6682\ : Span4Mux_s2_h
    port map (
            O => \N__31030\,
            I => \N__31027\
        );

    \I__6681\ : Odrv4
    port map (
            O => \N__31027\,
            I => \b2v_inst36.un2_count_1_cry_4_THRU_CO\
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__31024\,
            I => \b2v_inst36.countZ0Z_5_cascade_\
        );

    \I__6679\ : InMux
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__31018\,
            I => \b2v_inst36.count_2_5\
        );

    \I__6677\ : InMux
    port map (
            O => \N__31015\,
            I => \N__31010\
        );

    \I__6676\ : InMux
    port map (
            O => \N__31014\,
            I => \N__31005\
        );

    \I__6675\ : InMux
    port map (
            O => \N__31013\,
            I => \N__31005\
        );

    \I__6674\ : LocalMux
    port map (
            O => \N__31010\,
            I => \N__30999\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__31005\,
            I => \N__30999\
        );

    \I__6672\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30996\
        );

    \I__6671\ : Span4Mux_s3_h
    port map (
            O => \N__30999\,
            I => \N__30993\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__30996\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__30993\,
            I => \b2v_inst36.countZ0Z_7\
        );

    \I__6668\ : CascadeMux
    port map (
            O => \N__30988\,
            I => \N__30982\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30987\,
            I => \N__30970\
        );

    \I__6666\ : InMux
    port map (
            O => \N__30986\,
            I => \N__30961\
        );

    \I__6665\ : InMux
    port map (
            O => \N__30985\,
            I => \N__30961\
        );

    \I__6664\ : InMux
    port map (
            O => \N__30982\,
            I => \N__30961\
        );

    \I__6663\ : InMux
    port map (
            O => \N__30981\,
            I => \N__30961\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__30980\,
            I => \N__30953\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30979\,
            I => \N__30945\
        );

    \I__6660\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30945\
        );

    \I__6659\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30938\
        );

    \I__6658\ : InMux
    port map (
            O => \N__30976\,
            I => \N__30938\
        );

    \I__6657\ : InMux
    port map (
            O => \N__30975\,
            I => \N__30938\
        );

    \I__6656\ : InMux
    port map (
            O => \N__30974\,
            I => \N__30933\
        );

    \I__6655\ : InMux
    port map (
            O => \N__30973\,
            I => \N__30933\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__30970\,
            I => \N__30928\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30928\
        );

    \I__6652\ : CascadeMux
    port map (
            O => \N__30960\,
            I => \N__30924\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30959\,
            I => \N__30917\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30958\,
            I => \N__30917\
        );

    \I__6649\ : InMux
    port map (
            O => \N__30957\,
            I => \N__30917\
        );

    \I__6648\ : CascadeMux
    port map (
            O => \N__30956\,
            I => \N__30913\
        );

    \I__6647\ : InMux
    port map (
            O => \N__30953\,
            I => \N__30909\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30952\,
            I => \N__30902\
        );

    \I__6645\ : InMux
    port map (
            O => \N__30951\,
            I => \N__30902\
        );

    \I__6644\ : InMux
    port map (
            O => \N__30950\,
            I => \N__30902\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__30945\,
            I => \N__30899\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__30938\,
            I => \N__30892\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30892\
        );

    \I__6640\ : Span4Mux_s3_h
    port map (
            O => \N__30928\,
            I => \N__30892\
        );

    \I__6639\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30887\
        );

    \I__6638\ : InMux
    port map (
            O => \N__30924\,
            I => \N__30887\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__30917\,
            I => \N__30884\
        );

    \I__6636\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30877\
        );

    \I__6635\ : InMux
    port map (
            O => \N__30913\,
            I => \N__30877\
        );

    \I__6634\ : InMux
    port map (
            O => \N__30912\,
            I => \N__30877\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__30909\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__30902\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6631\ : Odrv4
    port map (
            O => \N__30899\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6630\ : Odrv4
    port map (
            O => \N__30892\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6629\ : LocalMux
    port map (
            O => \N__30887\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__30884\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6627\ : LocalMux
    port map (
            O => \N__30877\,
            I => \b2v_inst36.N_2942_i\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__30862\,
            I => \N__30849\
        );

    \I__6625\ : CascadeMux
    port map (
            O => \N__30861\,
            I => \N__30846\
        );

    \I__6624\ : InMux
    port map (
            O => \N__30860\,
            I => \N__30835\
        );

    \I__6623\ : InMux
    port map (
            O => \N__30859\,
            I => \N__30835\
        );

    \I__6622\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30835\
        );

    \I__6621\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30828\
        );

    \I__6620\ : InMux
    port map (
            O => \N__30856\,
            I => \N__30828\
        );

    \I__6619\ : InMux
    port map (
            O => \N__30855\,
            I => \N__30828\
        );

    \I__6618\ : InMux
    port map (
            O => \N__30854\,
            I => \N__30821\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30853\,
            I => \N__30821\
        );

    \I__6616\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30821\
        );

    \I__6615\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30816\
        );

    \I__6614\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30816\
        );

    \I__6613\ : InMux
    port map (
            O => \N__30845\,
            I => \N__30804\
        );

    \I__6612\ : InMux
    port map (
            O => \N__30844\,
            I => \N__30804\
        );

    \I__6611\ : InMux
    port map (
            O => \N__30843\,
            I => \N__30804\
        );

    \I__6610\ : InMux
    port map (
            O => \N__30842\,
            I => \N__30801\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__30835\,
            I => \N__30796\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__30828\,
            I => \N__30796\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__30821\,
            I => \N__30791\
        );

    \I__6606\ : LocalMux
    port map (
            O => \N__30816\,
            I => \N__30791\
        );

    \I__6605\ : InMux
    port map (
            O => \N__30815\,
            I => \N__30780\
        );

    \I__6604\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30780\
        );

    \I__6603\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30780\
        );

    \I__6602\ : InMux
    port map (
            O => \N__30812\,
            I => \N__30780\
        );

    \I__6601\ : InMux
    port map (
            O => \N__30811\,
            I => \N__30780\
        );

    \I__6600\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30777\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__30801\,
            I => \b2v_inst36.N_1_i\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__30796\,
            I => \b2v_inst36.N_1_i\
        );

    \I__6597\ : Odrv12
    port map (
            O => \N__30791\,
            I => \b2v_inst36.N_1_i\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__30780\,
            I => \b2v_inst36.N_1_i\
        );

    \I__6595\ : Odrv4
    port map (
            O => \N__30777\,
            I => \b2v_inst36.N_1_i\
        );

    \I__6594\ : InMux
    port map (
            O => \N__30766\,
            I => \N__30762\
        );

    \I__6593\ : InMux
    port map (
            O => \N__30765\,
            I => \N__30759\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__30762\,
            I => \N__30756\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__30759\,
            I => \N__30753\
        );

    \I__6590\ : Span4Mux_s1_h
    port map (
            O => \N__30756\,
            I => \N__30750\
        );

    \I__6589\ : Odrv4
    port map (
            O => \N__30753\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__30750\,
            I => \b2v_inst36.un2_count_1_cry_6_THRU_CO\
        );

    \I__6587\ : InMux
    port map (
            O => \N__30745\,
            I => \N__30742\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__30742\,
            I => \N__30739\
        );

    \I__6585\ : Span4Mux_h
    port map (
            O => \N__30739\,
            I => \N__30736\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__30736\,
            I => \b2v_inst36.count_2_7\
        );

    \I__6583\ : CEMux
    port map (
            O => \N__30733\,
            I => \N__30727\
        );

    \I__6582\ : CEMux
    port map (
            O => \N__30732\,
            I => \N__30721\
        );

    \I__6581\ : CEMux
    port map (
            O => \N__30731\,
            I => \N__30718\
        );

    \I__6580\ : CEMux
    port map (
            O => \N__30730\,
            I => \N__30715\
        );

    \I__6579\ : LocalMux
    port map (
            O => \N__30727\,
            I => \N__30712\
        );

    \I__6578\ : InMux
    port map (
            O => \N__30726\,
            I => \N__30702\
        );

    \I__6577\ : InMux
    port map (
            O => \N__30725\,
            I => \N__30702\
        );

    \I__6576\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30690\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__30721\,
            I => \N__30687\
        );

    \I__6574\ : LocalMux
    port map (
            O => \N__30718\,
            I => \N__30684\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__30715\,
            I => \N__30681\
        );

    \I__6572\ : IoSpan4Mux
    port map (
            O => \N__30712\,
            I => \N__30677\
        );

    \I__6571\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30672\
        );

    \I__6570\ : CEMux
    port map (
            O => \N__30710\,
            I => \N__30672\
        );

    \I__6569\ : InMux
    port map (
            O => \N__30709\,
            I => \N__30665\
        );

    \I__6568\ : InMux
    port map (
            O => \N__30708\,
            I => \N__30665\
        );

    \I__6567\ : InMux
    port map (
            O => \N__30707\,
            I => \N__30665\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__30702\,
            I => \N__30662\
        );

    \I__6565\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30655\
        );

    \I__6564\ : CEMux
    port map (
            O => \N__30700\,
            I => \N__30655\
        );

    \I__6563\ : CEMux
    port map (
            O => \N__30699\,
            I => \N__30644\
        );

    \I__6562\ : InMux
    port map (
            O => \N__30698\,
            I => \N__30644\
        );

    \I__6561\ : InMux
    port map (
            O => \N__30697\,
            I => \N__30644\
        );

    \I__6560\ : InMux
    port map (
            O => \N__30696\,
            I => \N__30644\
        );

    \I__6559\ : InMux
    port map (
            O => \N__30695\,
            I => \N__30644\
        );

    \I__6558\ : InMux
    port map (
            O => \N__30694\,
            I => \N__30639\
        );

    \I__6557\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30639\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30634\
        );

    \I__6555\ : Span4Mux_s2_v
    port map (
            O => \N__30687\,
            I => \N__30634\
        );

    \I__6554\ : Span4Mux_s2_v
    port map (
            O => \N__30684\,
            I => \N__30629\
        );

    \I__6553\ : Span4Mux_s2_v
    port map (
            O => \N__30681\,
            I => \N__30629\
        );

    \I__6552\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30626\
        );

    \I__6551\ : Span4Mux_s0_v
    port map (
            O => \N__30677\,
            I => \N__30617\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__30672\,
            I => \N__30617\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__30665\,
            I => \N__30617\
        );

    \I__6548\ : Span4Mux_s3_h
    port map (
            O => \N__30662\,
            I => \N__30617\
        );

    \I__6547\ : InMux
    port map (
            O => \N__30661\,
            I => \N__30612\
        );

    \I__6546\ : InMux
    port map (
            O => \N__30660\,
            I => \N__30612\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__30655\,
            I => \N__30605\
        );

    \I__6544\ : LocalMux
    port map (
            O => \N__30644\,
            I => \N__30605\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__30639\,
            I => \N__30605\
        );

    \I__6542\ : Odrv4
    port map (
            O => \N__30634\,
            I => \b2v_inst36.count_en\
        );

    \I__6541\ : Odrv4
    port map (
            O => \N__30629\,
            I => \b2v_inst36.count_en\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__30626\,
            I => \b2v_inst36.count_en\
        );

    \I__6539\ : Odrv4
    port map (
            O => \N__30617\,
            I => \b2v_inst36.count_en\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__30612\,
            I => \b2v_inst36.count_en\
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__30605\,
            I => \b2v_inst36.count_en\
        );

    \I__6536\ : SRMux
    port map (
            O => \N__30592\,
            I => \N__30584\
        );

    \I__6535\ : SRMux
    port map (
            O => \N__30591\,
            I => \N__30581\
        );

    \I__6534\ : SRMux
    port map (
            O => \N__30590\,
            I => \N__30577\
        );

    \I__6533\ : SRMux
    port map (
            O => \N__30589\,
            I => \N__30574\
        );

    \I__6532\ : SRMux
    port map (
            O => \N__30588\,
            I => \N__30571\
        );

    \I__6531\ : SRMux
    port map (
            O => \N__30587\,
            I => \N__30568\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__30584\,
            I => \N__30565\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__30581\,
            I => \N__30562\
        );

    \I__6528\ : SRMux
    port map (
            O => \N__30580\,
            I => \N__30559\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__30577\,
            I => \N__30556\
        );

    \I__6526\ : LocalMux
    port map (
            O => \N__30574\,
            I => \N__30553\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__30571\,
            I => \N__30550\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__30568\,
            I => \N__30547\
        );

    \I__6523\ : Span4Mux_s2_v
    port map (
            O => \N__30565\,
            I => \N__30540\
        );

    \I__6522\ : Span4Mux_s2_v
    port map (
            O => \N__30562\,
            I => \N__30540\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__30559\,
            I => \N__30540\
        );

    \I__6520\ : Span4Mux_s3_v
    port map (
            O => \N__30556\,
            I => \N__30537\
        );

    \I__6519\ : Span4Mux_s2_v
    port map (
            O => \N__30553\,
            I => \N__30532\
        );

    \I__6518\ : Span4Mux_h
    port map (
            O => \N__30550\,
            I => \N__30527\
        );

    \I__6517\ : Span4Mux_h
    port map (
            O => \N__30547\,
            I => \N__30527\
        );

    \I__6516\ : Span4Mux_h
    port map (
            O => \N__30540\,
            I => \N__30524\
        );

    \I__6515\ : Span4Mux_v
    port map (
            O => \N__30537\,
            I => \N__30521\
        );

    \I__6514\ : InMux
    port map (
            O => \N__30536\,
            I => \N__30516\
        );

    \I__6513\ : InMux
    port map (
            O => \N__30535\,
            I => \N__30516\
        );

    \I__6512\ : Odrv4
    port map (
            O => \N__30532\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6511\ : Odrv4
    port map (
            O => \N__30527\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6510\ : Odrv4
    port map (
            O => \N__30524\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6509\ : Odrv4
    port map (
            O => \N__30521\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__30516\,
            I => \b2v_inst36.count_0_sqmuxa\
        );

    \I__6507\ : InMux
    port map (
            O => \N__30505\,
            I => \N__30502\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__30502\,
            I => \b2v_inst6.count_0_14\
        );

    \I__6505\ : CascadeMux
    port map (
            O => \N__30499\,
            I => \b2v_inst6.countZ0Z_14_cascade_\
        );

    \I__6504\ : InMux
    port map (
            O => \N__30496\,
            I => \N__30493\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__30493\,
            I => \b2v_inst6.count_0_6\
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__30490\,
            I => \N__30485\
        );

    \I__6501\ : CascadeMux
    port map (
            O => \N__30489\,
            I => \N__30482\
        );

    \I__6500\ : CascadeMux
    port map (
            O => \N__30488\,
            I => \N__30479\
        );

    \I__6499\ : InMux
    port map (
            O => \N__30485\,
            I => \N__30476\
        );

    \I__6498\ : InMux
    port map (
            O => \N__30482\,
            I => \N__30471\
        );

    \I__6497\ : InMux
    port map (
            O => \N__30479\,
            I => \N__30471\
        );

    \I__6496\ : LocalMux
    port map (
            O => \N__30476\,
            I => \b2v_inst11.mult1_un152_sum_i_0_8\
        );

    \I__6495\ : LocalMux
    port map (
            O => \N__30471\,
            I => \b2v_inst11.mult1_un152_sum_i_0_8\
        );

    \I__6494\ : InMux
    port map (
            O => \N__30466\,
            I => \N__30463\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__30463\,
            I => \N__30460\
        );

    \I__6492\ : Span4Mux_s2_v
    port map (
            O => \N__30460\,
            I => \N__30457\
        );

    \I__6491\ : Odrv4
    port map (
            O => \N__30457\,
            I => \b2v_inst5.N_51\
        );

    \I__6490\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30451\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__30451\,
            I => \N__30448\
        );

    \I__6488\ : Span4Mux_h
    port map (
            O => \N__30448\,
            I => \N__30445\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__30445\,
            I => \b2v_inst5.curr_state_0_1\
        );

    \I__6486\ : IoInMux
    port map (
            O => \N__30442\,
            I => \N__30439\
        );

    \I__6485\ : LocalMux
    port map (
            O => \N__30439\,
            I => \N__30433\
        );

    \I__6484\ : InMux
    port map (
            O => \N__30438\,
            I => \N__30430\
        );

    \I__6483\ : InMux
    port map (
            O => \N__30437\,
            I => \N__30427\
        );

    \I__6482\ : InMux
    port map (
            O => \N__30436\,
            I => \N__30424\
        );

    \I__6481\ : Span12Mux_s0_v
    port map (
            O => \N__30433\,
            I => \N__30421\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__30430\,
            I => \N__30416\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__30427\,
            I => \N__30416\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30413\
        );

    \I__6477\ : Odrv12
    port map (
            O => \N__30421\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6476\ : Odrv4
    port map (
            O => \N__30416\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6475\ : Odrv4
    port map (
            O => \N__30413\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6474\ : InMux
    port map (
            O => \N__30406\,
            I => \N__30403\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__30403\,
            I => \N__30400\
        );

    \I__6472\ : Span4Mux_s1_v
    port map (
            O => \N__30400\,
            I => \N__30395\
        );

    \I__6471\ : InMux
    port map (
            O => \N__30399\,
            I => \N__30392\
        );

    \I__6470\ : InMux
    port map (
            O => \N__30398\,
            I => \N__30389\
        );

    \I__6469\ : Odrv4
    port map (
            O => \N__30395\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__6468\ : LocalMux
    port map (
            O => \N__30392\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__30389\,
            I => \b2v_inst36.countZ0Z_2\
        );

    \I__6466\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30379\
        );

    \I__6465\ : LocalMux
    port map (
            O => \N__30379\,
            I => \N__30376\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__30376\,
            I => \N__30373\
        );

    \I__6463\ : Odrv4
    port map (
            O => \N__30373\,
            I => \b2v_inst36.un12_clk_100khz_11\
        );

    \I__6462\ : CascadeMux
    port map (
            O => \N__30370\,
            I => \b2v_inst36.count_rst_11_cascade_\
        );

    \I__6461\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30360\
        );

    \I__6460\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30360\
        );

    \I__6459\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30357\
        );

    \I__6458\ : LocalMux
    port map (
            O => \N__30360\,
            I => \N__30352\
        );

    \I__6457\ : LocalMux
    port map (
            O => \N__30357\,
            I => \N__30352\
        );

    \I__6456\ : Odrv4
    port map (
            O => \N__30352\,
            I => \b2v_inst36.countZ0Z_3\
        );

    \I__6455\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30343\
        );

    \I__6454\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30343\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__30343\,
            I => \N__30340\
        );

    \I__6452\ : Odrv4
    port map (
            O => \N__30340\,
            I => \b2v_inst36.un2_count_1_cry_2_THRU_CO\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \b2v_inst36.countZ0Z_3_cascade_\
        );

    \I__6450\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30331\
        );

    \I__6449\ : LocalMux
    port map (
            O => \N__30331\,
            I => \b2v_inst36.count_2_3\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__30328\,
            I => \b2v_inst36.count_rst_9_cascade_\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__30325\,
            I => \N__30322\
        );

    \I__6446\ : InMux
    port map (
            O => \N__30322\,
            I => \N__30317\
        );

    \I__6445\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30314\
        );

    \I__6444\ : InMux
    port map (
            O => \N__30320\,
            I => \N__30311\
        );

    \I__6443\ : LocalMux
    port map (
            O => \N__30317\,
            I => \N__30308\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__30314\,
            I => \N__30305\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__30311\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__6440\ : Odrv4
    port map (
            O => \N__30308\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__6439\ : Odrv4
    port map (
            O => \N__30305\,
            I => \b2v_inst36.countZ0Z_5\
        );

    \I__6438\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30292\
        );

    \I__6437\ : CascadeMux
    port map (
            O => \N__30297\,
            I => \N__30288\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__30296\,
            I => \N__30284\
        );

    \I__6435\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30280\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30275\
        );

    \I__6433\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30272\
        );

    \I__6432\ : InMux
    port map (
            O => \N__30288\,
            I => \N__30269\
        );

    \I__6431\ : InMux
    port map (
            O => \N__30287\,
            I => \N__30266\
        );

    \I__6430\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30261\
        );

    \I__6429\ : InMux
    port map (
            O => \N__30283\,
            I => \N__30261\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__30280\,
            I => \N__30258\
        );

    \I__6427\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30255\
        );

    \I__6426\ : CascadeMux
    port map (
            O => \N__30278\,
            I => \N__30252\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__30275\,
            I => \N__30249\
        );

    \I__6424\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30246\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__30269\,
            I => \N__30243\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__30266\,
            I => \N__30238\
        );

    \I__6421\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30235\
        );

    \I__6420\ : Span4Mux_s2_h
    port map (
            O => \N__30258\,
            I => \N__30230\
        );

    \I__6419\ : LocalMux
    port map (
            O => \N__30255\,
            I => \N__30230\
        );

    \I__6418\ : InMux
    port map (
            O => \N__30252\,
            I => \N__30227\
        );

    \I__6417\ : Span4Mux_v
    port map (
            O => \N__30249\,
            I => \N__30224\
        );

    \I__6416\ : Span4Mux_v
    port map (
            O => \N__30246\,
            I => \N__30219\
        );

    \I__6415\ : Span4Mux_v
    port map (
            O => \N__30243\,
            I => \N__30219\
        );

    \I__6414\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30216\
        );

    \I__6413\ : InMux
    port map (
            O => \N__30241\,
            I => \N__30213\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__30238\,
            I => \N__30206\
        );

    \I__6411\ : Span4Mux_h
    port map (
            O => \N__30235\,
            I => \N__30206\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__30230\,
            I => \N__30206\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__30227\,
            I => \N__30203\
        );

    \I__6408\ : Odrv4
    port map (
            O => \N__30224\,
            I => \dutycycle_RNIU8G3G_0_2\
        );

    \I__6407\ : Odrv4
    port map (
            O => \N__30219\,
            I => \dutycycle_RNIU8G3G_0_2\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__30216\,
            I => \dutycycle_RNIU8G3G_0_2\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__30213\,
            I => \dutycycle_RNIU8G3G_0_2\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__30206\,
            I => \dutycycle_RNIU8G3G_0_2\
        );

    \I__6403\ : Odrv4
    port map (
            O => \N__30203\,
            I => \dutycycle_RNIU8G3G_0_2\
        );

    \I__6402\ : InMux
    port map (
            O => \N__30190\,
            I => \N__30187\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__30187\,
            I => \b2v_inst11.mult1_un152_sum_i\
        );

    \I__6400\ : InMux
    port map (
            O => \N__30184\,
            I => \b2v_inst11.mult1_un159_sum_cry_1\
        );

    \I__6399\ : InMux
    port map (
            O => \N__30181\,
            I => \N__30178\
        );

    \I__6398\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30175\
        );

    \I__6397\ : Span12Mux_s6_h
    port map (
            O => \N__30175\,
            I => \N__30172\
        );

    \I__6396\ : Odrv12
    port map (
            O => \N__30172\,
            I => \b2v_inst11.mult1_un152_sum_cry_3_s\
        );

    \I__6395\ : InMux
    port map (
            O => \N__30169\,
            I => \b2v_inst11.mult1_un159_sum_cry_2\
        );

    \I__6394\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30163\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__6392\ : Span4Mux_s2_v
    port map (
            O => \N__30160\,
            I => \N__30157\
        );

    \I__6391\ : Span4Mux_v
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__30154\,
            I => \N__30151\
        );

    \I__6389\ : Odrv4
    port map (
            O => \N__30151\,
            I => \b2v_inst11.mult1_un152_sum_cry_4_s\
        );

    \I__6388\ : InMux
    port map (
            O => \N__30148\,
            I => \b2v_inst11.mult1_un159_sum_cry_3\
        );

    \I__6387\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30142\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__30142\,
            I => \N__30139\
        );

    \I__6385\ : Span4Mux_s2_v
    port map (
            O => \N__30139\,
            I => \N__30136\
        );

    \I__6384\ : Span4Mux_v
    port map (
            O => \N__30136\,
            I => \N__30133\
        );

    \I__6383\ : Span4Mux_v
    port map (
            O => \N__30133\,
            I => \N__30130\
        );

    \I__6382\ : Odrv4
    port map (
            O => \N__30130\,
            I => \b2v_inst11.mult1_un152_sum_cry_5_s\
        );

    \I__6381\ : InMux
    port map (
            O => \N__30127\,
            I => \b2v_inst11.mult1_un159_sum_cry_4\
        );

    \I__6380\ : InMux
    port map (
            O => \N__30124\,
            I => \N__30121\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__30121\,
            I => \N__30118\
        );

    \I__6378\ : Span4Mux_s2_v
    port map (
            O => \N__30118\,
            I => \N__30115\
        );

    \I__6377\ : Span4Mux_v
    port map (
            O => \N__30115\,
            I => \N__30112\
        );

    \I__6376\ : Span4Mux_v
    port map (
            O => \N__30112\,
            I => \N__30109\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__30109\,
            I => \b2v_inst11.mult1_un152_sum_cry_6_s\
        );

    \I__6374\ : InMux
    port map (
            O => \N__30106\,
            I => \b2v_inst11.mult1_un159_sum_cry_5\
        );

    \I__6373\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30100\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__30100\,
            I => \N__30097\
        );

    \I__6371\ : Span12Mux_s10_v
    port map (
            O => \N__30097\,
            I => \N__30094\
        );

    \I__6370\ : Odrv12
    port map (
            O => \N__30094\,
            I => \b2v_inst11.mult1_un159_sum_axb_7\
        );

    \I__6369\ : InMux
    port map (
            O => \N__30091\,
            I => \b2v_inst11.mult1_un159_sum_cry_6\
        );

    \I__6368\ : InMux
    port map (
            O => \N__30088\,
            I => \N__30083\
        );

    \I__6367\ : InMux
    port map (
            O => \N__30087\,
            I => \N__30080\
        );

    \I__6366\ : InMux
    port map (
            O => \N__30086\,
            I => \N__30077\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__30083\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__30080\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__6363\ : LocalMux
    port map (
            O => \N__30077\,
            I => \b2v_inst11.mult1_un47_sum_s_6\
        );

    \I__6362\ : CascadeMux
    port map (
            O => \N__30070\,
            I => \N__30067\
        );

    \I__6361\ : InMux
    port map (
            O => \N__30067\,
            I => \N__30064\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__30064\,
            I => \b2v_inst11.mult1_un47_sum_l_fx_6\
        );

    \I__6359\ : InMux
    port map (
            O => \N__30061\,
            I => \b2v_inst11.mult1_un54_sum_cry_6\
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__30058\,
            I => \N__30055\
        );

    \I__6357\ : InMux
    port map (
            O => \N__30055\,
            I => \N__30051\
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__30054\,
            I => \N__30048\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__30051\,
            I => \N__30045\
        );

    \I__6354\ : InMux
    port map (
            O => \N__30048\,
            I => \N__30042\
        );

    \I__6353\ : Odrv4
    port map (
            O => \N__30045\,
            I => \b2v_inst11.mult1_un40_sum_i_5\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__30042\,
            I => \b2v_inst11.mult1_un40_sum_i_5\
        );

    \I__6351\ : InMux
    port map (
            O => \N__30037\,
            I => \b2v_inst11.mult1_un54_sum_cry_7\
        );

    \I__6350\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30031\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__30031\,
            I => \b2v_inst11.mult1_un47_sum_l_fx_3\
        );

    \I__6348\ : CascadeMux
    port map (
            O => \N__30028\,
            I => \N__30025\
        );

    \I__6347\ : InMux
    port map (
            O => \N__30025\,
            I => \N__30021\
        );

    \I__6346\ : InMux
    port map (
            O => \N__30024\,
            I => \N__30018\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__30021\,
            I => \N__30015\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__30018\,
            I => \b2v_inst11.mult1_un47_sum\
        );

    \I__6343\ : Odrv12
    port map (
            O => \N__30015\,
            I => \b2v_inst11.mult1_un47_sum\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__30010\,
            I => \N__30007\
        );

    \I__6341\ : InMux
    port map (
            O => \N__30007\,
            I => \N__30000\
        );

    \I__6340\ : InMux
    port map (
            O => \N__30006\,
            I => \N__30000\
        );

    \I__6339\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29997\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__30000\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__29997\,
            I => \b2v_inst11.mult1_un47_sum_cry_3_s\
        );

    \I__6336\ : InMux
    port map (
            O => \N__29992\,
            I => \b2v_inst11.mult1_un47_sum_cry_2\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__29989\,
            I => \N__29986\
        );

    \I__6334\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29983\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__29983\,
            I => \N__29980\
        );

    \I__6332\ : Odrv4
    port map (
            O => \N__29980\,
            I => \b2v_inst11.mult1_un47_sum_s_4_sf\
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__29977\,
            I => \N__29974\
        );

    \I__6330\ : InMux
    port map (
            O => \N__29974\,
            I => \N__29971\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__29971\,
            I => \b2v_inst11.mult1_un47_sum_cry_4_s\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29968\,
            I => \b2v_inst11.mult1_un47_sum_cry_3\
        );

    \I__6327\ : CascadeMux
    port map (
            O => \N__29965\,
            I => \N__29962\
        );

    \I__6326\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29959\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__29959\,
            I => \N__29956\
        );

    \I__6324\ : Odrv4
    port map (
            O => \N__29956\,
            I => \b2v_inst11.mult1_un40_sum_i_l_ofx_4\
        );

    \I__6323\ : CascadeMux
    port map (
            O => \N__29953\,
            I => \N__29950\
        );

    \I__6322\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29947\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__29947\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_s\
        );

    \I__6320\ : InMux
    port map (
            O => \N__29944\,
            I => \b2v_inst11.mult1_un47_sum_cry_4\
        );

    \I__6319\ : InMux
    port map (
            O => \N__29941\,
            I => \b2v_inst11.mult1_un47_sum_cry_5\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29934\
        );

    \I__6317\ : InMux
    port map (
            O => \N__29937\,
            I => \N__29931\
        );

    \I__6316\ : LocalMux
    port map (
            O => \N__29934\,
            I => \N__29928\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__29931\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__6314\ : Odrv4
    port map (
            O => \N__29928\,
            I => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\
        );

    \I__6313\ : CascadeMux
    port map (
            O => \N__29923\,
            I => \N__29917\
        );

    \I__6312\ : InMux
    port map (
            O => \N__29922\,
            I => \N__29914\
        );

    \I__6311\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29911\
        );

    \I__6310\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29906\
        );

    \I__6309\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29906\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__29914\,
            I => \N__29901\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__29911\,
            I => \N__29901\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__29906\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\
        );

    \I__6305\ : Odrv12
    port map (
            O => \N__29901\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__29896\,
            I => \N__29893\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29893\,
            I => \N__29890\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__29890\,
            I => \b2v_inst11.un1_dutycycle_53_i_29\
        );

    \I__6301\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29884\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29884\,
            I => \N__29880\
        );

    \I__6299\ : CascadeMux
    port map (
            O => \N__29883\,
            I => \N__29871\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29868\
        );

    \I__6297\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29863\
        );

    \I__6296\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29863\
        );

    \I__6295\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29856\
        );

    \I__6294\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29856\
        );

    \I__6293\ : InMux
    port map (
            O => \N__29875\,
            I => \N__29856\
        );

    \I__6292\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29851\
        );

    \I__6291\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29851\
        );

    \I__6290\ : Span4Mux_s3_h
    port map (
            O => \N__29868\,
            I => \N__29846\
        );

    \I__6289\ : LocalMux
    port map (
            O => \N__29863\,
            I => \N__29846\
        );

    \I__6288\ : LocalMux
    port map (
            O => \N__29856\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__29851\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__29846\,
            I => \b2v_inst11.curr_stateZ0Z_0\
        );

    \I__6285\ : InMux
    port map (
            O => \N__29839\,
            I => \N__29833\
        );

    \I__6284\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29829\
        );

    \I__6283\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29824\
        );

    \I__6282\ : InMux
    port map (
            O => \N__29836\,
            I => \N__29824\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__29833\,
            I => \N__29821\
        );

    \I__6280\ : InMux
    port map (
            O => \N__29832\,
            I => \N__29818\
        );

    \I__6279\ : LocalMux
    port map (
            O => \N__29829\,
            I => \N__29813\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__29824\,
            I => \N__29813\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__29821\,
            I => \b2v_inst11.count_RNIZ0Z_13\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__29818\,
            I => \b2v_inst11.count_RNIZ0Z_13\
        );

    \I__6275\ : Odrv4
    port map (
            O => \N__29813\,
            I => \b2v_inst11.count_RNIZ0Z_13\
        );

    \I__6274\ : InMux
    port map (
            O => \N__29806\,
            I => \N__29803\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__29803\,
            I => \N__29800\
        );

    \I__6272\ : Span4Mux_s3_v
    port map (
            O => \N__29800\,
            I => \N__29797\
        );

    \I__6271\ : Odrv4
    port map (
            O => \N__29797\,
            I => \b2v_inst11.curr_state_4_0\
        );

    \I__6270\ : CascadeMux
    port map (
            O => \N__29794\,
            I => \N__29790\
        );

    \I__6269\ : InMux
    port map (
            O => \N__29793\,
            I => \N__29787\
        );

    \I__6268\ : InMux
    port map (
            O => \N__29790\,
            I => \N__29784\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__29787\,
            I => \b2v_inst11.CO2_THRU_CO\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__29784\,
            I => \b2v_inst11.CO2_THRU_CO\
        );

    \I__6265\ : CascadeMux
    port map (
            O => \N__29779\,
            I => \N__29775\
        );

    \I__6264\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29771\
        );

    \I__6263\ : InMux
    port map (
            O => \N__29775\,
            I => \N__29766\
        );

    \I__6262\ : InMux
    port map (
            O => \N__29774\,
            I => \N__29766\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__29771\,
            I => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__29766\,
            I => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\
        );

    \I__6259\ : CascadeMux
    port map (
            O => \N__29761\,
            I => \N__29758\
        );

    \I__6258\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29755\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__29755\,
            I => \N__29752\
        );

    \I__6256\ : Odrv4
    port map (
            O => \N__29752\,
            I => \b2v_inst11.mult1_un47_sum_i\
        );

    \I__6255\ : InMux
    port map (
            O => \N__29749\,
            I => \b2v_inst11.mult1_un54_sum_cry_2\
        );

    \I__6254\ : InMux
    port map (
            O => \N__29746\,
            I => \b2v_inst11.mult1_un54_sum_cry_3\
        );

    \I__6253\ : InMux
    port map (
            O => \N__29743\,
            I => \b2v_inst11.mult1_un54_sum_cry_4\
        );

    \I__6252\ : InMux
    port map (
            O => \N__29740\,
            I => \b2v_inst11.mult1_un54_sum_cry_5\
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__29737\,
            I => \N__29733\
        );

    \I__6250\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29727\
        );

    \I__6249\ : InMux
    port map (
            O => \N__29733\,
            I => \N__29722\
        );

    \I__6248\ : InMux
    port map (
            O => \N__29732\,
            I => \N__29719\
        );

    \I__6247\ : InMux
    port map (
            O => \N__29731\,
            I => \N__29716\
        );

    \I__6246\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29713\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__29727\,
            I => \N__29710\
        );

    \I__6244\ : InMux
    port map (
            O => \N__29726\,
            I => \N__29707\
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__29725\,
            I => \N__29702\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29699\
        );

    \I__6241\ : LocalMux
    port map (
            O => \N__29719\,
            I => \N__29696\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__29716\,
            I => \N__29691\
        );

    \I__6239\ : LocalMux
    port map (
            O => \N__29713\,
            I => \N__29691\
        );

    \I__6238\ : Span4Mux_h
    port map (
            O => \N__29710\,
            I => \N__29688\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__29707\,
            I => \N__29685\
        );

    \I__6236\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29680\
        );

    \I__6235\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29680\
        );

    \I__6234\ : InMux
    port map (
            O => \N__29702\,
            I => \N__29677\
        );

    \I__6233\ : Span4Mux_h
    port map (
            O => \N__29699\,
            I => \N__29670\
        );

    \I__6232\ : Span4Mux_v
    port map (
            O => \N__29696\,
            I => \N__29670\
        );

    \I__6231\ : Span4Mux_v
    port map (
            O => \N__29691\,
            I => \N__29670\
        );

    \I__6230\ : Odrv4
    port map (
            O => \N__29688\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__6229\ : Odrv4
    port map (
            O => \N__29685\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__6228\ : LocalMux
    port map (
            O => \N__29680\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__29677\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__6226\ : Odrv4
    port map (
            O => \N__29670\,
            I => \b2v_inst11.dutycycleZ0Z_12\
        );

    \I__6225\ : CascadeMux
    port map (
            O => \N__29659\,
            I => \N__29656\
        );

    \I__6224\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29653\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__29653\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_13\
        );

    \I__6222\ : InMux
    port map (
            O => \N__29650\,
            I => \b2v_inst11.un1_dutycycle_53_cry_13\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__29647\,
            I => \N__29644\
        );

    \I__6220\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29641\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__29641\,
            I => \N__29638\
        );

    \I__6218\ : Span4Mux_h
    port map (
            O => \N__29638\,
            I => \N__29635\
        );

    \I__6217\ : Span4Mux_v
    port map (
            O => \N__29635\,
            I => \N__29632\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__29632\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_15\
        );

    \I__6215\ : InMux
    port map (
            O => \N__29629\,
            I => \b2v_inst11.un1_dutycycle_53_cry_14\
        );

    \I__6214\ : InMux
    port map (
            O => \N__29626\,
            I => \N__29623\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__29623\,
            I => \N__29620\
        );

    \I__6212\ : Span4Mux_v
    port map (
            O => \N__29620\,
            I => \N__29617\
        );

    \I__6211\ : Odrv4
    port map (
            O => \N__29617\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_14\
        );

    \I__6210\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29609\
        );

    \I__6209\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29604\
        );

    \I__6208\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29601\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__29609\,
            I => \N__29598\
        );

    \I__6206\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29595\
        );

    \I__6205\ : CascadeMux
    port map (
            O => \N__29607\,
            I => \N__29591\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__29604\,
            I => \N__29586\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__29601\,
            I => \N__29583\
        );

    \I__6202\ : Span4Mux_h
    port map (
            O => \N__29598\,
            I => \N__29580\
        );

    \I__6201\ : LocalMux
    port map (
            O => \N__29595\,
            I => \N__29577\
        );

    \I__6200\ : InMux
    port map (
            O => \N__29594\,
            I => \N__29574\
        );

    \I__6199\ : InMux
    port map (
            O => \N__29591\,
            I => \N__29571\
        );

    \I__6198\ : InMux
    port map (
            O => \N__29590\,
            I => \N__29568\
        );

    \I__6197\ : InMux
    port map (
            O => \N__29589\,
            I => \N__29565\
        );

    \I__6196\ : Span4Mux_h
    port map (
            O => \N__29586\,
            I => \N__29560\
        );

    \I__6195\ : Span4Mux_h
    port map (
            O => \N__29583\,
            I => \N__29560\
        );

    \I__6194\ : Odrv4
    port map (
            O => \N__29580\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6193\ : Odrv12
    port map (
            O => \N__29577\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6192\ : LocalMux
    port map (
            O => \N__29574\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__29571\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__29568\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__29565\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__29560\,
            I => \b2v_inst11.dutycycleZ0Z_11\
        );

    \I__6187\ : InMux
    port map (
            O => \N__29545\,
            I => \bfn_9_11_0_\
        );

    \I__6186\ : InMux
    port map (
            O => \N__29542\,
            I => \b2v_inst11.CO2\
        );

    \I__6185\ : CascadeMux
    port map (
            O => \N__29539\,
            I => \N__29527\
        );

    \I__6184\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29519\
        );

    \I__6183\ : InMux
    port map (
            O => \N__29537\,
            I => \N__29519\
        );

    \I__6182\ : CascadeMux
    port map (
            O => \N__29536\,
            I => \N__29513\
        );

    \I__6181\ : CascadeMux
    port map (
            O => \N__29535\,
            I => \N__29510\
        );

    \I__6180\ : InMux
    port map (
            O => \N__29534\,
            I => \N__29506\
        );

    \I__6179\ : InMux
    port map (
            O => \N__29533\,
            I => \N__29503\
        );

    \I__6178\ : CascadeMux
    port map (
            O => \N__29532\,
            I => \N__29500\
        );

    \I__6177\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29495\
        );

    \I__6176\ : CascadeMux
    port map (
            O => \N__29530\,
            I => \N__29492\
        );

    \I__6175\ : InMux
    port map (
            O => \N__29527\,
            I => \N__29483\
        );

    \I__6174\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29483\
        );

    \I__6173\ : InMux
    port map (
            O => \N__29525\,
            I => \N__29483\
        );

    \I__6172\ : InMux
    port map (
            O => \N__29524\,
            I => \N__29479\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__29519\,
            I => \N__29476\
        );

    \I__6170\ : InMux
    port map (
            O => \N__29518\,
            I => \N__29465\
        );

    \I__6169\ : InMux
    port map (
            O => \N__29517\,
            I => \N__29465\
        );

    \I__6168\ : InMux
    port map (
            O => \N__29516\,
            I => \N__29465\
        );

    \I__6167\ : InMux
    port map (
            O => \N__29513\,
            I => \N__29465\
        );

    \I__6166\ : InMux
    port map (
            O => \N__29510\,
            I => \N__29465\
        );

    \I__6165\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29462\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__29506\,
            I => \N__29459\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29456\
        );

    \I__6162\ : InMux
    port map (
            O => \N__29500\,
            I => \N__29449\
        );

    \I__6161\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29449\
        );

    \I__6160\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29449\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__29495\,
            I => \N__29446\
        );

    \I__6158\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29439\
        );

    \I__6157\ : InMux
    port map (
            O => \N__29491\,
            I => \N__29439\
        );

    \I__6156\ : InMux
    port map (
            O => \N__29490\,
            I => \N__29439\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__29483\,
            I => \N__29436\
        );

    \I__6154\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29433\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__29479\,
            I => \N__29426\
        );

    \I__6152\ : Span4Mux_v
    port map (
            O => \N__29476\,
            I => \N__29426\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29426\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29417\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__29459\,
            I => \N__29417\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__29456\,
            I => \N__29417\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__29449\,
            I => \N__29417\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__29446\,
            I => \N__29410\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__29439\,
            I => \N__29410\
        );

    \I__6144\ : Span4Mux_h
    port map (
            O => \N__29436\,
            I => \N__29410\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__29433\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__6142\ : Odrv4
    port map (
            O => \N__29426\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__29417\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__29410\,
            I => \b2v_inst11.dutycycleZ0Z_7\
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__29401\,
            I => \N__29394\
        );

    \I__6138\ : CascadeMux
    port map (
            O => \N__29400\,
            I => \N__29385\
        );

    \I__6137\ : InMux
    port map (
            O => \N__29399\,
            I => \N__29382\
        );

    \I__6136\ : InMux
    port map (
            O => \N__29398\,
            I => \N__29379\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__29397\,
            I => \N__29376\
        );

    \I__6134\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29371\
        );

    \I__6133\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29371\
        );

    \I__6132\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29368\
        );

    \I__6131\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29365\
        );

    \I__6130\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29362\
        );

    \I__6129\ : CascadeMux
    port map (
            O => \N__29389\,
            I => \N__29359\
        );

    \I__6128\ : InMux
    port map (
            O => \N__29388\,
            I => \N__29356\
        );

    \I__6127\ : InMux
    port map (
            O => \N__29385\,
            I => \N__29353\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__29382\,
            I => \N__29348\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__29379\,
            I => \N__29348\
        );

    \I__6124\ : InMux
    port map (
            O => \N__29376\,
            I => \N__29345\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__29371\,
            I => \N__29341\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__29368\,
            I => \N__29334\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__29365\,
            I => \N__29334\
        );

    \I__6120\ : LocalMux
    port map (
            O => \N__29362\,
            I => \N__29334\
        );

    \I__6119\ : InMux
    port map (
            O => \N__29359\,
            I => \N__29331\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__29356\,
            I => \N__29326\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__29353\,
            I => \N__29323\
        );

    \I__6116\ : Span4Mux_h
    port map (
            O => \N__29348\,
            I => \N__29320\
        );

    \I__6115\ : LocalMux
    port map (
            O => \N__29345\,
            I => \N__29317\
        );

    \I__6114\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29314\
        );

    \I__6113\ : Span4Mux_s3_h
    port map (
            O => \N__29341\,
            I => \N__29307\
        );

    \I__6112\ : Span4Mux_v
    port map (
            O => \N__29334\,
            I => \N__29307\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__29331\,
            I => \N__29307\
        );

    \I__6110\ : InMux
    port map (
            O => \N__29330\,
            I => \N__29304\
        );

    \I__6109\ : InMux
    port map (
            O => \N__29329\,
            I => \N__29301\
        );

    \I__6108\ : Span4Mux_h
    port map (
            O => \N__29326\,
            I => \N__29298\
        );

    \I__6107\ : Span12Mux_s4_h
    port map (
            O => \N__29323\,
            I => \N__29295\
        );

    \I__6106\ : Span4Mux_v
    port map (
            O => \N__29320\,
            I => \N__29292\
        );

    \I__6105\ : Span4Mux_h
    port map (
            O => \N__29317\,
            I => \N__29285\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__29314\,
            I => \N__29285\
        );

    \I__6103\ : Span4Mux_h
    port map (
            O => \N__29307\,
            I => \N__29285\
        );

    \I__6102\ : LocalMux
    port map (
            O => \N__29304\,
            I => \dutycycle_RNISSAOS1_0_5\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__29301\,
            I => \dutycycle_RNISSAOS1_0_5\
        );

    \I__6100\ : Odrv4
    port map (
            O => \N__29298\,
            I => \dutycycle_RNISSAOS1_0_5\
        );

    \I__6099\ : Odrv12
    port map (
            O => \N__29295\,
            I => \dutycycle_RNISSAOS1_0_5\
        );

    \I__6098\ : Odrv4
    port map (
            O => \N__29292\,
            I => \dutycycle_RNISSAOS1_0_5\
        );

    \I__6097\ : Odrv4
    port map (
            O => \N__29285\,
            I => \dutycycle_RNISSAOS1_0_5\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__29272\,
            I => \N__29269\
        );

    \I__6095\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29266\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__29266\,
            I => \N__29263\
        );

    \I__6093\ : Odrv4
    port map (
            O => \N__29263\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_1\
        );

    \I__6092\ : InMux
    port map (
            O => \N__29260\,
            I => \N__29257\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__6090\ : Odrv4
    port map (
            O => \N__29254\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_9\
        );

    \I__6089\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29247\
        );

    \I__6088\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29244\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__29247\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__29244\,
            I => \b2v_inst11.mult1_un103_sum\
        );

    \I__6085\ : InMux
    port map (
            O => \N__29239\,
            I => \b2v_inst11.un1_dutycycle_53_cry_5\
        );

    \I__6084\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29233\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29230\
        );

    \I__6082\ : Span4Mux_h
    port map (
            O => \N__29230\,
            I => \N__29227\
        );

    \I__6081\ : Odrv4
    port map (
            O => \N__29227\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_9\
        );

    \I__6080\ : CascadeMux
    port map (
            O => \N__29224\,
            I => \N__29220\
        );

    \I__6079\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29212\
        );

    \I__6078\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29209\
        );

    \I__6077\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29204\
        );

    \I__6076\ : InMux
    port map (
            O => \N__29218\,
            I => \N__29204\
        );

    \I__6075\ : CascadeMux
    port map (
            O => \N__29217\,
            I => \N__29201\
        );

    \I__6074\ : InMux
    port map (
            O => \N__29216\,
            I => \N__29195\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__29215\,
            I => \N__29192\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__29212\,
            I => \N__29186\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__29209\,
            I => \N__29181\
        );

    \I__6070\ : LocalMux
    port map (
            O => \N__29204\,
            I => \N__29181\
        );

    \I__6069\ : InMux
    port map (
            O => \N__29201\,
            I => \N__29178\
        );

    \I__6068\ : InMux
    port map (
            O => \N__29200\,
            I => \N__29173\
        );

    \I__6067\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29173\
        );

    \I__6066\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29170\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__29195\,
            I => \N__29167\
        );

    \I__6064\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29164\
        );

    \I__6063\ : InMux
    port map (
            O => \N__29191\,
            I => \N__29157\
        );

    \I__6062\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29157\
        );

    \I__6061\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29157\
        );

    \I__6060\ : Span4Mux_v
    port map (
            O => \N__29186\,
            I => \N__29152\
        );

    \I__6059\ : Span4Mux_h
    port map (
            O => \N__29181\,
            I => \N__29152\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__29178\,
            I => \N__29143\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__29173\,
            I => \N__29143\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__29170\,
            I => \N__29143\
        );

    \I__6055\ : Span4Mux_h
    port map (
            O => \N__29167\,
            I => \N__29143\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__29164\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__29157\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__29152\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__6051\ : Odrv4
    port map (
            O => \N__29143\,
            I => \b2v_inst11.dutycycleZ0Z_4\
        );

    \I__6050\ : InMux
    port map (
            O => \N__29134\,
            I => \b2v_inst11.un1_dutycycle_53_cry_6\
        );

    \I__6049\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29125\
        );

    \I__6048\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29120\
        );

    \I__6047\ : InMux
    port map (
            O => \N__29129\,
            I => \N__29120\
        );

    \I__6046\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29117\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__29125\,
            I => \N__29112\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__29120\,
            I => \N__29109\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__29117\,
            I => \N__29106\
        );

    \I__6042\ : InMux
    port map (
            O => \N__29116\,
            I => \N__29103\
        );

    \I__6041\ : InMux
    port map (
            O => \N__29115\,
            I => \N__29098\
        );

    \I__6040\ : Span4Mux_h
    port map (
            O => \N__29112\,
            I => \N__29095\
        );

    \I__6039\ : Span4Mux_v
    port map (
            O => \N__29109\,
            I => \N__29088\
        );

    \I__6038\ : Span4Mux_h
    port map (
            O => \N__29106\,
            I => \N__29088\
        );

    \I__6037\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29088\
        );

    \I__6036\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29083\
        );

    \I__6035\ : InMux
    port map (
            O => \N__29101\,
            I => \N__29083\
        );

    \I__6034\ : LocalMux
    port map (
            O => \N__29098\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__6033\ : Odrv4
    port map (
            O => \N__29095\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__6032\ : Odrv4
    port map (
            O => \N__29088\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__29083\,
            I => \b2v_inst11.dutycycleZ0Z_6\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__29074\,
            I => \N__29071\
        );

    \I__6029\ : InMux
    port map (
            O => \N__29071\,
            I => \N__29068\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__29068\,
            I => \N__29065\
        );

    \I__6027\ : Span4Mux_h
    port map (
            O => \N__29065\,
            I => \N__29062\
        );

    \I__6026\ : Odrv4
    port map (
            O => \N__29062\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_11\
        );

    \I__6025\ : InMux
    port map (
            O => \N__29059\,
            I => \bfn_9_10_0_\
        );

    \I__6024\ : InMux
    port map (
            O => \N__29056\,
            I => \N__29053\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__29053\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_12\
        );

    \I__6022\ : InMux
    port map (
            O => \N__29050\,
            I => \N__29041\
        );

    \I__6021\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29041\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__29048\,
            I => \N__29038\
        );

    \I__6019\ : InMux
    port map (
            O => \N__29047\,
            I => \N__29034\
        );

    \I__6018\ : CascadeMux
    port map (
            O => \N__29046\,
            I => \N__29030\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__29041\,
            I => \N__29024\
        );

    \I__6016\ : InMux
    port map (
            O => \N__29038\,
            I => \N__29021\
        );

    \I__6015\ : InMux
    port map (
            O => \N__29037\,
            I => \N__29018\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__29034\,
            I => \N__29015\
        );

    \I__6013\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29012\
        );

    \I__6012\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29009\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__29029\,
            I => \N__29006\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__29028\,
            I => \N__29002\
        );

    \I__6009\ : CascadeMux
    port map (
            O => \N__29027\,
            I => \N__28997\
        );

    \I__6008\ : Span4Mux_v
    port map (
            O => \N__29024\,
            I => \N__28994\
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__29021\,
            I => \N__28989\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__29018\,
            I => \N__28989\
        );

    \I__6005\ : Span4Mux_h
    port map (
            O => \N__29015\,
            I => \N__28986\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__29012\,
            I => \N__28983\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__29009\,
            I => \N__28980\
        );

    \I__6002\ : InMux
    port map (
            O => \N__29006\,
            I => \N__28977\
        );

    \I__6001\ : InMux
    port map (
            O => \N__29005\,
            I => \N__28974\
        );

    \I__6000\ : InMux
    port map (
            O => \N__29002\,
            I => \N__28965\
        );

    \I__5999\ : InMux
    port map (
            O => \N__29001\,
            I => \N__28965\
        );

    \I__5998\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28965\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28997\,
            I => \N__28965\
        );

    \I__5996\ : Span4Mux_h
    port map (
            O => \N__28994\,
            I => \N__28960\
        );

    \I__5995\ : Span4Mux_h
    port map (
            O => \N__28989\,
            I => \N__28960\
        );

    \I__5994\ : Odrv4
    port map (
            O => \N__28986\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5993\ : Odrv4
    port map (
            O => \N__28983\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5992\ : Odrv12
    port map (
            O => \N__28980\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__28977\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__28974\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__28965\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5988\ : Odrv4
    port map (
            O => \N__28960\,
            I => \b2v_inst11.dutycycleZ0Z_9\
        );

    \I__5987\ : InMux
    port map (
            O => \N__28945\,
            I => \b2v_inst11.un1_dutycycle_53_cry_8\
        );

    \I__5986\ : CascadeMux
    port map (
            O => \N__28942\,
            I => \N__28939\
        );

    \I__5985\ : InMux
    port map (
            O => \N__28939\,
            I => \N__28936\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__28936\,
            I => \N__28933\
        );

    \I__5983\ : Span4Mux_v
    port map (
            O => \N__28933\,
            I => \N__28930\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__28930\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_13\
        );

    \I__5981\ : InMux
    port map (
            O => \N__28927\,
            I => \b2v_inst11.un1_dutycycle_53_cry_9\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__28924\,
            I => \N__28921\
        );

    \I__5979\ : InMux
    port map (
            O => \N__28921\,
            I => \N__28918\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__28918\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_14\
        );

    \I__5977\ : InMux
    port map (
            O => \N__28915\,
            I => \b2v_inst11.un1_dutycycle_53_cry_10\
        );

    \I__5976\ : CascadeMux
    port map (
            O => \N__28912\,
            I => \N__28909\
        );

    \I__5975\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28906\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__28906\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_11\
        );

    \I__5973\ : InMux
    port map (
            O => \N__28903\,
            I => \b2v_inst11.un1_dutycycle_53_cry_11\
        );

    \I__5972\ : InMux
    port map (
            O => \N__28900\,
            I => \N__28892\
        );

    \I__5971\ : InMux
    port map (
            O => \N__28899\,
            I => \N__28889\
        );

    \I__5970\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28886\
        );

    \I__5969\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28883\
        );

    \I__5968\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28878\
        );

    \I__5967\ : InMux
    port map (
            O => \N__28895\,
            I => \N__28875\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__28892\,
            I => \N__28872\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__28889\,
            I => \N__28865\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__28886\,
            I => \N__28865\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__28883\,
            I => \N__28865\
        );

    \I__5962\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28860\
        );

    \I__5961\ : InMux
    port map (
            O => \N__28881\,
            I => \N__28860\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__28878\,
            I => \N__28855\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__28875\,
            I => \N__28855\
        );

    \I__5958\ : Odrv12
    port map (
            O => \N__28872\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__5957\ : Odrv4
    port map (
            O => \N__28865\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__28860\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__28855\,
            I => \b2v_inst11.dutycycleZ0Z_8\
        );

    \I__5954\ : CascadeMux
    port map (
            O => \N__28846\,
            I => \N__28843\
        );

    \I__5953\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28840\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__28840\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_13\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28837\,
            I => \b2v_inst11.un1_dutycycle_53_cry_12\
        );

    \I__5950\ : InMux
    port map (
            O => \N__28834\,
            I => \b2v_inst11.mult1_un103_sum_cry_7\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__28831\,
            I => \N__28826\
        );

    \I__5948\ : InMux
    port map (
            O => \N__28830\,
            I => \N__28822\
        );

    \I__5947\ : InMux
    port map (
            O => \N__28829\,
            I => \N__28817\
        );

    \I__5946\ : InMux
    port map (
            O => \N__28826\,
            I => \N__28817\
        );

    \I__5945\ : InMux
    port map (
            O => \N__28825\,
            I => \N__28814\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__28822\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__28817\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__28814\,
            I => \b2v_inst11.mult1_un103_sum_s_8\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__28807\,
            I => \b2v_inst11.mult1_un103_sum_s_8_cascade_\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__28804\,
            I => \N__28800\
        );

    \I__5939\ : CascadeMux
    port map (
            O => \N__28803\,
            I => \N__28796\
        );

    \I__5938\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28789\
        );

    \I__5937\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28789\
        );

    \I__5936\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28789\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__28789\,
            I => \b2v_inst11.mult1_un103_sum_i_0_8\
        );

    \I__5934\ : InMux
    port map (
            O => \N__28786\,
            I => \N__28781\
        );

    \I__5933\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28776\
        );

    \I__5932\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28776\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__28781\,
            I => \N__28769\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__28776\,
            I => \N__28766\
        );

    \I__5929\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28759\
        );

    \I__5928\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28759\
        );

    \I__5927\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28759\
        );

    \I__5926\ : InMux
    port map (
            O => \N__28772\,
            I => \N__28751\
        );

    \I__5925\ : Span4Mux_v
    port map (
            O => \N__28769\,
            I => \N__28744\
        );

    \I__5924\ : Span4Mux_v
    port map (
            O => \N__28766\,
            I => \N__28744\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__28759\,
            I => \N__28744\
        );

    \I__5922\ : CascadeMux
    port map (
            O => \N__28758\,
            I => \N__28741\
        );

    \I__5921\ : CascadeMux
    port map (
            O => \N__28757\,
            I => \N__28738\
        );

    \I__5920\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28735\
        );

    \I__5919\ : InMux
    port map (
            O => \N__28755\,
            I => \N__28730\
        );

    \I__5918\ : InMux
    port map (
            O => \N__28754\,
            I => \N__28730\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__28751\,
            I => \N__28725\
        );

    \I__5916\ : Span4Mux_h
    port map (
            O => \N__28744\,
            I => \N__28725\
        );

    \I__5915\ : InMux
    port map (
            O => \N__28741\,
            I => \N__28722\
        );

    \I__5914\ : InMux
    port map (
            O => \N__28738\,
            I => \N__28719\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__28735\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5912\ : LocalMux
    port map (
            O => \N__28730\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5911\ : Odrv4
    port map (
            O => \N__28725\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__28722\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__28719\,
            I => \b2v_inst11.dutycycleZ0Z_3\
        );

    \I__5908\ : InMux
    port map (
            O => \N__28708\,
            I => \N__28704\
        );

    \I__5907\ : InMux
    port map (
            O => \N__28707\,
            I => \N__28701\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__28704\,
            I => \N__28696\
        );

    \I__5905\ : LocalMux
    port map (
            O => \N__28701\,
            I => \N__28696\
        );

    \I__5904\ : Odrv4
    port map (
            O => \N__28696\,
            I => \b2v_inst11.un1_dutycycle_53_axb_0\
        );

    \I__5903\ : InMux
    port map (
            O => \N__28693\,
            I => \N__28690\
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__28690\,
            I => \N__28687\
        );

    \I__5901\ : Span4Mux_h
    port map (
            O => \N__28687\,
            I => \N__28684\
        );

    \I__5900\ : Odrv4
    port map (
            O => \N__28684\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_1\
        );

    \I__5899\ : InMux
    port map (
            O => \N__28681\,
            I => \N__28678\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__28678\,
            I => \N__28674\
        );

    \I__5897\ : InMux
    port map (
            O => \N__28677\,
            I => \N__28671\
        );

    \I__5896\ : Span4Mux_h
    port map (
            O => \N__28674\,
            I => \N__28666\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__28671\,
            I => \N__28666\
        );

    \I__5894\ : Span4Mux_v
    port map (
            O => \N__28666\,
            I => \N__28663\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__28663\,
            I => \b2v_inst11.mult1_un138_sum\
        );

    \I__5892\ : InMux
    port map (
            O => \N__28660\,
            I => \b2v_inst11.un1_dutycycle_53_cry_0\
        );

    \I__5891\ : InMux
    port map (
            O => \N__28657\,
            I => \N__28653\
        );

    \I__5890\ : InMux
    port map (
            O => \N__28656\,
            I => \N__28650\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__28653\,
            I => \N__28647\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__28650\,
            I => \N__28642\
        );

    \I__5887\ : Span4Mux_h
    port map (
            O => \N__28647\,
            I => \N__28642\
        );

    \I__5886\ : Odrv4
    port map (
            O => \N__28642\,
            I => \b2v_inst11.mult1_un131_sum\
        );

    \I__5885\ : InMux
    port map (
            O => \N__28639\,
            I => \b2v_inst11.un1_dutycycle_53_cry_1\
        );

    \I__5884\ : InMux
    port map (
            O => \N__28636\,
            I => \N__28633\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__28633\,
            I => \N__28630\
        );

    \I__5882\ : Odrv4
    port map (
            O => \N__28630\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_2\
        );

    \I__5881\ : InMux
    port map (
            O => \N__28627\,
            I => \N__28623\
        );

    \I__5880\ : InMux
    port map (
            O => \N__28626\,
            I => \N__28620\
        );

    \I__5879\ : LocalMux
    port map (
            O => \N__28623\,
            I => \N__28615\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__28620\,
            I => \N__28615\
        );

    \I__5877\ : Span4Mux_h
    port map (
            O => \N__28615\,
            I => \N__28612\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__28612\,
            I => \b2v_inst11.mult1_un124_sum\
        );

    \I__5875\ : InMux
    port map (
            O => \N__28609\,
            I => \b2v_inst11.un1_dutycycle_53_cry_2\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__28606\,
            I => \N__28602\
        );

    \I__5873\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28599\
        );

    \I__5872\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28596\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28593\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__28596\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_3\
        );

    \I__5869\ : Odrv4
    port map (
            O => \N__28593\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_3\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__28588\,
            I => \N__28585\
        );

    \I__5867\ : InMux
    port map (
            O => \N__28585\,
            I => \N__28582\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__28582\,
            I => \N__28579\
        );

    \I__5865\ : Odrv4
    port map (
            O => \N__28579\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_3\
        );

    \I__5864\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28572\
        );

    \I__5863\ : InMux
    port map (
            O => \N__28575\,
            I => \N__28569\
        );

    \I__5862\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28564\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__28569\,
            I => \N__28564\
        );

    \I__5860\ : Odrv4
    port map (
            O => \N__28564\,
            I => \b2v_inst11.mult1_un117_sum\
        );

    \I__5859\ : InMux
    port map (
            O => \N__28561\,
            I => \b2v_inst11.un1_dutycycle_53_cry_3\
        );

    \I__5858\ : CascadeMux
    port map (
            O => \N__28558\,
            I => \N__28555\
        );

    \I__5857\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28552\
        );

    \I__5856\ : LocalMux
    port map (
            O => \N__28552\,
            I => \N__28549\
        );

    \I__5855\ : Span4Mux_s3_h
    port map (
            O => \N__28549\,
            I => \N__28546\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__28546\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_8\
        );

    \I__5853\ : InMux
    port map (
            O => \N__28543\,
            I => \N__28539\
        );

    \I__5852\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28536\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28533\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__28536\,
            I => \b2v_inst11.mult1_un110_sum\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__28533\,
            I => \b2v_inst11.mult1_un110_sum\
        );

    \I__5848\ : InMux
    port map (
            O => \N__28528\,
            I => \b2v_inst11.un1_dutycycle_53_cry_4\
        );

    \I__5847\ : CascadeMux
    port map (
            O => \N__28525\,
            I => \N__28522\
        );

    \I__5846\ : InMux
    port map (
            O => \N__28522\,
            I => \N__28519\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__28519\,
            I => \b2v_inst11.mult1_un117_sum_axb_8\
        );

    \I__5844\ : InMux
    port map (
            O => \N__28516\,
            I => \b2v_inst11.mult1_un110_sum_cry_6\
        );

    \I__5843\ : InMux
    port map (
            O => \N__28513\,
            I => \b2v_inst11.mult1_un110_sum_cry_7\
        );

    \I__5842\ : CascadeMux
    port map (
            O => \N__28510\,
            I => \b2v_inst11.mult1_un110_sum_s_8_cascade_\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__28507\,
            I => \N__28503\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__28506\,
            I => \N__28499\
        );

    \I__5839\ : InMux
    port map (
            O => \N__28503\,
            I => \N__28492\
        );

    \I__5838\ : InMux
    port map (
            O => \N__28502\,
            I => \N__28492\
        );

    \I__5837\ : InMux
    port map (
            O => \N__28499\,
            I => \N__28492\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__28492\,
            I => \b2v_inst11.mult1_un110_sum_i_0_8\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__28489\,
            I => \N__28486\
        );

    \I__5834\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28483\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__28483\,
            I => \b2v_inst11.mult1_un103_sum_cry_3_s\
        );

    \I__5832\ : InMux
    port map (
            O => \N__28480\,
            I => \b2v_inst11.mult1_un103_sum_cry_2\
        );

    \I__5831\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28474\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__28474\,
            I => \b2v_inst11.mult1_un103_sum_cry_4_s\
        );

    \I__5829\ : InMux
    port map (
            O => \N__28471\,
            I => \b2v_inst11.mult1_un103_sum_cry_3\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__28468\,
            I => \N__28465\
        );

    \I__5827\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28462\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__28462\,
            I => \b2v_inst11.mult1_un103_sum_cry_5_s\
        );

    \I__5825\ : InMux
    port map (
            O => \N__28459\,
            I => \b2v_inst11.mult1_un103_sum_cry_4\
        );

    \I__5824\ : InMux
    port map (
            O => \N__28456\,
            I => \N__28453\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__28453\,
            I => \b2v_inst11.mult1_un103_sum_cry_6_s\
        );

    \I__5822\ : InMux
    port map (
            O => \N__28450\,
            I => \b2v_inst11.mult1_un103_sum_cry_5\
        );

    \I__5821\ : CascadeMux
    port map (
            O => \N__28447\,
            I => \N__28443\
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__28446\,
            I => \N__28439\
        );

    \I__5819\ : InMux
    port map (
            O => \N__28443\,
            I => \N__28432\
        );

    \I__5818\ : InMux
    port map (
            O => \N__28442\,
            I => \N__28432\
        );

    \I__5817\ : InMux
    port map (
            O => \N__28439\,
            I => \N__28432\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__28432\,
            I => \b2v_inst11.mult1_un96_sum_i_0_8\
        );

    \I__5815\ : CascadeMux
    port map (
            O => \N__28429\,
            I => \N__28426\
        );

    \I__5814\ : InMux
    port map (
            O => \N__28426\,
            I => \N__28423\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__28423\,
            I => \b2v_inst11.mult1_un110_sum_axb_8\
        );

    \I__5812\ : InMux
    port map (
            O => \N__28420\,
            I => \b2v_inst11.mult1_un103_sum_cry_6\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__28417\,
            I => \N__28414\
        );

    \I__5810\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28411\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__28411\,
            I => \b2v_inst11.mult1_un138_sum_cry_6_s\
        );

    \I__5808\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28405\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__28405\,
            I => \N__28402\
        );

    \I__5806\ : Odrv4
    port map (
            O => \N__28402\,
            I => \b2v_inst11.mult1_un152_sum_axb_8\
        );

    \I__5805\ : InMux
    port map (
            O => \N__28399\,
            I => \b2v_inst11.mult1_un145_sum_cry_6\
        );

    \I__5804\ : InMux
    port map (
            O => \N__28396\,
            I => \N__28393\
        );

    \I__5803\ : LocalMux
    port map (
            O => \N__28393\,
            I => \b2v_inst11.mult1_un145_sum_axb_8\
        );

    \I__5802\ : InMux
    port map (
            O => \N__28390\,
            I => \b2v_inst11.mult1_un145_sum_cry_7\
        );

    \I__5801\ : CascadeMux
    port map (
            O => \N__28387\,
            I => \N__28382\
        );

    \I__5800\ : CascadeMux
    port map (
            O => \N__28386\,
            I => \N__28379\
        );

    \I__5799\ : InMux
    port map (
            O => \N__28385\,
            I => \N__28374\
        );

    \I__5798\ : InMux
    port map (
            O => \N__28382\,
            I => \N__28374\
        );

    \I__5797\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28371\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__28374\,
            I => \b2v_inst11.mult1_un138_sum_i_0_8\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__28371\,
            I => \b2v_inst11.mult1_un138_sum_i_0_8\
        );

    \I__5794\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28363\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__28363\,
            I => \b2v_inst11.mult1_un103_sum_i\
        );

    \I__5792\ : CascadeMux
    port map (
            O => \N__28360\,
            I => \N__28357\
        );

    \I__5791\ : InMux
    port map (
            O => \N__28357\,
            I => \N__28354\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__28354\,
            I => \b2v_inst11.mult1_un110_sum_cry_3_s\
        );

    \I__5789\ : InMux
    port map (
            O => \N__28351\,
            I => \b2v_inst11.mult1_un110_sum_cry_2\
        );

    \I__5788\ : InMux
    port map (
            O => \N__28348\,
            I => \N__28345\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__28345\,
            I => \b2v_inst11.mult1_un110_sum_cry_4_s\
        );

    \I__5786\ : InMux
    port map (
            O => \N__28342\,
            I => \b2v_inst11.mult1_un110_sum_cry_3\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__28339\,
            I => \N__28336\
        );

    \I__5784\ : InMux
    port map (
            O => \N__28336\,
            I => \N__28333\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__28333\,
            I => \b2v_inst11.mult1_un110_sum_cry_5_s\
        );

    \I__5782\ : InMux
    port map (
            O => \N__28330\,
            I => \b2v_inst11.mult1_un110_sum_cry_4\
        );

    \I__5781\ : InMux
    port map (
            O => \N__28327\,
            I => \N__28324\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__28324\,
            I => \b2v_inst11.mult1_un110_sum_cry_6_s\
        );

    \I__5779\ : InMux
    port map (
            O => \N__28321\,
            I => \b2v_inst11.mult1_un110_sum_cry_5\
        );

    \I__5778\ : CascadeMux
    port map (
            O => \N__28318\,
            I => \b2v_inst5.un2_count_1_axb_13_cascade_\
        );

    \I__5777\ : InMux
    port map (
            O => \N__28315\,
            I => \N__28312\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__28312\,
            I => \b2v_inst5.count_rst_1\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__28309\,
            I => \N__28306\
        );

    \I__5774\ : InMux
    port map (
            O => \N__28306\,
            I => \N__28302\
        );

    \I__5773\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28299\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__28302\,
            I => \b2v_inst5.count_1_13\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__28299\,
            I => \b2v_inst5.count_1_13\
        );

    \I__5770\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28291\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__28291\,
            I => \N__28288\
        );

    \I__5768\ : Span4Mux_v
    port map (
            O => \N__28288\,
            I => \N__28285\
        );

    \I__5767\ : Odrv4
    port map (
            O => \N__28285\,
            I => \b2v_inst5.un12_clk_100khz_5\
        );

    \I__5766\ : InMux
    port map (
            O => \N__28282\,
            I => \N__28279\
        );

    \I__5765\ : LocalMux
    port map (
            O => \N__28279\,
            I => \N__28276\
        );

    \I__5764\ : Span4Mux_h
    port map (
            O => \N__28276\,
            I => \N__28273\
        );

    \I__5763\ : Odrv4
    port map (
            O => \N__28273\,
            I => \b2v_inst5.count_rst_6\
        );

    \I__5762\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28267\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__28267\,
            I => \N__28264\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__28264\,
            I => \b2v_inst5.un12_clk_100khz_8\
        );

    \I__5759\ : InMux
    port map (
            O => \N__28261\,
            I => \N__28258\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__28258\,
            I => \N__28255\
        );

    \I__5757\ : Span4Mux_v
    port map (
            O => \N__28255\,
            I => \N__28252\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__28252\,
            I => \b2v_inst11.mult1_un138_sum_i\
        );

    \I__5755\ : InMux
    port map (
            O => \N__28249\,
            I => \N__28246\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__28246\,
            I => \N__28243\
        );

    \I__5753\ : Odrv12
    port map (
            O => \N__28243\,
            I => \b2v_inst11.mult1_un145_sum_cry_3_s\
        );

    \I__5752\ : InMux
    port map (
            O => \N__28240\,
            I => \b2v_inst11.mult1_un145_sum_cry_2\
        );

    \I__5751\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__28234\,
            I => \b2v_inst11.mult1_un138_sum_cry_3_s\
        );

    \I__5749\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__28228\,
            I => \N__28225\
        );

    \I__5747\ : Odrv12
    port map (
            O => \N__28225\,
            I => \b2v_inst11.mult1_un145_sum_cry_4_s\
        );

    \I__5746\ : InMux
    port map (
            O => \N__28222\,
            I => \b2v_inst11.mult1_un145_sum_cry_3\
        );

    \I__5745\ : CascadeMux
    port map (
            O => \N__28219\,
            I => \N__28216\
        );

    \I__5744\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__28213\,
            I => \b2v_inst11.mult1_un138_sum_cry_4_s\
        );

    \I__5742\ : InMux
    port map (
            O => \N__28210\,
            I => \N__28207\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__28207\,
            I => \N__28204\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__28204\,
            I => \b2v_inst11.mult1_un145_sum_cry_5_s\
        );

    \I__5739\ : InMux
    port map (
            O => \N__28201\,
            I => \b2v_inst11.mult1_un145_sum_cry_4\
        );

    \I__5738\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28195\
        );

    \I__5737\ : LocalMux
    port map (
            O => \N__28195\,
            I => \b2v_inst11.mult1_un138_sum_cry_5_s\
        );

    \I__5736\ : InMux
    port map (
            O => \N__28192\,
            I => \N__28189\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__28189\,
            I => \N__28186\
        );

    \I__5734\ : Odrv4
    port map (
            O => \N__28186\,
            I => \b2v_inst11.mult1_un145_sum_cry_6_s\
        );

    \I__5733\ : InMux
    port map (
            O => \N__28183\,
            I => \b2v_inst11.mult1_un145_sum_cry_5\
        );

    \I__5732\ : CascadeMux
    port map (
            O => \N__28180\,
            I => \b2v_inst5.count_RNIZ0Z_1_cascade_\
        );

    \I__5731\ : InMux
    port map (
            O => \N__28177\,
            I => \N__28174\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__28174\,
            I => \b2v_inst5.count_1_3\
        );

    \I__5729\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28168\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__28168\,
            I => \b2v_inst5.count_RNIZ0Z_1\
        );

    \I__5727\ : InMux
    port map (
            O => \N__28165\,
            I => \N__28162\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__28162\,
            I => \b2v_inst5.count_1_1\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__28159\,
            I => \b2v_inst5.count_rst_14_cascade_\
        );

    \I__5724\ : CascadeMux
    port map (
            O => \N__28156\,
            I => \b2v_inst5.count_rst_1_cascade_\
        );

    \I__5723\ : CascadeMux
    port map (
            O => \N__28153\,
            I => \b2v_inst36.count_rst_4_cascade_\
        );

    \I__5722\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28146\
        );

    \I__5721\ : CascadeMux
    port map (
            O => \N__28149\,
            I => \N__28143\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__28146\,
            I => \N__28139\
        );

    \I__5719\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28136\
        );

    \I__5718\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28133\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__28139\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__28136\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__28133\,
            I => \b2v_inst36.countZ0Z_10\
        );

    \I__5714\ : InMux
    port map (
            O => \N__28126\,
            I => \N__28120\
        );

    \I__5713\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28120\
        );

    \I__5712\ : LocalMux
    port map (
            O => \N__28120\,
            I => \b2v_inst36.un2_count_1_cry_9_THRU_CO\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__28117\,
            I => \b2v_inst36.countZ0Z_10_cascade_\
        );

    \I__5710\ : InMux
    port map (
            O => \N__28114\,
            I => \N__28111\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__28111\,
            I => \b2v_inst36.count_2_10\
        );

    \I__5708\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28104\
        );

    \I__5707\ : InMux
    port map (
            O => \N__28107\,
            I => \N__28101\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__28104\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__28101\,
            I => \b2v_inst36.countZ0Z_13\
        );

    \I__5704\ : InMux
    port map (
            O => \N__28096\,
            I => \N__28090\
        );

    \I__5703\ : InMux
    port map (
            O => \N__28095\,
            I => \N__28090\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__28090\,
            I => \b2v_inst36.count_rst_1\
        );

    \I__5701\ : InMux
    port map (
            O => \N__28087\,
            I => \N__28084\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__28084\,
            I => \b2v_inst36.count_2_13\
        );

    \I__5699\ : InMux
    port map (
            O => \N__28081\,
            I => \N__28078\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__28078\,
            I => \N__28075\
        );

    \I__5697\ : Odrv12
    port map (
            O => \N__28075\,
            I => \b2v_inst36.count_2_15\
        );

    \I__5696\ : InMux
    port map (
            O => \N__28072\,
            I => \N__28068\
        );

    \I__5695\ : InMux
    port map (
            O => \N__28071\,
            I => \N__28065\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__28068\,
            I => \b2v_inst36.count_rst\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__28065\,
            I => \b2v_inst36.count_rst\
        );

    \I__5692\ : InMux
    port map (
            O => \N__28060\,
            I => \N__28056\
        );

    \I__5691\ : InMux
    port map (
            O => \N__28059\,
            I => \N__28053\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__28056\,
            I => \b2v_inst36.countZ0Z_15\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__28053\,
            I => \b2v_inst36.countZ0Z_15\
        );

    \I__5688\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28045\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__28045\,
            I => \N__28042\
        );

    \I__5686\ : Span4Mux_v
    port map (
            O => \N__28042\,
            I => \N__28039\
        );

    \I__5685\ : Odrv4
    port map (
            O => \N__28039\,
            I => \b2v_inst5.un12_clk_100khz_4\
        );

    \I__5684\ : InMux
    port map (
            O => \N__28036\,
            I => \N__28030\
        );

    \I__5683\ : InMux
    port map (
            O => \N__28035\,
            I => \N__28030\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__28030\,
            I => \b2v_inst5.count_1_2\
        );

    \I__5681\ : InMux
    port map (
            O => \N__28027\,
            I => \N__28022\
        );

    \I__5680\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28019\
        );

    \I__5679\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28016\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__28022\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__28019\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__28016\,
            I => \b2v_inst36.countZ0Z_11\
        );

    \I__5675\ : InMux
    port map (
            O => \N__28009\,
            I => \N__28003\
        );

    \I__5674\ : InMux
    port map (
            O => \N__28008\,
            I => \N__28003\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__28003\,
            I => \b2v_inst36.un2_count_1_cry_10_THRU_CO\
        );

    \I__5672\ : InMux
    port map (
            O => \N__28000\,
            I => \b2v_inst36.un2_count_1_cry_10\
        );

    \I__5671\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27993\
        );

    \I__5670\ : CascadeMux
    port map (
            O => \N__27996\,
            I => \N__27990\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27987\
        );

    \I__5668\ : InMux
    port map (
            O => \N__27990\,
            I => \N__27984\
        );

    \I__5667\ : Span4Mux_h
    port map (
            O => \N__27987\,
            I => \N__27981\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__27984\,
            I => \b2v_inst36.countZ0Z_12\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__27981\,
            I => \b2v_inst36.countZ0Z_12\
        );

    \I__5664\ : InMux
    port map (
            O => \N__27976\,
            I => \N__27972\
        );

    \I__5663\ : InMux
    port map (
            O => \N__27975\,
            I => \N__27969\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27972\,
            I => \N__27964\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__27969\,
            I => \N__27964\
        );

    \I__5660\ : Span4Mux_s1_v
    port map (
            O => \N__27964\,
            I => \N__27961\
        );

    \I__5659\ : Odrv4
    port map (
            O => \N__27961\,
            I => \b2v_inst36.count_rst_2\
        );

    \I__5658\ : InMux
    port map (
            O => \N__27958\,
            I => \b2v_inst36.un2_count_1_cry_11\
        );

    \I__5657\ : InMux
    port map (
            O => \N__27955\,
            I => \b2v_inst36.un2_count_1_cry_12\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__27952\,
            I => \N__27949\
        );

    \I__5655\ : InMux
    port map (
            O => \N__27949\,
            I => \N__27945\
        );

    \I__5654\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27942\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__27945\,
            I => \N__27937\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27937\
        );

    \I__5651\ : Odrv4
    port map (
            O => \N__27937\,
            I => \b2v_inst36.countZ0Z_14\
        );

    \I__5650\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27930\
        );

    \I__5649\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27927\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__27930\,
            I => \N__27924\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27927\,
            I => \N__27921\
        );

    \I__5646\ : Odrv4
    port map (
            O => \N__27924\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__5645\ : Odrv4
    port map (
            O => \N__27921\,
            I => \b2v_inst36.count_rst_0\
        );

    \I__5644\ : InMux
    port map (
            O => \N__27916\,
            I => \b2v_inst36.un2_count_1_cry_13\
        );

    \I__5643\ : InMux
    port map (
            O => \N__27913\,
            I => \b2v_inst36.un2_count_1_cry_14\
        );

    \I__5642\ : InMux
    port map (
            O => \N__27910\,
            I => \N__27907\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__27907\,
            I => \b2v_inst36.count_rst_6\
        );

    \I__5640\ : InMux
    port map (
            O => \N__27904\,
            I => \N__27899\
        );

    \I__5639\ : InMux
    port map (
            O => \N__27903\,
            I => \N__27896\
        );

    \I__5638\ : InMux
    port map (
            O => \N__27902\,
            I => \N__27893\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__27899\,
            I => \N__27890\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27887\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__27893\,
            I => \N__27884\
        );

    \I__5634\ : Odrv4
    port map (
            O => \N__27890\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__5633\ : Odrv12
    port map (
            O => \N__27887\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__5632\ : Odrv4
    port map (
            O => \N__27884\,
            I => \b2v_inst36.countZ0Z_8\
        );

    \I__5631\ : InMux
    port map (
            O => \N__27877\,
            I => \N__27873\
        );

    \I__5630\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27870\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__27873\,
            I => \N__27865\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__27870\,
            I => \N__27865\
        );

    \I__5627\ : Span4Mux_h
    port map (
            O => \N__27865\,
            I => \N__27862\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__27862\,
            I => \b2v_inst36.un2_count_1_cry_7_THRU_CO\
        );

    \I__5625\ : CascadeMux
    port map (
            O => \N__27859\,
            I => \b2v_inst36.countZ0Z_8_cascade_\
        );

    \I__5624\ : InMux
    port map (
            O => \N__27856\,
            I => \N__27853\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__27853\,
            I => \b2v_inst36.count_2_8\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27850\,
            I => \N__27844\
        );

    \I__5621\ : InMux
    port map (
            O => \N__27849\,
            I => \N__27844\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__27844\,
            I => \b2v_inst36.un2_count_1_cry_1_THRU_CO\
        );

    \I__5619\ : InMux
    port map (
            O => \N__27841\,
            I => \b2v_inst36.un2_count_1_cry_1\
        );

    \I__5618\ : InMux
    port map (
            O => \N__27838\,
            I => \b2v_inst36.un2_count_1_cry_2\
        );

    \I__5617\ : InMux
    port map (
            O => \N__27835\,
            I => \N__27831\
        );

    \I__5616\ : InMux
    port map (
            O => \N__27834\,
            I => \N__27828\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27825\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__27828\,
            I => \b2v_inst36.countZ0Z_4\
        );

    \I__5613\ : Odrv12
    port map (
            O => \N__27825\,
            I => \b2v_inst36.countZ0Z_4\
        );

    \I__5612\ : InMux
    port map (
            O => \N__27820\,
            I => \N__27814\
        );

    \I__5611\ : InMux
    port map (
            O => \N__27819\,
            I => \N__27814\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__27814\,
            I => \N__27811\
        );

    \I__5609\ : Odrv4
    port map (
            O => \N__27811\,
            I => \b2v_inst36.count_rst_10\
        );

    \I__5608\ : InMux
    port map (
            O => \N__27808\,
            I => \b2v_inst36.un2_count_1_cry_3\
        );

    \I__5607\ : InMux
    port map (
            O => \N__27805\,
            I => \b2v_inst36.un2_count_1_cry_4\
        );

    \I__5606\ : InMux
    port map (
            O => \N__27802\,
            I => \N__27798\
        );

    \I__5605\ : InMux
    port map (
            O => \N__27801\,
            I => \N__27795\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__27798\,
            I => \N__27790\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__27795\,
            I => \N__27790\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__27790\,
            I => \b2v_inst36.countZ0Z_6\
        );

    \I__5601\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27781\
        );

    \I__5600\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27781\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__27781\,
            I => \N__27778\
        );

    \I__5598\ : Odrv12
    port map (
            O => \N__27778\,
            I => \b2v_inst36.count_rst_8\
        );

    \I__5597\ : InMux
    port map (
            O => \N__27775\,
            I => \b2v_inst36.un2_count_1_cry_5\
        );

    \I__5596\ : InMux
    port map (
            O => \N__27772\,
            I => \b2v_inst36.un2_count_1_cry_6\
        );

    \I__5595\ : InMux
    port map (
            O => \N__27769\,
            I => \b2v_inst36.un2_count_1_cry_7\
        );

    \I__5594\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27763\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__27763\,
            I => \N__27759\
        );

    \I__5592\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27756\
        );

    \I__5591\ : Span4Mux_h
    port map (
            O => \N__27759\,
            I => \N__27753\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__27756\,
            I => \b2v_inst36.countZ0Z_9\
        );

    \I__5589\ : Odrv4
    port map (
            O => \N__27753\,
            I => \b2v_inst36.countZ0Z_9\
        );

    \I__5588\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27744\
        );

    \I__5587\ : InMux
    port map (
            O => \N__27747\,
            I => \N__27741\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__27744\,
            I => \N__27736\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__27741\,
            I => \N__27736\
        );

    \I__5584\ : Span4Mux_s1_v
    port map (
            O => \N__27736\,
            I => \N__27733\
        );

    \I__5583\ : Odrv4
    port map (
            O => \N__27733\,
            I => \b2v_inst36.count_rst_5\
        );

    \I__5582\ : InMux
    port map (
            O => \N__27730\,
            I => \bfn_9_2_0_\
        );

    \I__5581\ : InMux
    port map (
            O => \N__27727\,
            I => \b2v_inst36.un2_count_1_cry_9\
        );

    \I__5580\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27715\
        );

    \I__5579\ : InMux
    port map (
            O => \N__27723\,
            I => \N__27711\
        );

    \I__5578\ : InMux
    port map (
            O => \N__27722\,
            I => \N__27707\
        );

    \I__5577\ : InMux
    port map (
            O => \N__27721\,
            I => \N__27702\
        );

    \I__5576\ : InMux
    port map (
            O => \N__27720\,
            I => \N__27702\
        );

    \I__5575\ : InMux
    port map (
            O => \N__27719\,
            I => \N__27695\
        );

    \I__5574\ : InMux
    port map (
            O => \N__27718\,
            I => \N__27695\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__27715\,
            I => \N__27692\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__27714\,
            I => \N__27689\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__27711\,
            I => \N__27684\
        );

    \I__5570\ : InMux
    port map (
            O => \N__27710\,
            I => \N__27681\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__27707\,
            I => \N__27676\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__27702\,
            I => \N__27676\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__27701\,
            I => \N__27673\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__27700\,
            I => \N__27665\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__27695\,
            I => \N__27660\
        );

    \I__5564\ : Span4Mux_h
    port map (
            O => \N__27692\,
            I => \N__27654\
        );

    \I__5563\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27651\
        );

    \I__5562\ : InMux
    port map (
            O => \N__27688\,
            I => \N__27646\
        );

    \I__5561\ : InMux
    port map (
            O => \N__27687\,
            I => \N__27646\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__27684\,
            I => \N__27639\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__27681\,
            I => \N__27639\
        );

    \I__5558\ : Span4Mux_h
    port map (
            O => \N__27676\,
            I => \N__27639\
        );

    \I__5557\ : InMux
    port map (
            O => \N__27673\,
            I => \N__27634\
        );

    \I__5556\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27634\
        );

    \I__5555\ : InMux
    port map (
            O => \N__27671\,
            I => \N__27629\
        );

    \I__5554\ : InMux
    port map (
            O => \N__27670\,
            I => \N__27629\
        );

    \I__5553\ : InMux
    port map (
            O => \N__27669\,
            I => \N__27624\
        );

    \I__5552\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27624\
        );

    \I__5551\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27617\
        );

    \I__5550\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27617\
        );

    \I__5549\ : InMux
    port map (
            O => \N__27663\,
            I => \N__27617\
        );

    \I__5548\ : Span4Mux_h
    port map (
            O => \N__27660\,
            I => \N__27614\
        );

    \I__5547\ : InMux
    port map (
            O => \N__27659\,
            I => \N__27607\
        );

    \I__5546\ : InMux
    port map (
            O => \N__27658\,
            I => \N__27607\
        );

    \I__5545\ : InMux
    port map (
            O => \N__27657\,
            I => \N__27607\
        );

    \I__5544\ : Span4Mux_v
    port map (
            O => \N__27654\,
            I => \N__27604\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__27651\,
            I => \N__27596\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__27646\,
            I => \N__27596\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__27639\,
            I => \N__27596\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__27634\,
            I => \N__27586\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__27629\,
            I => \N__27586\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27586\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__27617\,
            I => \N__27586\
        );

    \I__5536\ : Span4Mux_v
    port map (
            O => \N__27614\,
            I => \N__27581\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__27607\,
            I => \N__27581\
        );

    \I__5534\ : Span4Mux_v
    port map (
            O => \N__27604\,
            I => \N__27578\
        );

    \I__5533\ : IoInMux
    port map (
            O => \N__27603\,
            I => \N__27575\
        );

    \I__5532\ : Span4Mux_v
    port map (
            O => \N__27596\,
            I => \N__27572\
        );

    \I__5531\ : InMux
    port map (
            O => \N__27595\,
            I => \N__27569\
        );

    \I__5530\ : Span4Mux_v
    port map (
            O => \N__27586\,
            I => \N__27564\
        );

    \I__5529\ : Span4Mux_h
    port map (
            O => \N__27581\,
            I => \N__27564\
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__27578\,
            I => \G_146\
        );

    \I__5527\ : LocalMux
    port map (
            O => \N__27575\,
            I => \G_146\
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__27572\,
            I => \G_146\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__27569\,
            I => \G_146\
        );

    \I__5524\ : Odrv4
    port map (
            O => \N__27564\,
            I => \G_146\
        );

    \I__5523\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27549\
        );

    \I__5522\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27546\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__27549\,
            I => \N__27543\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__27546\,
            I => \N__27538\
        );

    \I__5519\ : Span4Mux_h
    port map (
            O => \N__27543\,
            I => \N__27538\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__27538\,
            I => \N_15_i_0_a4_1\
        );

    \I__5517\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27531\
        );

    \I__5516\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27528\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__27531\,
            I => \N__27525\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27522\
        );

    \I__5513\ : Span4Mux_h
    port map (
            O => \N__27525\,
            I => \N__27519\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__27522\,
            I => \N__27516\
        );

    \I__5511\ : Odrv4
    port map (
            O => \N__27519\,
            I => \N_73_mux_i_i_a7_0_0\
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__27516\,
            I => \N_73_mux_i_i_a7_0_0\
        );

    \I__5509\ : InMux
    port map (
            O => \N__27511\,
            I => \N__27505\
        );

    \I__5508\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27505\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__27505\,
            I => \N__27502\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__27502\,
            I => \b2v_inst11.count_1_8\
        );

    \I__5505\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27496\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__27496\,
            I => \b2v_inst11.count_0_8\
        );

    \I__5503\ : InMux
    port map (
            O => \N__27493\,
            I => \N__27490\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27487\
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__27487\,
            I => \b2v_inst11.g0_2_1\
        );

    \I__5500\ : InMux
    port map (
            O => \N__27484\,
            I => \N__27480\
        );

    \I__5499\ : InMux
    port map (
            O => \N__27483\,
            I => \N__27477\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__27480\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__27477\,
            I => \b2v_inst11.pwm_outZ0\
        );

    \I__5496\ : SRMux
    port map (
            O => \N__27472\,
            I => \N__27469\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__27469\,
            I => \N__27466\
        );

    \I__5494\ : Odrv12
    port map (
            O => \N__27466\,
            I => \b2v_inst11.pwm_out_1_sqmuxa\
        );

    \I__5493\ : CascadeMux
    port map (
            O => \N__27463\,
            I => \b2v_inst11.curr_state_3_0_cascade_\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__27460\,
            I => \b2v_inst11.curr_stateZ0Z_0_cascade_\
        );

    \I__5491\ : InMux
    port map (
            O => \N__27457\,
            I => \N__27441\
        );

    \I__5490\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27441\
        );

    \I__5489\ : InMux
    port map (
            O => \N__27455\,
            I => \N__27441\
        );

    \I__5488\ : InMux
    port map (
            O => \N__27454\,
            I => \N__27430\
        );

    \I__5487\ : InMux
    port map (
            O => \N__27453\,
            I => \N__27430\
        );

    \I__5486\ : InMux
    port map (
            O => \N__27452\,
            I => \N__27430\
        );

    \I__5485\ : InMux
    port map (
            O => \N__27451\,
            I => \N__27421\
        );

    \I__5484\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27421\
        );

    \I__5483\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27421\
        );

    \I__5482\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27421\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__27441\,
            I => \N__27415\
        );

    \I__5480\ : InMux
    port map (
            O => \N__27440\,
            I => \N__27406\
        );

    \I__5479\ : InMux
    port map (
            O => \N__27439\,
            I => \N__27406\
        );

    \I__5478\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27406\
        );

    \I__5477\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27406\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__27430\,
            I => \N__27403\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__27421\,
            I => \N__27400\
        );

    \I__5474\ : InMux
    port map (
            O => \N__27420\,
            I => \N__27395\
        );

    \I__5473\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27395\
        );

    \I__5472\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27392\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__27415\,
            I => \N__27389\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__27406\,
            I => \N__27382\
        );

    \I__5469\ : Span4Mux_h
    port map (
            O => \N__27403\,
            I => \N__27382\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__27400\,
            I => \N__27382\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__27395\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__27392\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5465\ : Odrv4
    port map (
            O => \N__27389\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__27382\,
            I => \b2v_inst11.count_0_sqmuxa_i\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__27373\,
            I => \b2v_inst11.count_0_sqmuxa_i_cascade_\
        );

    \I__5462\ : InMux
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__27367\,
            I => \b2v_inst11.count_1_0\
        );

    \I__5460\ : InMux
    port map (
            O => \N__27364\,
            I => \N__27360\
        );

    \I__5459\ : InMux
    port map (
            O => \N__27363\,
            I => \N__27357\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__27360\,
            I => \b2v_inst36.un2_count_1_axb_1\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__27357\,
            I => \b2v_inst36.un2_count_1_axb_1\
        );

    \I__5456\ : CascadeMux
    port map (
            O => \N__27352\,
            I => \N__27345\
        );

    \I__5455\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27340\
        );

    \I__5454\ : InMux
    port map (
            O => \N__27350\,
            I => \N__27340\
        );

    \I__5453\ : InMux
    port map (
            O => \N__27349\,
            I => \N__27335\
        );

    \I__5452\ : InMux
    port map (
            O => \N__27348\,
            I => \N__27335\
        );

    \I__5451\ : InMux
    port map (
            O => \N__27345\,
            I => \N__27332\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__27340\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__27335\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__27332\,
            I => \b2v_inst36.countZ0Z_0\
        );

    \I__5447\ : InMux
    port map (
            O => \N__27325\,
            I => \N__27322\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__27322\,
            I => \b2v_inst11.un79_clk_100khzlt6\
        );

    \I__5445\ : CascadeMux
    port map (
            O => \N__27319\,
            I => \b2v_inst11.un79_clk_100khzlto15_4_cascade_\
        );

    \I__5444\ : InMux
    port map (
            O => \N__27316\,
            I => \N__27313\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__27313\,
            I => \b2v_inst11.un79_clk_100khzlto15_7\
        );

    \I__5442\ : CascadeMux
    port map (
            O => \N__27310\,
            I => \b2v_inst11.count_RNIZ0Z_13_cascade_\
        );

    \I__5441\ : CascadeMux
    port map (
            O => \N__27307\,
            I => \b2v_inst11.countZ0Z_0_cascade_\
        );

    \I__5440\ : CascadeMux
    port map (
            O => \N__27304\,
            I => \b2v_inst11.count_1_1_cascade_\
        );

    \I__5439\ : CascadeMux
    port map (
            O => \N__27301\,
            I => \b2v_inst11.countZ0Z_1_cascade_\
        );

    \I__5438\ : InMux
    port map (
            O => \N__27298\,
            I => \N__27295\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__27295\,
            I => \b2v_inst11.count_0_1\
        );

    \I__5436\ : InMux
    port map (
            O => \N__27292\,
            I => \N__27289\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__27289\,
            I => \b2v_inst11.count_0_0\
        );

    \I__5434\ : InMux
    port map (
            O => \N__27286\,
            I => \N__27282\
        );

    \I__5433\ : CascadeMux
    port map (
            O => \N__27285\,
            I => \N__27279\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__27282\,
            I => \N__27276\
        );

    \I__5431\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27273\
        );

    \I__5430\ : Span4Mux_h
    port map (
            O => \N__27276\,
            I => \N__27268\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__27273\,
            I => \N__27268\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__27268\,
            I => \N__27265\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__27265\,
            I => \N__27262\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__27262\,
            I => \N__27259\
        );

    \I__5425\ : Odrv4
    port map (
            O => \N__27259\,
            I => b2v_inst11_dutycycle_set_1
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__27256\,
            I => \N__27253\
        );

    \I__5423\ : InMux
    port map (
            O => \N__27253\,
            I => \N__27247\
        );

    \I__5422\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27247\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__27247\,
            I => \b2v_inst11.count_1_3\
        );

    \I__5420\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27241\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__27241\,
            I => \b2v_inst11.count_0_3\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__27238\,
            I => \N__27235\
        );

    \I__5417\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27229\
        );

    \I__5416\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27229\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__27229\,
            I => \b2v_inst11.count_1_13\
        );

    \I__5414\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27223\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__27223\,
            I => \b2v_inst11.count_0_13\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__27220\,
            I => \N__27217\
        );

    \I__5411\ : InMux
    port map (
            O => \N__27217\,
            I => \N__27211\
        );

    \I__5410\ : InMux
    port map (
            O => \N__27216\,
            I => \N__27211\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__27211\,
            I => \b2v_inst11.count_1_4\
        );

    \I__5408\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27205\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__27205\,
            I => \b2v_inst11.count_0_4\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__27202\,
            I => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\
        );

    \I__5405\ : InMux
    port map (
            O => \N__27199\,
            I => \N__27196\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__27193\,
            I => \N__27190\
        );

    \I__5402\ : Odrv4
    port map (
            O => \N__27190\,
            I => \b2v_inst11.g2_0_0\
        );

    \I__5401\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__27184\,
            I => b2v_inst11_un1_dutycycle_164_0
        );

    \I__5399\ : CascadeMux
    port map (
            O => \N__27181\,
            I => \N__27178\
        );

    \I__5398\ : InMux
    port map (
            O => \N__27178\,
            I => \N__27172\
        );

    \I__5397\ : InMux
    port map (
            O => \N__27177\,
            I => \N__27172\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__5395\ : Odrv12
    port map (
            O => \N__27169\,
            I => \b2v_inst5.N_6\
        );

    \I__5394\ : CascadeMux
    port map (
            O => \N__27166\,
            I => \b2v_inst11_un1_dutycycle_164_0_cascade_\
        );

    \I__5393\ : InMux
    port map (
            O => \N__27163\,
            I => \N__27160\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__27160\,
            I => \N__27157\
        );

    \I__5391\ : Span4Mux_h
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__27154\,
            I => \b2v_inst5.N_13\
        );

    \I__5389\ : CascadeMux
    port map (
            O => \N__27151\,
            I => \N__27143\
        );

    \I__5388\ : CascadeMux
    port map (
            O => \N__27150\,
            I => \N__27139\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__27149\,
            I => \N__27136\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__27148\,
            I => \N__27133\
        );

    \I__5385\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27126\
        );

    \I__5384\ : CascadeMux
    port map (
            O => \N__27146\,
            I => \N__27123\
        );

    \I__5383\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27120\
        );

    \I__5382\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27117\
        );

    \I__5381\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27114\
        );

    \I__5380\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27109\
        );

    \I__5379\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27109\
        );

    \I__5378\ : CascadeMux
    port map (
            O => \N__27132\,
            I => \N__27105\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__27131\,
            I => \N__27097\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__27130\,
            I => \N__27093\
        );

    \I__5375\ : CascadeMux
    port map (
            O => \N__27129\,
            I => \N__27089\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__27126\,
            I => \N__27085\
        );

    \I__5373\ : InMux
    port map (
            O => \N__27123\,
            I => \N__27082\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__27120\,
            I => \N__27079\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__27117\,
            I => \N__27075\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__27114\,
            I => \N__27070\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__27109\,
            I => \N__27070\
        );

    \I__5368\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27065\
        );

    \I__5367\ : InMux
    port map (
            O => \N__27105\,
            I => \N__27065\
        );

    \I__5366\ : CascadeMux
    port map (
            O => \N__27104\,
            I => \N__27060\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__27103\,
            I => \N__27055\
        );

    \I__5364\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27051\
        );

    \I__5363\ : InMux
    port map (
            O => \N__27101\,
            I => \N__27034\
        );

    \I__5362\ : InMux
    port map (
            O => \N__27100\,
            I => \N__27034\
        );

    \I__5361\ : InMux
    port map (
            O => \N__27097\,
            I => \N__27034\
        );

    \I__5360\ : InMux
    port map (
            O => \N__27096\,
            I => \N__27034\
        );

    \I__5359\ : InMux
    port map (
            O => \N__27093\,
            I => \N__27034\
        );

    \I__5358\ : InMux
    port map (
            O => \N__27092\,
            I => \N__27034\
        );

    \I__5357\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27034\
        );

    \I__5356\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27034\
        );

    \I__5355\ : Span4Mux_v
    port map (
            O => \N__27085\,
            I => \N__27029\
        );

    \I__5354\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27029\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__27079\,
            I => \N__27026\
        );

    \I__5352\ : InMux
    port map (
            O => \N__27078\,
            I => \N__27023\
        );

    \I__5351\ : Span4Mux_v
    port map (
            O => \N__27075\,
            I => \N__27018\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__27070\,
            I => \N__27018\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__27065\,
            I => \N__27015\
        );

    \I__5348\ : InMux
    port map (
            O => \N__27064\,
            I => \N__27010\
        );

    \I__5347\ : InMux
    port map (
            O => \N__27063\,
            I => \N__27010\
        );

    \I__5346\ : InMux
    port map (
            O => \N__27060\,
            I => \N__26999\
        );

    \I__5345\ : InMux
    port map (
            O => \N__27059\,
            I => \N__26999\
        );

    \I__5344\ : InMux
    port map (
            O => \N__27058\,
            I => \N__26999\
        );

    \I__5343\ : InMux
    port map (
            O => \N__27055\,
            I => \N__26999\
        );

    \I__5342\ : InMux
    port map (
            O => \N__27054\,
            I => \N__26999\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__27051\,
            I => \N__26992\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__27034\,
            I => \N__26992\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__27029\,
            I => \N__26992\
        );

    \I__5338\ : Odrv4
    port map (
            O => \N__27026\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__27023\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5336\ : Odrv4
    port map (
            O => \N__27018\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__27015\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__27010\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__26999\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__26992\,
            I => \b2v_inst11.N_3060_i\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26977\,
            I => \N__26971\
        );

    \I__5330\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26971\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__26971\,
            I => \N__26968\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__26968\,
            I => \N__26965\
        );

    \I__5327\ : Odrv4
    port map (
            O => \N__26965\,
            I => \b2v_inst11.un1_dutycycle_96_0_a3_1\
        );

    \I__5326\ : InMux
    port map (
            O => \N__26962\,
            I => \N__26959\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__26959\,
            I => \N__26956\
        );

    \I__5324\ : Span4Mux_h
    port map (
            O => \N__26956\,
            I => \N__26953\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__5322\ : Odrv4
    port map (
            O => \N__26950\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_7\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__5320\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26938\
        );

    \I__5319\ : InMux
    port map (
            O => \N__26943\,
            I => \N__26935\
        );

    \I__5318\ : InMux
    port map (
            O => \N__26942\,
            I => \N__26932\
        );

    \I__5317\ : InMux
    port map (
            O => \N__26941\,
            I => \N__26928\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__26938\,
            I => \N__26925\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__26935\,
            I => \N__26922\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__26932\,
            I => \N__26919\
        );

    \I__5313\ : CascadeMux
    port map (
            O => \N__26931\,
            I => \N__26916\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__26928\,
            I => \N__26912\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__26925\,
            I => \N__26909\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__26922\,
            I => \N__26904\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__26919\,
            I => \N__26904\
        );

    \I__5308\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26899\
        );

    \I__5307\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26899\
        );

    \I__5306\ : Span4Mux_h
    port map (
            O => \N__26912\,
            I => \N__26896\
        );

    \I__5305\ : Odrv4
    port map (
            O => \N__26909\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__26904\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__26899\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__26896\,
            I => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\
        );

    \I__5301\ : CascadeMux
    port map (
            O => \N__26887\,
            I => \N__26883\
        );

    \I__5300\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26880\
        );

    \I__5299\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26877\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__26880\,
            I => \N__26873\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__26877\,
            I => \N__26870\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26876\,
            I => \N__26867\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__26873\,
            I => \N__26864\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__26870\,
            I => \N__26861\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__26867\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5\
        );

    \I__5292\ : Odrv4
    port map (
            O => \N__26864\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__26861\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5\
        );

    \I__5290\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26848\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26848\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__26848\,
            I => \N_73_mux_i_i_o3_1_1\
        );

    \I__5287\ : CascadeMux
    port map (
            O => \N__26845\,
            I => \N__26839\
        );

    \I__5286\ : CascadeMux
    port map (
            O => \N__26844\,
            I => \N__26827\
        );

    \I__5285\ : CascadeMux
    port map (
            O => \N__26843\,
            I => \N__26824\
        );

    \I__5284\ : CascadeMux
    port map (
            O => \N__26842\,
            I => \N__26820\
        );

    \I__5283\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26817\
        );

    \I__5282\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26812\
        );

    \I__5281\ : InMux
    port map (
            O => \N__26837\,
            I => \N__26812\
        );

    \I__5280\ : CascadeMux
    port map (
            O => \N__26836\,
            I => \N__26809\
        );

    \I__5279\ : InMux
    port map (
            O => \N__26835\,
            I => \N__26801\
        );

    \I__5278\ : InMux
    port map (
            O => \N__26834\,
            I => \N__26801\
        );

    \I__5277\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26801\
        );

    \I__5276\ : CascadeMux
    port map (
            O => \N__26832\,
            I => \N__26795\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__26831\,
            I => \N__26792\
        );

    \I__5274\ : InMux
    port map (
            O => \N__26830\,
            I => \N__26784\
        );

    \I__5273\ : InMux
    port map (
            O => \N__26827\,
            I => \N__26784\
        );

    \I__5272\ : InMux
    port map (
            O => \N__26824\,
            I => \N__26781\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__26823\,
            I => \N__26778\
        );

    \I__5270\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26773\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__26817\,
            I => \N__26768\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__26812\,
            I => \N__26768\
        );

    \I__5267\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26763\
        );

    \I__5266\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26763\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__26801\,
            I => \N__26760\
        );

    \I__5264\ : InMux
    port map (
            O => \N__26800\,
            I => \N__26751\
        );

    \I__5263\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26751\
        );

    \I__5262\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26751\
        );

    \I__5261\ : InMux
    port map (
            O => \N__26795\,
            I => \N__26751\
        );

    \I__5260\ : InMux
    port map (
            O => \N__26792\,
            I => \N__26745\
        );

    \I__5259\ : InMux
    port map (
            O => \N__26791\,
            I => \N__26745\
        );

    \I__5258\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26740\
        );

    \I__5257\ : InMux
    port map (
            O => \N__26789\,
            I => \N__26740\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__26784\,
            I => \N__26737\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__26781\,
            I => \N__26734\
        );

    \I__5254\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26731\
        );

    \I__5253\ : InMux
    port map (
            O => \N__26777\,
            I => \N__26726\
        );

    \I__5252\ : InMux
    port map (
            O => \N__26776\,
            I => \N__26726\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__26773\,
            I => \N__26723\
        );

    \I__5250\ : Span4Mux_v
    port map (
            O => \N__26768\,
            I => \N__26718\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__26763\,
            I => \N__26718\
        );

    \I__5248\ : Span4Mux_h
    port map (
            O => \N__26760\,
            I => \N__26713\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26713\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__26750\,
            I => \N__26709\
        );

    \I__5245\ : LocalMux
    port map (
            O => \N__26745\,
            I => \N__26706\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__26740\,
            I => \N__26703\
        );

    \I__5243\ : Span4Mux_h
    port map (
            O => \N__26737\,
            I => \N__26700\
        );

    \I__5242\ : Span4Mux_v
    port map (
            O => \N__26734\,
            I => \N__26693\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26693\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__26726\,
            I => \N__26693\
        );

    \I__5239\ : Span4Mux_h
    port map (
            O => \N__26723\,
            I => \N__26688\
        );

    \I__5238\ : Span4Mux_h
    port map (
            O => \N__26718\,
            I => \N__26688\
        );

    \I__5237\ : Span4Mux_v
    port map (
            O => \N__26713\,
            I => \N__26685\
        );

    \I__5236\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26680\
        );

    \I__5235\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26680\
        );

    \I__5234\ : Odrv12
    port map (
            O => \N__26706\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5233\ : Odrv4
    port map (
            O => \N__26703\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__26700\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__26693\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5230\ : Odrv4
    port map (
            O => \N__26688\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5229\ : Odrv4
    port map (
            O => \N__26685\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__26680\,
            I => \b2v_inst11.dutycycleZ1Z_3\
        );

    \I__5227\ : CascadeMux
    port map (
            O => \N__26665\,
            I => \N__26662\
        );

    \I__5226\ : InMux
    port map (
            O => \N__26662\,
            I => \N__26659\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__26659\,
            I => \N__26656\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__26656\,
            I => \N__26653\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__26653\,
            I => \b2v_inst11.g3_0_1\
        );

    \I__5222\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26638\
        );

    \I__5221\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26629\
        );

    \I__5220\ : InMux
    port map (
            O => \N__26648\,
            I => \N__26626\
        );

    \I__5219\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26623\
        );

    \I__5218\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26616\
        );

    \I__5217\ : InMux
    port map (
            O => \N__26645\,
            I => \N__26616\
        );

    \I__5216\ : InMux
    port map (
            O => \N__26644\,
            I => \N__26616\
        );

    \I__5215\ : InMux
    port map (
            O => \N__26643\,
            I => \N__26613\
        );

    \I__5214\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26608\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__26641\,
            I => \N__26605\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__26638\,
            I => \N__26602\
        );

    \I__5211\ : InMux
    port map (
            O => \N__26637\,
            I => \N__26597\
        );

    \I__5210\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26597\
        );

    \I__5209\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26594\
        );

    \I__5208\ : InMux
    port map (
            O => \N__26634\,
            I => \N__26591\
        );

    \I__5207\ : CascadeMux
    port map (
            O => \N__26633\,
            I => \N__26588\
        );

    \I__5206\ : InMux
    port map (
            O => \N__26632\,
            I => \N__26584\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__26629\,
            I => \N__26579\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__26626\,
            I => \N__26579\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26576\
        );

    \I__5202\ : LocalMux
    port map (
            O => \N__26616\,
            I => \N__26571\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__26613\,
            I => \N__26571\
        );

    \I__5200\ : InMux
    port map (
            O => \N__26612\,
            I => \N__26563\
        );

    \I__5199\ : InMux
    port map (
            O => \N__26611\,
            I => \N__26563\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__26608\,
            I => \N__26560\
        );

    \I__5197\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26557\
        );

    \I__5196\ : Span4Mux_v
    port map (
            O => \N__26602\,
            I => \N__26552\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__26597\,
            I => \N__26552\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__26594\,
            I => \N__26547\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__26591\,
            I => \N__26547\
        );

    \I__5192\ : InMux
    port map (
            O => \N__26588\,
            I => \N__26542\
        );

    \I__5191\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26542\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26539\
        );

    \I__5189\ : Span4Mux_v
    port map (
            O => \N__26579\,
            I => \N__26534\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__26576\,
            I => \N__26534\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__26571\,
            I => \N__26531\
        );

    \I__5186\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26526\
        );

    \I__5185\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26526\
        );

    \I__5184\ : InMux
    port map (
            O => \N__26568\,
            I => \N__26523\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__26563\,
            I => \N__26520\
        );

    \I__5182\ : Span4Mux_s3_v
    port map (
            O => \N__26560\,
            I => \N__26517\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__26557\,
            I => \N__26508\
        );

    \I__5180\ : Span4Mux_h
    port map (
            O => \N__26552\,
            I => \N__26508\
        );

    \I__5179\ : Span4Mux_v
    port map (
            O => \N__26547\,
            I => \N__26508\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__26542\,
            I => \N__26508\
        );

    \I__5177\ : Span4Mux_v
    port map (
            O => \N__26539\,
            I => \N__26505\
        );

    \I__5176\ : Sp12to4
    port map (
            O => \N__26534\,
            I => \N__26496\
        );

    \I__5175\ : Sp12to4
    port map (
            O => \N__26531\,
            I => \N__26496\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__26526\,
            I => \N__26496\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__26523\,
            I => \N__26496\
        );

    \I__5172\ : Span4Mux_v
    port map (
            O => \N__26520\,
            I => \N__26489\
        );

    \I__5171\ : Span4Mux_h
    port map (
            O => \N__26517\,
            I => \N__26489\
        );

    \I__5170\ : Span4Mux_h
    port map (
            O => \N__26508\,
            I => \N__26489\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__26505\,
            I => \b2v_inst11.N_3038_i\
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__26496\,
            I => \b2v_inst11.N_3038_i\
        );

    \I__5167\ : Odrv4
    port map (
            O => \N__26489\,
            I => \b2v_inst11.N_3038_i\
        );

    \I__5166\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26478\
        );

    \I__5165\ : InMux
    port map (
            O => \N__26481\,
            I => \N__26475\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__26478\,
            I => g3_0_4
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__26475\,
            I => g3_0_4
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__26470\,
            I => \N__26467\
        );

    \I__5161\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26461\
        );

    \I__5160\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26461\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__26461\,
            I => \b2v_inst11.count_1_12\
        );

    \I__5158\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26455\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__26455\,
            I => \b2v_inst11.count_0_12\
        );

    \I__5156\ : InMux
    port map (
            O => \N__26452\,
            I => \N__26442\
        );

    \I__5155\ : CascadeMux
    port map (
            O => \N__26451\,
            I => \N__26439\
        );

    \I__5154\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26427\
        );

    \I__5153\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26427\
        );

    \I__5152\ : InMux
    port map (
            O => \N__26448\,
            I => \N__26422\
        );

    \I__5151\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26415\
        );

    \I__5150\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26415\
        );

    \I__5149\ : InMux
    port map (
            O => \N__26445\,
            I => \N__26415\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__26442\,
            I => \N__26412\
        );

    \I__5147\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26409\
        );

    \I__5146\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26406\
        );

    \I__5145\ : InMux
    port map (
            O => \N__26437\,
            I => \N__26403\
        );

    \I__5144\ : InMux
    port map (
            O => \N__26436\,
            I => \N__26398\
        );

    \I__5143\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26398\
        );

    \I__5142\ : InMux
    port map (
            O => \N__26434\,
            I => \N__26391\
        );

    \I__5141\ : InMux
    port map (
            O => \N__26433\,
            I => \N__26391\
        );

    \I__5140\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26391\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__26427\,
            I => \N__26388\
        );

    \I__5138\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26383\
        );

    \I__5137\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26383\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__26422\,
            I => \N__26380\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__26415\,
            I => \N__26375\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__26412\,
            I => \N__26375\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__26409\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__26406\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__26403\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__26398\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__26391\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__26388\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__26383\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5126\ : Odrv4
    port map (
            O => \N__26380\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5125\ : Odrv4
    port map (
            O => \N__26375\,
            I => \b2v_inst11.dutycycleZ0Z_1\
        );

    \I__5124\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26353\
        );

    \I__5123\ : LocalMux
    port map (
            O => \N__26353\,
            I => \b2v_inst11.un1_dutycycle_53_50_1_i_0_1\
        );

    \I__5122\ : InMux
    port map (
            O => \N__26350\,
            I => \N__26347\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__26347\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_1\
        );

    \I__5120\ : CascadeMux
    port map (
            O => \N__26344\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_1_cascade_\
        );

    \I__5119\ : CascadeMux
    port map (
            O => \N__26341\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_3_cascade_\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__26338\,
            I => \N__26330\
        );

    \I__5117\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26323\
        );

    \I__5116\ : CascadeMux
    port map (
            O => \N__26336\,
            I => \N__26320\
        );

    \I__5115\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26317\
        );

    \I__5114\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26310\
        );

    \I__5113\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26310\
        );

    \I__5112\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26310\
        );

    \I__5111\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26305\
        );

    \I__5110\ : InMux
    port map (
            O => \N__26328\,
            I => \N__26302\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__26327\,
            I => \N__26296\
        );

    \I__5108\ : InMux
    port map (
            O => \N__26326\,
            I => \N__26293\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__26323\,
            I => \N__26290\
        );

    \I__5106\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26287\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__26317\,
            I => \N__26284\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__26310\,
            I => \N__26281\
        );

    \I__5103\ : CascadeMux
    port map (
            O => \N__26309\,
            I => \N__26277\
        );

    \I__5102\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26272\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__26305\,
            I => \N__26269\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26266\
        );

    \I__5099\ : InMux
    port map (
            O => \N__26301\,
            I => \N__26257\
        );

    \I__5098\ : InMux
    port map (
            O => \N__26300\,
            I => \N__26257\
        );

    \I__5097\ : InMux
    port map (
            O => \N__26299\,
            I => \N__26257\
        );

    \I__5096\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26257\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__26293\,
            I => \N__26254\
        );

    \I__5094\ : Span4Mux_v
    port map (
            O => \N__26290\,
            I => \N__26251\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26244\
        );

    \I__5092\ : Span4Mux_v
    port map (
            O => \N__26284\,
            I => \N__26244\
        );

    \I__5091\ : Span4Mux_h
    port map (
            O => \N__26281\,
            I => \N__26244\
        );

    \I__5090\ : InMux
    port map (
            O => \N__26280\,
            I => \N__26241\
        );

    \I__5089\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26238\
        );

    \I__5088\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26233\
        );

    \I__5087\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26233\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__26272\,
            I => \N__26228\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__26269\,
            I => \N__26228\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__26266\,
            I => \N__26221\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26221\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__26254\,
            I => \N__26221\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__26251\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__26244\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__26241\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__26238\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__26233\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__26228\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__26221\,
            I => \b2v_inst11.dutycycleZ0Z_5\
        );

    \I__5074\ : InMux
    port map (
            O => \N__26206\,
            I => \N__26203\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26200\
        );

    \I__5072\ : Odrv4
    port map (
            O => \N__26200\,
            I => \b2v_inst11.m6_0_1\
        );

    \I__5071\ : CascadeMux
    port map (
            O => \N__26197\,
            I => \N__26193\
        );

    \I__5070\ : CascadeMux
    port map (
            O => \N__26196\,
            I => \N__26185\
        );

    \I__5069\ : InMux
    port map (
            O => \N__26193\,
            I => \N__26180\
        );

    \I__5068\ : InMux
    port map (
            O => \N__26192\,
            I => \N__26171\
        );

    \I__5067\ : InMux
    port map (
            O => \N__26191\,
            I => \N__26171\
        );

    \I__5066\ : InMux
    port map (
            O => \N__26190\,
            I => \N__26171\
        );

    \I__5065\ : InMux
    port map (
            O => \N__26189\,
            I => \N__26168\
        );

    \I__5064\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26161\
        );

    \I__5063\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26158\
        );

    \I__5062\ : InMux
    port map (
            O => \N__26184\,
            I => \N__26148\
        );

    \I__5061\ : InMux
    port map (
            O => \N__26183\,
            I => \N__26148\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26145\
        );

    \I__5059\ : InMux
    port map (
            O => \N__26179\,
            I => \N__26140\
        );

    \I__5058\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26140\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26137\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__26168\,
            I => \N__26134\
        );

    \I__5055\ : InMux
    port map (
            O => \N__26167\,
            I => \N__26125\
        );

    \I__5054\ : InMux
    port map (
            O => \N__26166\,
            I => \N__26125\
        );

    \I__5053\ : InMux
    port map (
            O => \N__26165\,
            I => \N__26125\
        );

    \I__5052\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26125\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26122\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__26158\,
            I => \N__26119\
        );

    \I__5049\ : InMux
    port map (
            O => \N__26157\,
            I => \N__26116\
        );

    \I__5048\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26107\
        );

    \I__5047\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26107\
        );

    \I__5046\ : InMux
    port map (
            O => \N__26154\,
            I => \N__26107\
        );

    \I__5045\ : InMux
    port map (
            O => \N__26153\,
            I => \N__26107\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__26148\,
            I => \N__26104\
        );

    \I__5043\ : Span4Mux_v
    port map (
            O => \N__26145\,
            I => \N__26099\
        );

    \I__5042\ : LocalMux
    port map (
            O => \N__26140\,
            I => \N__26096\
        );

    \I__5041\ : Span4Mux_v
    port map (
            O => \N__26137\,
            I => \N__26087\
        );

    \I__5040\ : Span4Mux_v
    port map (
            O => \N__26134\,
            I => \N__26087\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__26125\,
            I => \N__26087\
        );

    \I__5038\ : Span4Mux_v
    port map (
            O => \N__26122\,
            I => \N__26087\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__26119\,
            I => \N__26084\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__26116\,
            I => \N__26077\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26077\
        );

    \I__5034\ : Span4Mux_h
    port map (
            O => \N__26104\,
            I => \N__26077\
        );

    \I__5033\ : InMux
    port map (
            O => \N__26103\,
            I => \N__26072\
        );

    \I__5032\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26072\
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__26099\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5030\ : Odrv12
    port map (
            O => \N__26096\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5029\ : Odrv4
    port map (
            O => \N__26087\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5028\ : Odrv4
    port map (
            O => \N__26084\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__26077\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__26072\,
            I => \b2v_inst11.dutycycleZ1Z_6\
        );

    \I__5025\ : InMux
    port map (
            O => \N__26059\,
            I => \N__26056\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__26056\,
            I => \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_0_1\
        );

    \I__5023\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26050\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__26047\
        );

    \I__5021\ : Span4Mux_h
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__26044\,
            I => \N_18\
        );

    \I__5019\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26038\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__26038\,
            I => \b2v_inst11.N_15_mux\
        );

    \I__5017\ : InMux
    port map (
            O => \N__26035\,
            I => \N__26032\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__26032\,
            I => \b2v_inst11.i6_mux_i_1\
        );

    \I__5015\ : InMux
    port map (
            O => \N__26029\,
            I => \N__26026\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__26026\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_11\
        );

    \I__5013\ : InMux
    port map (
            O => \N__26023\,
            I => \N__26017\
        );

    \I__5012\ : InMux
    port map (
            O => \N__26022\,
            I => \N__26017\
        );

    \I__5011\ : LocalMux
    port map (
            O => \N__26017\,
            I => \N__26014\
        );

    \I__5010\ : Span4Mux_h
    port map (
            O => \N__26014\,
            I => \N__26011\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__26011\,
            I => \b2v_inst11.dutycycle_RNI9R6T4Z0Z_12\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__26008\,
            I => \N__26005\
        );

    \I__5007\ : InMux
    port map (
            O => \N__26005\,
            I => \N__25999\
        );

    \I__5006\ : InMux
    port map (
            O => \N__26004\,
            I => \N__25999\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__5004\ : Odrv12
    port map (
            O => \N__25996\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5\
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__25993\,
            I => \N__25990\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25984\
        );

    \I__5001\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25984\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__25984\,
            I => \b2v_inst11.dutycycleZ1Z_12\
        );

    \I__4999\ : SRMux
    port map (
            O => \N__25981\,
            I => \N__25977\
        );

    \I__4998\ : SRMux
    port map (
            O => \N__25980\,
            I => \N__25973\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25977\,
            I => \N__25969\
        );

    \I__4996\ : SRMux
    port map (
            O => \N__25976\,
            I => \N__25966\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__25973\,
            I => \N__25963\
        );

    \I__4994\ : SRMux
    port map (
            O => \N__25972\,
            I => \N__25960\
        );

    \I__4993\ : Span4Mux_h
    port map (
            O => \N__25969\,
            I => \N__25955\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__25966\,
            I => \N__25955\
        );

    \I__4991\ : Span4Mux_h
    port map (
            O => \N__25963\,
            I => \N__25952\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__25960\,
            I => \N__25949\
        );

    \I__4989\ : Span4Mux_v
    port map (
            O => \N__25955\,
            I => \N__25938\
        );

    \I__4988\ : Span4Mux_h
    port map (
            O => \N__25952\,
            I => \N__25938\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__25949\,
            I => \N__25938\
        );

    \I__4986\ : SRMux
    port map (
            O => \N__25948\,
            I => \N__25934\
        );

    \I__4985\ : SRMux
    port map (
            O => \N__25947\,
            I => \N__25931\
        );

    \I__4984\ : SRMux
    port map (
            O => \N__25946\,
            I => \N__25928\
        );

    \I__4983\ : SRMux
    port map (
            O => \N__25945\,
            I => \N__25925\
        );

    \I__4982\ : Span4Mux_v
    port map (
            O => \N__25938\,
            I => \N__25922\
        );

    \I__4981\ : SRMux
    port map (
            O => \N__25937\,
            I => \N__25919\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__25934\,
            I => \N__25916\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__25931\,
            I => \N__25909\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__25928\,
            I => \N__25909\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__25925\,
            I => \N__25909\
        );

    \I__4976\ : IoSpan4Mux
    port map (
            O => \N__25922\,
            I => \N__25904\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25904\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__25916\,
            I => \N__25901\
        );

    \I__4973\ : Span4Mux_v
    port map (
            O => \N__25909\,
            I => \N__25898\
        );

    \I__4972\ : Span4Mux_s3_v
    port map (
            O => \N__25904\,
            I => \N__25894\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__25901\,
            I => \N__25891\
        );

    \I__4970\ : Sp12to4
    port map (
            O => \N__25898\,
            I => \N__25888\
        );

    \I__4969\ : SRMux
    port map (
            O => \N__25897\,
            I => \N__25885\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__25894\,
            I => \N__25882\
        );

    \I__4967\ : Odrv4
    port map (
            O => \N__25891\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__4966\ : Odrv12
    port map (
            O => \N__25888\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__25885\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__4964\ : Odrv4
    port map (
            O => \N__25882\,
            I => \b2v_inst11.N_224_iZ0\
        );

    \I__4963\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25867\
        );

    \I__4962\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25867\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__25867\,
            I => \b2v_inst11.dutycycleZ0Z_15\
        );

    \I__4960\ : InMux
    port map (
            O => \N__25864\,
            I => \N__25854\
        );

    \I__4959\ : InMux
    port map (
            O => \N__25863\,
            I => \N__25844\
        );

    \I__4958\ : InMux
    port map (
            O => \N__25862\,
            I => \N__25844\
        );

    \I__4957\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25844\
        );

    \I__4956\ : InMux
    port map (
            O => \N__25860\,
            I => \N__25844\
        );

    \I__4955\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25841\
        );

    \I__4954\ : InMux
    port map (
            O => \N__25858\,
            I => \N__25831\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__25857\,
            I => \N__25827\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25820\
        );

    \I__4951\ : CascadeMux
    port map (
            O => \N__25853\,
            I => \N__25812\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__25844\,
            I => \N__25808\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25805\
        );

    \I__4948\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25802\
        );

    \I__4947\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25789\
        );

    \I__4946\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25789\
        );

    \I__4945\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25789\
        );

    \I__4944\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25789\
        );

    \I__4943\ : InMux
    port map (
            O => \N__25835\,
            I => \N__25789\
        );

    \I__4942\ : InMux
    port map (
            O => \N__25834\,
            I => \N__25789\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__25831\,
            I => \N__25786\
        );

    \I__4940\ : InMux
    port map (
            O => \N__25830\,
            I => \N__25777\
        );

    \I__4939\ : InMux
    port map (
            O => \N__25827\,
            I => \N__25777\
        );

    \I__4938\ : InMux
    port map (
            O => \N__25826\,
            I => \N__25777\
        );

    \I__4937\ : InMux
    port map (
            O => \N__25825\,
            I => \N__25777\
        );

    \I__4936\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25772\
        );

    \I__4935\ : InMux
    port map (
            O => \N__25823\,
            I => \N__25772\
        );

    \I__4934\ : Span4Mux_v
    port map (
            O => \N__25820\,
            I => \N__25769\
        );

    \I__4933\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25758\
        );

    \I__4932\ : InMux
    port map (
            O => \N__25818\,
            I => \N__25758\
        );

    \I__4931\ : InMux
    port map (
            O => \N__25817\,
            I => \N__25758\
        );

    \I__4930\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25758\
        );

    \I__4929\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25758\
        );

    \I__4928\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25753\
        );

    \I__4927\ : InMux
    port map (
            O => \N__25811\,
            I => \N__25753\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__25808\,
            I => \N__25746\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__25805\,
            I => \N__25746\
        );

    \I__4924\ : LocalMux
    port map (
            O => \N__25802\,
            I => \N__25746\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__25789\,
            I => \N__25739\
        );

    \I__4922\ : Span12Mux_s6_v
    port map (
            O => \N__25786\,
            I => \N__25739\
        );

    \I__4921\ : LocalMux
    port map (
            O => \N__25777\,
            I => \N__25739\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__25772\,
            I => \N__25736\
        );

    \I__4919\ : Odrv4
    port map (
            O => \N__25769\,
            I => \func_state_RNIVS8U1_3_1\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__25758\,
            I => \func_state_RNIVS8U1_3_1\
        );

    \I__4917\ : LocalMux
    port map (
            O => \N__25753\,
            I => \func_state_RNIVS8U1_3_1\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__25746\,
            I => \func_state_RNIVS8U1_3_1\
        );

    \I__4915\ : Odrv12
    port map (
            O => \N__25739\,
            I => \func_state_RNIVS8U1_3_1\
        );

    \I__4914\ : Odrv4
    port map (
            O => \N__25736\,
            I => \func_state_RNIVS8U1_3_1\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \N__25720\
        );

    \I__4912\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25714\
        );

    \I__4911\ : InMux
    port map (
            O => \N__25719\,
            I => \N__25714\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__25714\,
            I => \N__25711\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__25711\,
            I => \N__25708\
        );

    \I__4908\ : Odrv4
    port map (
            O => \N__25708\,
            I => \b2v_inst11.dutycycle_en_12\
        );

    \I__4907\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25699\
        );

    \I__4906\ : InMux
    port map (
            O => \N__25704\,
            I => \N__25699\
        );

    \I__4905\ : LocalMux
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__25696\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\
        );

    \I__4903\ : InMux
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__25690\,
            I => \N__25687\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__4900\ : Odrv4
    port map (
            O => \N__25684\,
            I => \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_3_1\
        );

    \I__4899\ : CascadeMux
    port map (
            O => \N__25681\,
            I => \b2v_inst11.un1_dutycycle_53_50_1_i_i_1_cascade_\
        );

    \I__4898\ : CascadeMux
    port map (
            O => \N__25678\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\
        );

    \I__4897\ : InMux
    port map (
            O => \N__25675\,
            I => \N__25672\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__25672\,
            I => \b2v_inst11.mult1_un110_sum_i\
        );

    \I__4895\ : InMux
    port map (
            O => \N__25669\,
            I => \N__25666\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__25666\,
            I => \b2v_inst5.un12_clk_100khz_13\
        );

    \I__4893\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25660\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__25660\,
            I => \b2v_inst11.un1_dutycycle_53_axb_11\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__25657\,
            I => \b2v_inst11.i7_mux_cascade_\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__25654\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_11_cascade_\
        );

    \I__4889\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__25648\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_9\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__25645\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_8_cascade_\
        );

    \I__4886\ : InMux
    port map (
            O => \N__25642\,
            I => \N__25639\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__25639\,
            I => \b2v_inst11.mult1_un117_sum_cry_4_s\
        );

    \I__4884\ : InMux
    port map (
            O => \N__25636\,
            I => \b2v_inst11.mult1_un117_sum_cry_3\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__4882\ : InMux
    port map (
            O => \N__25630\,
            I => \N__25627\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__25627\,
            I => \b2v_inst11.mult1_un117_sum_cry_5_s\
        );

    \I__4880\ : InMux
    port map (
            O => \N__25624\,
            I => \b2v_inst11.mult1_un117_sum_cry_4\
        );

    \I__4879\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25618\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__25618\,
            I => \b2v_inst11.mult1_un117_sum_cry_6_s\
        );

    \I__4877\ : InMux
    port map (
            O => \N__25615\,
            I => \b2v_inst11.mult1_un117_sum_cry_5\
        );

    \I__4876\ : CascadeMux
    port map (
            O => \N__25612\,
            I => \N__25609\
        );

    \I__4875\ : InMux
    port map (
            O => \N__25609\,
            I => \N__25606\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__25606\,
            I => \b2v_inst11.mult1_un124_sum_axb_8\
        );

    \I__4873\ : InMux
    port map (
            O => \N__25603\,
            I => \b2v_inst11.mult1_un117_sum_cry_6\
        );

    \I__4872\ : InMux
    port map (
            O => \N__25600\,
            I => \b2v_inst11.mult1_un117_sum_cry_7\
        );

    \I__4871\ : CascadeMux
    port map (
            O => \N__25597\,
            I => \b2v_inst11.mult1_un117_sum_s_8_cascade_\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__25594\,
            I => \N__25590\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__25593\,
            I => \N__25586\
        );

    \I__4868\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25579\
        );

    \I__4867\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25579\
        );

    \I__4866\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25579\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__25579\,
            I => \b2v_inst11.mult1_un117_sum_i_0_8\
        );

    \I__4864\ : InMux
    port map (
            O => \N__25576\,
            I => \N__25573\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__25573\,
            I => \N__25570\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__25570\,
            I => \N__25566\
        );

    \I__4861\ : InMux
    port map (
            O => \N__25569\,
            I => \N__25563\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__25566\,
            I => \N__25560\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__25563\,
            I => \b2v_inst5.curr_stateZ0Z_1\
        );

    \I__4858\ : Odrv4
    port map (
            O => \N__25560\,
            I => \b2v_inst5.curr_stateZ0Z_1\
        );

    \I__4857\ : CascadeMux
    port map (
            O => \N__25555\,
            I => \N__25552\
        );

    \I__4856\ : InMux
    port map (
            O => \N__25552\,
            I => \N__25549\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__25549\,
            I => \N__25544\
        );

    \I__4854\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25539\
        );

    \I__4853\ : InMux
    port map (
            O => \N__25547\,
            I => \N__25539\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__25544\,
            I => \N__25534\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__25539\,
            I => \N__25534\
        );

    \I__4850\ : Span4Mux_v
    port map (
            O => \N__25534\,
            I => \N__25531\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__25531\,
            I => \N_413\
        );

    \I__4848\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25525\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__25525\,
            I => \b2v_inst11.mult1_un138_sum_axb_8\
        );

    \I__4846\ : InMux
    port map (
            O => \N__25522\,
            I => \b2v_inst11.mult1_un138_sum_cry_7\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__25519\,
            I => \N__25514\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__25518\,
            I => \N__25511\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__25517\,
            I => \N__25508\
        );

    \I__4842\ : InMux
    port map (
            O => \N__25514\,
            I => \N__25505\
        );

    \I__4841\ : InMux
    port map (
            O => \N__25511\,
            I => \N__25500\
        );

    \I__4840\ : InMux
    port map (
            O => \N__25508\,
            I => \N__25500\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__25505\,
            I => \b2v_inst11.mult1_un131_sum_i_0_8\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__25500\,
            I => \b2v_inst11.mult1_un131_sum_i_0_8\
        );

    \I__4837\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25492\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__25492\,
            I => \b2v_inst11.mult1_un117_sum_i\
        );

    \I__4835\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25486\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__25486\,
            I => \b2v_inst11.mult1_un131_sum_i\
        );

    \I__4833\ : CascadeMux
    port map (
            O => \N__25483\,
            I => \N__25479\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__25482\,
            I => \N__25476\
        );

    \I__4831\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25470\
        );

    \I__4830\ : InMux
    port map (
            O => \N__25476\,
            I => \N__25465\
        );

    \I__4829\ : InMux
    port map (
            O => \N__25475\,
            I => \N__25465\
        );

    \I__4828\ : InMux
    port map (
            O => \N__25474\,
            I => \N__25462\
        );

    \I__4827\ : InMux
    port map (
            O => \N__25473\,
            I => \N__25459\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__25470\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__25465\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__25462\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__25459\,
            I => \b2v_inst11.mult1_un131_sum_s_8\
        );

    \I__4822\ : InMux
    port map (
            O => \N__25450\,
            I => \N__25447\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__25447\,
            I => \b2v_inst11.mult1_un124_sum_i\
        );

    \I__4820\ : InMux
    port map (
            O => \N__25444\,
            I => \N__25441\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__25441\,
            I => \N__25438\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__25438\,
            I => \b2v_inst11.mult1_un145_sum_i\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__4816\ : InMux
    port map (
            O => \N__25432\,
            I => \N__25429\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__25429\,
            I => \b2v_inst11.mult1_un117_sum_cry_3_s\
        );

    \I__4814\ : InMux
    port map (
            O => \N__25426\,
            I => \b2v_inst11.mult1_un117_sum_cry_2\
        );

    \I__4813\ : InMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__25420\,
            I => \N__25417\
        );

    \I__4811\ : Odrv4
    port map (
            O => \N__25417\,
            I => \b2v_inst5.count_1_12\
        );

    \I__4810\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25411\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__25411\,
            I => \b2v_inst5.count_1_14\
        );

    \I__4808\ : InMux
    port map (
            O => \N__25408\,
            I => \b2v_inst11.mult1_un138_sum_cry_2\
        );

    \I__4807\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25402\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__25402\,
            I => \b2v_inst11.mult1_un131_sum_cry_3_s\
        );

    \I__4805\ : InMux
    port map (
            O => \N__25399\,
            I => \b2v_inst11.mult1_un138_sum_cry_3\
        );

    \I__4804\ : InMux
    port map (
            O => \N__25396\,
            I => \N__25393\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__25393\,
            I => \b2v_inst11.mult1_un131_sum_cry_4_s\
        );

    \I__4802\ : InMux
    port map (
            O => \N__25390\,
            I => \b2v_inst11.mult1_un138_sum_cry_4\
        );

    \I__4801\ : InMux
    port map (
            O => \N__25387\,
            I => \N__25384\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__25384\,
            I => \b2v_inst11.mult1_un131_sum_cry_5_s\
        );

    \I__4799\ : InMux
    port map (
            O => \N__25381\,
            I => \b2v_inst11.mult1_un138_sum_cry_5\
        );

    \I__4798\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25375\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__25375\,
            I => \b2v_inst11.mult1_un131_sum_cry_6_s\
        );

    \I__4796\ : InMux
    port map (
            O => \N__25372\,
            I => \b2v_inst11.mult1_un138_sum_cry_6\
        );

    \I__4795\ : CascadeMux
    port map (
            O => \N__25369\,
            I => \N__25366\
        );

    \I__4794\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25357\
        );

    \I__4793\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25357\
        );

    \I__4792\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25357\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__25357\,
            I => \b2v_inst36.N_2939_i\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__25354\,
            I => \N__25348\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__25353\,
            I => \N__25344\
        );

    \I__4788\ : CascadeMux
    port map (
            O => \N__25352\,
            I => \N__25341\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__25351\,
            I => \N__25337\
        );

    \I__4786\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25325\
        );

    \I__4785\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25325\
        );

    \I__4784\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25325\
        );

    \I__4783\ : InMux
    port map (
            O => \N__25341\,
            I => \N__25325\
        );

    \I__4782\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25325\
        );

    \I__4781\ : InMux
    port map (
            O => \N__25337\,
            I => \N__25320\
        );

    \I__4780\ : InMux
    port map (
            O => \N__25336\,
            I => \N__25320\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__25325\,
            I => \N__25317\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__25320\,
            I => \N__25314\
        );

    \I__4777\ : Span4Mux_h
    port map (
            O => \N__25317\,
            I => \N__25311\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__25314\,
            I => \N__25308\
        );

    \I__4775\ : Sp12to4
    port map (
            O => \N__25311\,
            I => \N__25305\
        );

    \I__4774\ : Span4Mux_v
    port map (
            O => \N__25308\,
            I => \N__25302\
        );

    \I__4773\ : Span12Mux_v
    port map (
            O => \N__25305\,
            I => \N__25299\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__25302\,
            I => \N__25296\
        );

    \I__4771\ : Odrv12
    port map (
            O => \N__25299\,
            I => \V33DSW_OK_c\
        );

    \I__4770\ : Odrv4
    port map (
            O => \N__25296\,
            I => \V33DSW_OK_c\
        );

    \I__4769\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25280\
        );

    \I__4768\ : InMux
    port map (
            O => \N__25290\,
            I => \N__25280\
        );

    \I__4767\ : InMux
    port map (
            O => \N__25289\,
            I => \N__25269\
        );

    \I__4766\ : InMux
    port map (
            O => \N__25288\,
            I => \N__25269\
        );

    \I__4765\ : InMux
    port map (
            O => \N__25287\,
            I => \N__25269\
        );

    \I__4764\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25269\
        );

    \I__4763\ : InMux
    port map (
            O => \N__25285\,
            I => \N__25269\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__25280\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__25269\,
            I => \b2v_inst36.curr_stateZ0Z_1\
        );

    \I__4760\ : CascadeMux
    port map (
            O => \N__25264\,
            I => \b2v_inst36.count_rst_7_cascade_\
        );

    \I__4759\ : CascadeMux
    port map (
            O => \N__25261\,
            I => \b2v_inst36.N_2942_i_cascade_\
        );

    \I__4758\ : InMux
    port map (
            O => \N__25258\,
            I => \N__25254\
        );

    \I__4757\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25251\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__25254\,
            I => \N__25246\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__25251\,
            I => \N__25246\
        );

    \I__4754\ : Span4Mux_h
    port map (
            O => \N__25246\,
            I => \N__25243\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__25243\,
            I => \b2v_inst200.countZ0Z_9\
        );

    \I__4752\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25234\
        );

    \I__4751\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25234\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__25234\,
            I => \N__25231\
        );

    \I__4749\ : Span4Mux_h
    port map (
            O => \N__25231\,
            I => \N__25228\
        );

    \I__4748\ : Odrv4
    port map (
            O => \N__25228\,
            I => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\
        );

    \I__4747\ : InMux
    port map (
            O => \N__25225\,
            I => \N__25222\
        );

    \I__4746\ : LocalMux
    port map (
            O => \N__25222\,
            I => \b2v_inst200.count_3_9\
        );

    \I__4745\ : InMux
    port map (
            O => \N__25219\,
            I => \N__25199\
        );

    \I__4744\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25192\
        );

    \I__4743\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25192\
        );

    \I__4742\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25192\
        );

    \I__4741\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25185\
        );

    \I__4740\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25185\
        );

    \I__4739\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25185\
        );

    \I__4738\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25178\
        );

    \I__4737\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25178\
        );

    \I__4736\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25178\
        );

    \I__4735\ : InMux
    port map (
            O => \N__25209\,
            I => \N__25169\
        );

    \I__4734\ : InMux
    port map (
            O => \N__25208\,
            I => \N__25169\
        );

    \I__4733\ : InMux
    port map (
            O => \N__25207\,
            I => \N__25169\
        );

    \I__4732\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25169\
        );

    \I__4731\ : InMux
    port map (
            O => \N__25205\,
            I => \N__25162\
        );

    \I__4730\ : InMux
    port map (
            O => \N__25204\,
            I => \N__25162\
        );

    \I__4729\ : InMux
    port map (
            O => \N__25203\,
            I => \N__25162\
        );

    \I__4728\ : InMux
    port map (
            O => \N__25202\,
            I => \N__25159\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__25199\,
            I => \N__25150\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__25192\,
            I => \N__25147\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__25185\,
            I => \N__25144\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__25178\,
            I => \N__25141\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__25169\,
            I => \N__25138\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__25162\,
            I => \N__25135\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__25159\,
            I => \N__25132\
        );

    \I__4720\ : CEMux
    port map (
            O => \N__25158\,
            I => \N__25105\
        );

    \I__4719\ : CEMux
    port map (
            O => \N__25157\,
            I => \N__25105\
        );

    \I__4718\ : CEMux
    port map (
            O => \N__25156\,
            I => \N__25105\
        );

    \I__4717\ : CEMux
    port map (
            O => \N__25155\,
            I => \N__25105\
        );

    \I__4716\ : CEMux
    port map (
            O => \N__25154\,
            I => \N__25105\
        );

    \I__4715\ : CEMux
    port map (
            O => \N__25153\,
            I => \N__25105\
        );

    \I__4714\ : Glb2LocalMux
    port map (
            O => \N__25150\,
            I => \N__25105\
        );

    \I__4713\ : Glb2LocalMux
    port map (
            O => \N__25147\,
            I => \N__25105\
        );

    \I__4712\ : Glb2LocalMux
    port map (
            O => \N__25144\,
            I => \N__25105\
        );

    \I__4711\ : Glb2LocalMux
    port map (
            O => \N__25141\,
            I => \N__25105\
        );

    \I__4710\ : Glb2LocalMux
    port map (
            O => \N__25138\,
            I => \N__25105\
        );

    \I__4709\ : Glb2LocalMux
    port map (
            O => \N__25135\,
            I => \N__25105\
        );

    \I__4708\ : Glb2LocalMux
    port map (
            O => \N__25132\,
            I => \N__25105\
        );

    \I__4707\ : GlobalMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__4706\ : gio2CtrlBuf
    port map (
            O => \N__25102\,
            I => \b2v_inst200.count_en_g\
        );

    \I__4705\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25096\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__25096\,
            I => \N__25093\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__25093\,
            I => \b2v_inst36.count_2_14\
        );

    \I__4702\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25087\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__25087\,
            I => \b2v_inst5.count_1_11\
        );

    \I__4700\ : CascadeMux
    port map (
            O => \N__25084\,
            I => \b2v_inst36.count_rst_3_cascade_\
        );

    \I__4699\ : CascadeMux
    port map (
            O => \N__25081\,
            I => \b2v_inst36.countZ0Z_11_cascade_\
        );

    \I__4698\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25075\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__25075\,
            I => \b2v_inst36.count_2_11\
        );

    \I__4696\ : CascadeMux
    port map (
            O => \N__25072\,
            I => \b2v_inst36.count_rst_12_cascade_\
        );

    \I__4695\ : CascadeMux
    port map (
            O => \N__25069\,
            I => \b2v_inst36.countZ0Z_2_cascade_\
        );

    \I__4694\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25063\
        );

    \I__4693\ : LocalMux
    port map (
            O => \N__25063\,
            I => \b2v_inst36.count_2_2\
        );

    \I__4692\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25057\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__25057\,
            I => \b2v_inst36.curr_state_7_1\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__25054\,
            I => \b2v_inst36.curr_stateZ0Z_1_cascade_\
        );

    \I__4689\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25048\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__25048\,
            I => \b2v_inst36.curr_state_0_1\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__25045\,
            I => \b2v_inst36.countZ0Z_1_cascade_\
        );

    \I__4686\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25039\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__25039\,
            I => \N__25036\
        );

    \I__4684\ : Odrv4
    port map (
            O => \N__25036\,
            I => \b2v_inst36.un12_clk_100khz_9\
        );

    \I__4683\ : CascadeMux
    port map (
            O => \N__25033\,
            I => \b2v_inst36.un12_clk_100khz_10_cascade_\
        );

    \I__4682\ : InMux
    port map (
            O => \N__25030\,
            I => \N__25027\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__25027\,
            I => \b2v_inst36.count_2_0\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__25024\,
            I => \b2v_inst36.countZ0Z_0_cascade_\
        );

    \I__4679\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__25018\,
            I => \b2v_inst36.count_rst_13\
        );

    \I__4677\ : CascadeMux
    port map (
            O => \N__25015\,
            I => \b2v_inst36.count_rst_13_cascade_\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__25012\,
            I => \b2v_inst36.un2_count_1_axb_1_cascade_\
        );

    \I__4675\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25003\
        );

    \I__4674\ : InMux
    port map (
            O => \N__25008\,
            I => \N__25003\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__25003\,
            I => \b2v_inst36.count_2_1\
        );

    \I__4672\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24997\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__24997\,
            I => \b2v_inst36.un12_clk_100khz_8\
        );

    \I__4670\ : InMux
    port map (
            O => \N__24994\,
            I => \N__24991\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__24991\,
            I => \b2v_inst36.count_rst_14\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__24988\,
            I => \N__24985\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24985\,
            I => \N__24979\
        );

    \I__4666\ : InMux
    port map (
            O => \N__24984\,
            I => \N__24979\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__24979\,
            I => \N__24976\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__24976\,
            I => \b2v_inst11.count_1_6\
        );

    \I__4663\ : InMux
    port map (
            O => \N__24973\,
            I => \N__24970\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__24970\,
            I => \b2v_inst11.count_0_6\
        );

    \I__4661\ : CascadeMux
    port map (
            O => \N__24967\,
            I => \N__24964\
        );

    \I__4660\ : InMux
    port map (
            O => \N__24964\,
            I => \N__24958\
        );

    \I__4659\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24958\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__24958\,
            I => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__24952\,
            I => \b2v_inst11.count_0_15\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__24949\,
            I => \b2v_inst11.pwm_out_en_cascade_\
        );

    \I__4654\ : IoInMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__24943\,
            I => \PWRBTN_LED_c\
        );

    \I__4652\ : InMux
    port map (
            O => \N__24940\,
            I => \N__24937\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__24937\,
            I => \b2v_inst11.pwm_out_1_sqmuxa_0\
        );

    \I__4650\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24928\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__24933\,
            I => \N__24925\
        );

    \I__4648\ : CascadeMux
    port map (
            O => \N__24932\,
            I => \N__24921\
        );

    \I__4647\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24917\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__24928\,
            I => \N__24914\
        );

    \I__4645\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24911\
        );

    \I__4644\ : InMux
    port map (
            O => \N__24924\,
            I => \N__24908\
        );

    \I__4643\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24905\
        );

    \I__4642\ : InMux
    port map (
            O => \N__24920\,
            I => \N__24902\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__24917\,
            I => \N__24895\
        );

    \I__4640\ : Span4Mux_h
    port map (
            O => \N__24914\,
            I => \N__24895\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24890\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__24908\,
            I => \N__24890\
        );

    \I__4637\ : LocalMux
    port map (
            O => \N__24905\,
            I => \N__24885\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__24902\,
            I => \N__24885\
        );

    \I__4635\ : InMux
    port map (
            O => \N__24901\,
            I => \N__24880\
        );

    \I__4634\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24880\
        );

    \I__4633\ : Span4Mux_v
    port map (
            O => \N__24895\,
            I => \N__24875\
        );

    \I__4632\ : Span4Mux_h
    port map (
            O => \N__24890\,
            I => \N__24875\
        );

    \I__4631\ : Span4Mux_h
    port map (
            O => \N__24885\,
            I => \N__24872\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__24880\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__24875\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__24872\,
            I => \SYNTHESIZED_WIRE_1keep_3_rep1\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__24865\,
            I => \N__24861\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__24864\,
            I => \N__24858\
        );

    \I__4625\ : InMux
    port map (
            O => \N__24861\,
            I => \N__24850\
        );

    \I__4624\ : InMux
    port map (
            O => \N__24858\,
            I => \N__24850\
        );

    \I__4623\ : InMux
    port map (
            O => \N__24857\,
            I => \N__24850\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__24850\,
            I => \N__24846\
        );

    \I__4621\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24842\
        );

    \I__4620\ : Span4Mux_v
    port map (
            O => \N__24846\,
            I => \N__24832\
        );

    \I__4619\ : InMux
    port map (
            O => \N__24845\,
            I => \N__24829\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__24842\,
            I => \N__24826\
        );

    \I__4617\ : InMux
    port map (
            O => \N__24841\,
            I => \N__24815\
        );

    \I__4616\ : InMux
    port map (
            O => \N__24840\,
            I => \N__24815\
        );

    \I__4615\ : InMux
    port map (
            O => \N__24839\,
            I => \N__24815\
        );

    \I__4614\ : InMux
    port map (
            O => \N__24838\,
            I => \N__24815\
        );

    \I__4613\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24815\
        );

    \I__4612\ : InMux
    port map (
            O => \N__24836\,
            I => \N__24810\
        );

    \I__4611\ : InMux
    port map (
            O => \N__24835\,
            I => \N__24810\
        );

    \I__4610\ : Span4Mux_v
    port map (
            O => \N__24832\,
            I => \N__24805\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__24829\,
            I => \N__24805\
        );

    \I__4608\ : Span4Mux_v
    port map (
            O => \N__24826\,
            I => \N__24802\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__24815\,
            I => \N__24797\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__24810\,
            I => \N__24797\
        );

    \I__4605\ : Span4Mux_h
    port map (
            O => \N__24805\,
            I => \N__24794\
        );

    \I__4604\ : Odrv4
    port map (
            O => \N__24802\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4603\ : Odrv12
    port map (
            O => \N__24797\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__24794\,
            I => \b2v_inst20_un4_counter_7_THRU_CO\
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__24787\,
            I => \N__24784\
        );

    \I__4600\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24778\
        );

    \I__4599\ : InMux
    port map (
            O => \N__24783\,
            I => \N__24778\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__24778\,
            I => \b2v_inst11.count_1_11\
        );

    \I__4597\ : InMux
    port map (
            O => \N__24775\,
            I => \b2v_inst11.un1_count_cry_10\
        );

    \I__4596\ : InMux
    port map (
            O => \N__24772\,
            I => \b2v_inst11.un1_count_cry_11\
        );

    \I__4595\ : InMux
    port map (
            O => \N__24769\,
            I => \b2v_inst11.un1_count_cry_12\
        );

    \I__4594\ : InMux
    port map (
            O => \N__24766\,
            I => \b2v_inst11.un1_count_cry_13\
        );

    \I__4593\ : InMux
    port map (
            O => \N__24763\,
            I => \b2v_inst11.un1_count_cry_14\
        );

    \I__4592\ : CascadeMux
    port map (
            O => \N__24760\,
            I => \N__24757\
        );

    \I__4591\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24751\
        );

    \I__4590\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24751\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__24751\,
            I => \N__24748\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__24748\,
            I => \b2v_inst11.count_1_5\
        );

    \I__4587\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24742\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__24742\,
            I => \b2v_inst11.count_0_5\
        );

    \I__4585\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24735\
        );

    \I__4584\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24732\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__24735\,
            I => \b2v_inst11.count_1_14\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__24732\,
            I => \b2v_inst11.count_1_14\
        );

    \I__4581\ : InMux
    port map (
            O => \N__24727\,
            I => \N__24724\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__24724\,
            I => \b2v_inst11.count_0_14\
        );

    \I__4579\ : CascadeMux
    port map (
            O => \N__24721\,
            I => \N__24717\
        );

    \I__4578\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24712\
        );

    \I__4577\ : InMux
    port map (
            O => \N__24717\,
            I => \N__24712\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__24712\,
            I => \N__24709\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__24709\,
            I => \b2v_inst11.count_1_2\
        );

    \I__4574\ : InMux
    port map (
            O => \N__24706\,
            I => \b2v_inst11.un1_count_cry_1\
        );

    \I__4573\ : InMux
    port map (
            O => \N__24703\,
            I => \b2v_inst11.un1_count_cry_2\
        );

    \I__4572\ : InMux
    port map (
            O => \N__24700\,
            I => \b2v_inst11.un1_count_cry_3\
        );

    \I__4571\ : InMux
    port map (
            O => \N__24697\,
            I => \b2v_inst11.un1_count_cry_4\
        );

    \I__4570\ : InMux
    port map (
            O => \N__24694\,
            I => \b2v_inst11.un1_count_cry_5\
        );

    \I__4569\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24685\
        );

    \I__4568\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24685\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__24685\,
            I => \N__24682\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__24682\,
            I => \b2v_inst11.count_1_7\
        );

    \I__4565\ : InMux
    port map (
            O => \N__24679\,
            I => \b2v_inst11.un1_count_cry_6\
        );

    \I__4564\ : InMux
    port map (
            O => \N__24676\,
            I => \b2v_inst11.un1_count_cry_7\
        );

    \I__4563\ : CascadeMux
    port map (
            O => \N__24673\,
            I => \N__24670\
        );

    \I__4562\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24664\
        );

    \I__4561\ : InMux
    port map (
            O => \N__24669\,
            I => \N__24664\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__24664\,
            I => \b2v_inst11.count_1_9\
        );

    \I__4559\ : InMux
    port map (
            O => \N__24661\,
            I => \bfn_7_14_0_\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__24658\,
            I => \N__24654\
        );

    \I__4557\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24649\
        );

    \I__4556\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24649\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__24649\,
            I => \b2v_inst11.count_1_10\
        );

    \I__4554\ : InMux
    port map (
            O => \N__24646\,
            I => \b2v_inst11.un1_count_cry_9\
        );

    \I__4553\ : InMux
    port map (
            O => \N__24643\,
            I => \N__24634\
        );

    \I__4552\ : InMux
    port map (
            O => \N__24642\,
            I => \N__24631\
        );

    \I__4551\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24626\
        );

    \I__4550\ : InMux
    port map (
            O => \N__24640\,
            I => \N__24626\
        );

    \I__4549\ : InMux
    port map (
            O => \N__24639\,
            I => \N__24623\
        );

    \I__4548\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24619\
        );

    \I__4547\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24616\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__24634\,
            I => \N__24607\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__24631\,
            I => \N__24607\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__24626\,
            I => \N__24607\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__24623\,
            I => \N__24607\
        );

    \I__4542\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24601\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__24619\,
            I => \N__24596\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__24616\,
            I => \N__24596\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__24607\,
            I => \N__24593\
        );

    \I__4538\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24588\
        );

    \I__4537\ : InMux
    port map (
            O => \N__24605\,
            I => \N__24588\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__24604\,
            I => \N__24583\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__24601\,
            I => \N__24577\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__24596\,
            I => \N__24574\
        );

    \I__4533\ : Sp12to4
    port map (
            O => \N__24593\,
            I => \N__24569\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__24588\,
            I => \N__24569\
        );

    \I__4531\ : InMux
    port map (
            O => \N__24587\,
            I => \N__24566\
        );

    \I__4530\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24563\
        );

    \I__4529\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24555\
        );

    \I__4528\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24555\
        );

    \I__4527\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24555\
        );

    \I__4526\ : InMux
    port map (
            O => \N__24580\,
            I => \N__24552\
        );

    \I__4525\ : Sp12to4
    port map (
            O => \N__24577\,
            I => \N__24549\
        );

    \I__4524\ : Span4Mux_v
    port map (
            O => \N__24574\,
            I => \N__24546\
        );

    \I__4523\ : Span12Mux_s4_h
    port map (
            O => \N__24569\,
            I => \N__24539\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__24566\,
            I => \N__24539\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__24563\,
            I => \N__24539\
        );

    \I__4520\ : InMux
    port map (
            O => \N__24562\,
            I => \N__24536\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24531\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__24552\,
            I => \N__24531\
        );

    \I__4517\ : Odrv12
    port map (
            O => \N__24549\,
            I => \GPIO_FPGA_SoC_4_c\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__24546\,
            I => \GPIO_FPGA_SoC_4_c\
        );

    \I__4515\ : Odrv12
    port map (
            O => \N__24539\,
            I => \GPIO_FPGA_SoC_4_c\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__24536\,
            I => \GPIO_FPGA_SoC_4_c\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__24531\,
            I => \GPIO_FPGA_SoC_4_c\
        );

    \I__4512\ : CascadeMux
    port map (
            O => \N__24520\,
            I => \N__24516\
        );

    \I__4511\ : CascadeMux
    port map (
            O => \N__24519\,
            I => \N__24507\
        );

    \I__4510\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24504\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__24515\,
            I => \N__24501\
        );

    \I__4508\ : InMux
    port map (
            O => \N__24514\,
            I => \N__24497\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__24513\,
            I => \N__24494\
        );

    \I__4506\ : InMux
    port map (
            O => \N__24512\,
            I => \N__24491\
        );

    \I__4505\ : InMux
    port map (
            O => \N__24511\,
            I => \N__24488\
        );

    \I__4504\ : InMux
    port map (
            O => \N__24510\,
            I => \N__24485\
        );

    \I__4503\ : InMux
    port map (
            O => \N__24507\,
            I => \N__24481\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__24504\,
            I => \N__24478\
        );

    \I__4501\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24473\
        );

    \I__4500\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24473\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24470\
        );

    \I__4498\ : InMux
    port map (
            O => \N__24494\,
            I => \N__24466\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__24491\,
            I => \N__24461\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__24488\,
            I => \N__24461\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__24485\,
            I => \N__24458\
        );

    \I__4494\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24455\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__24481\,
            I => \N__24452\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__24478\,
            I => \N__24449\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__24473\,
            I => \N__24446\
        );

    \I__4490\ : Span4Mux_v
    port map (
            O => \N__24470\,
            I => \N__24443\
        );

    \I__4489\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24440\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24437\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__24461\,
            I => \N__24434\
        );

    \I__4486\ : Span4Mux_s2_v
    port map (
            O => \N__24458\,
            I => \N__24429\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__24455\,
            I => \N__24429\
        );

    \I__4484\ : Span4Mux_v
    port map (
            O => \N__24452\,
            I => \N__24426\
        );

    \I__4483\ : Span4Mux_v
    port map (
            O => \N__24449\,
            I => \N__24415\
        );

    \I__4482\ : Span4Mux_s2_h
    port map (
            O => \N__24446\,
            I => \N__24415\
        );

    \I__4481\ : Span4Mux_h
    port map (
            O => \N__24443\,
            I => \N__24415\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24415\
        );

    \I__4479\ : Span4Mux_h
    port map (
            O => \N__24437\,
            I => \N__24415\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__24434\,
            I => \N__24410\
        );

    \I__4477\ : Span4Mux_v
    port map (
            O => \N__24429\,
            I => \N__24410\
        );

    \I__4476\ : Span4Mux_s2_h
    port map (
            O => \N__24426\,
            I => \N__24405\
        );

    \I__4475\ : Span4Mux_v
    port map (
            O => \N__24415\,
            I => \N__24405\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__24410\,
            I => \N_161\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__24405\,
            I => \N_161\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__24400\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\
        );

    \I__4471\ : InMux
    port map (
            O => \N__24397\,
            I => \N__24376\
        );

    \I__4470\ : InMux
    port map (
            O => \N__24396\,
            I => \N__24376\
        );

    \I__4469\ : InMux
    port map (
            O => \N__24395\,
            I => \N__24376\
        );

    \I__4468\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24376\
        );

    \I__4467\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24376\
        );

    \I__4466\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24371\
        );

    \I__4465\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24371\
        );

    \I__4464\ : InMux
    port map (
            O => \N__24390\,
            I => \N__24367\
        );

    \I__4463\ : InMux
    port map (
            O => \N__24389\,
            I => \N__24362\
        );

    \I__4462\ : InMux
    port map (
            O => \N__24388\,
            I => \N__24358\
        );

    \I__4461\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24355\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__24376\,
            I => \N__24350\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__24371\,
            I => \N__24350\
        );

    \I__4458\ : InMux
    port map (
            O => \N__24370\,
            I => \N__24347\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__24367\,
            I => \N__24344\
        );

    \I__4456\ : InMux
    port map (
            O => \N__24366\,
            I => \N__24341\
        );

    \I__4455\ : InMux
    port map (
            O => \N__24365\,
            I => \N__24338\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__24362\,
            I => \N__24335\
        );

    \I__4453\ : InMux
    port map (
            O => \N__24361\,
            I => \N__24332\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__24358\,
            I => \N__24325\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__24355\,
            I => \N__24320\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__24350\,
            I => \N__24320\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__24347\,
            I => \N__24314\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__24344\,
            I => \N__24309\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__24341\,
            I => \N__24309\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__24338\,
            I => \N__24305\
        );

    \I__4445\ : Span4Mux_v
    port map (
            O => \N__24335\,
            I => \N__24300\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24300\
        );

    \I__4443\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24297\
        );

    \I__4442\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24290\
        );

    \I__4441\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24290\
        );

    \I__4440\ : InMux
    port map (
            O => \N__24328\,
            I => \N__24290\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__24325\,
            I => \N__24285\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__24320\,
            I => \N__24285\
        );

    \I__4437\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24278\
        );

    \I__4436\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24278\
        );

    \I__4435\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24278\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__24314\,
            I => \N__24275\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__24309\,
            I => \N__24272\
        );

    \I__4432\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24269\
        );

    \I__4431\ : Span4Mux_v
    port map (
            O => \N__24305\,
            I => \N__24266\
        );

    \I__4430\ : Span4Mux_h
    port map (
            O => \N__24300\,
            I => \N__24259\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__24297\,
            I => \N__24259\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__24290\,
            I => \N__24259\
        );

    \I__4427\ : Span4Mux_v
    port map (
            O => \N__24285\,
            I => \N__24254\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__24278\,
            I => \N__24254\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__24275\,
            I => \N__24251\
        );

    \I__4424\ : Span4Mux_v
    port map (
            O => \N__24272\,
            I => \N__24246\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__24269\,
            I => \N__24246\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__24266\,
            I => \N__24241\
        );

    \I__4421\ : Span4Mux_v
    port map (
            O => \N__24259\,
            I => \N__24241\
        );

    \I__4420\ : Span4Mux_h
    port map (
            O => \N__24254\,
            I => \N__24238\
        );

    \I__4419\ : Span4Mux_h
    port map (
            O => \N__24251\,
            I => \N__24233\
        );

    \I__4418\ : Span4Mux_h
    port map (
            O => \N__24246\,
            I => \N__24233\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__24241\,
            I => \SLP_S3n_c\
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__24238\,
            I => \SLP_S3n_c\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__24233\,
            I => \SLP_S3n_c\
        );

    \I__4414\ : InMux
    port map (
            O => \N__24226\,
            I => \N__24223\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__24223\,
            I => \N__24220\
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__24220\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIZ0\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__24217\,
            I => \N__24214\
        );

    \I__4410\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24208\
        );

    \I__4409\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24205\
        );

    \I__4408\ : InMux
    port map (
            O => \N__24212\,
            I => \N__24202\
        );

    \I__4407\ : InMux
    port map (
            O => \N__24211\,
            I => \N__24199\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__24208\,
            I => \N__24196\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__24205\,
            I => \N__24191\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24191\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__24199\,
            I => \N__24187\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__24196\,
            I => \N__24184\
        );

    \I__4401\ : Span4Mux_v
    port map (
            O => \N__24191\,
            I => \N__24181\
        );

    \I__4400\ : InMux
    port map (
            O => \N__24190\,
            I => \N__24178\
        );

    \I__4399\ : Span4Mux_s3_h
    port map (
            O => \N__24187\,
            I => \N__24175\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__24184\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__24181\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__24178\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__24175\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1\
        );

    \I__4394\ : CascadeMux
    port map (
            O => \N__24166\,
            I => \N__24163\
        );

    \I__4393\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24156\
        );

    \I__4392\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24156\
        );

    \I__4391\ : CascadeMux
    port map (
            O => \N__24161\,
            I => \N__24152\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__24156\,
            I => \N__24145\
        );

    \I__4389\ : InMux
    port map (
            O => \N__24155\,
            I => \N__24142\
        );

    \I__4388\ : InMux
    port map (
            O => \N__24152\,
            I => \N__24133\
        );

    \I__4387\ : InMux
    port map (
            O => \N__24151\,
            I => \N__24133\
        );

    \I__4386\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24133\
        );

    \I__4385\ : InMux
    port map (
            O => \N__24149\,
            I => \N__24133\
        );

    \I__4384\ : CascadeMux
    port map (
            O => \N__24148\,
            I => \N__24129\
        );

    \I__4383\ : Span4Mux_s3_h
    port map (
            O => \N__24145\,
            I => \N__24120\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__24142\,
            I => \N__24120\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__24133\,
            I => \N__24117\
        );

    \I__4380\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24114\
        );

    \I__4379\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24108\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__24128\,
            I => \N__24105\
        );

    \I__4377\ : InMux
    port map (
            O => \N__24127\,
            I => \N__24097\
        );

    \I__4376\ : InMux
    port map (
            O => \N__24126\,
            I => \N__24094\
        );

    \I__4375\ : InMux
    port map (
            O => \N__24125\,
            I => \N__24091\
        );

    \I__4374\ : Span4Mux_h
    port map (
            O => \N__24120\,
            I => \N__24086\
        );

    \I__4373\ : Span4Mux_s3_h
    port map (
            O => \N__24117\,
            I => \N__24086\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__24114\,
            I => \N__24083\
        );

    \I__4371\ : InMux
    port map (
            O => \N__24113\,
            I => \N__24076\
        );

    \I__4370\ : InMux
    port map (
            O => \N__24112\,
            I => \N__24076\
        );

    \I__4369\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24076\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24073\
        );

    \I__4367\ : InMux
    port map (
            O => \N__24105\,
            I => \N__24066\
        );

    \I__4366\ : InMux
    port map (
            O => \N__24104\,
            I => \N__24066\
        );

    \I__4365\ : InMux
    port map (
            O => \N__24103\,
            I => \N__24066\
        );

    \I__4364\ : InMux
    port map (
            O => \N__24102\,
            I => \N__24063\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__24101\,
            I => \N__24060\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__24100\,
            I => \N__24057\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__24097\,
            I => \N__24053\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__24094\,
            I => \N__24047\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__24091\,
            I => \N__24047\
        );

    \I__4358\ : Span4Mux_v
    port map (
            O => \N__24086\,
            I => \N__24040\
        );

    \I__4357\ : Span4Mux_s3_h
    port map (
            O => \N__24083\,
            I => \N__24040\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__24076\,
            I => \N__24040\
        );

    \I__4355\ : Span4Mux_s3_h
    port map (
            O => \N__24073\,
            I => \N__24035\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__24066\,
            I => \N__24035\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24032\
        );

    \I__4352\ : InMux
    port map (
            O => \N__24060\,
            I => \N__24029\
        );

    \I__4351\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24026\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__24056\,
            I => \N__24022\
        );

    \I__4349\ : Span4Mux_s3_h
    port map (
            O => \N__24053\,
            I => \N__24018\
        );

    \I__4348\ : InMux
    port map (
            O => \N__24052\,
            I => \N__24015\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__24047\,
            I => \N__24012\
        );

    \I__4346\ : Span4Mux_h
    port map (
            O => \N__24040\,
            I => \N__24009\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__24035\,
            I => \N__24000\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__24032\,
            I => \N__24000\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__24029\,
            I => \N__24000\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__24026\,
            I => \N__24000\
        );

    \I__4341\ : InMux
    port map (
            O => \N__24025\,
            I => \N__23995\
        );

    \I__4340\ : InMux
    port map (
            O => \N__24022\,
            I => \N__23995\
        );

    \I__4339\ : InMux
    port map (
            O => \N__24021\,
            I => \N__23992\
        );

    \I__4338\ : Sp12to4
    port map (
            O => \N__24018\,
            I => \N__23986\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__23986\
        );

    \I__4336\ : Span4Mux_v
    port map (
            O => \N__24012\,
            I => \N__23983\
        );

    \I__4335\ : Span4Mux_v
    port map (
            O => \N__24009\,
            I => \N__23980\
        );

    \I__4334\ : Span4Mux_v
    port map (
            O => \N__24000\,
            I => \N__23975\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__23995\,
            I => \N__23975\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__23992\,
            I => \N__23972\
        );

    \I__4331\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23969\
        );

    \I__4330\ : Odrv12
    port map (
            O => \N__23986\,
            I => \SLP_S4n_c\
        );

    \I__4329\ : Odrv4
    port map (
            O => \N__23983\,
            I => \SLP_S4n_c\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__23980\,
            I => \SLP_S4n_c\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__23975\,
            I => \SLP_S4n_c\
        );

    \I__4326\ : Odrv12
    port map (
            O => \N__23972\,
            I => \SLP_S4n_c\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__23969\,
            I => \SLP_S4n_c\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__23956\,
            I => \b2v_inst11.g1_0_0_cascade_\
        );

    \I__4323\ : InMux
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__23950\,
            I => \b2v_inst11.N_295\
        );

    \I__4321\ : CascadeMux
    port map (
            O => \N__23947\,
            I => \N__23944\
        );

    \I__4320\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23941\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__23941\,
            I => \b2v_inst11.g1\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__23938\,
            I => \b2v_inst11.g1_cascade_\
        );

    \I__4317\ : InMux
    port map (
            O => \N__23935\,
            I => \N__23929\
        );

    \I__4316\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23929\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23926\
        );

    \I__4314\ : Span4Mux_v
    port map (
            O => \N__23926\,
            I => \N__23923\
        );

    \I__4313\ : Odrv4
    port map (
            O => \N__23923\,
            I => \b2v_inst11.g1_0\
        );

    \I__4312\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23914\
        );

    \I__4311\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23914\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__23914\,
            I => \b2v_inst11.dutycycleZ0Z_2\
        );

    \I__4309\ : IoInMux
    port map (
            O => \N__23911\,
            I => \N__23908\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__23908\,
            I => \N__23900\
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__23907\,
            I => \N__23896\
        );

    \I__4306\ : CascadeMux
    port map (
            O => \N__23906\,
            I => \N__23891\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__23905\,
            I => \N__23888\
        );

    \I__4304\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23881\
        );

    \I__4303\ : InMux
    port map (
            O => \N__23903\,
            I => \N__23881\
        );

    \I__4302\ : IoSpan4Mux
    port map (
            O => \N__23900\,
            I => \N__23871\
        );

    \I__4301\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23866\
        );

    \I__4300\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23866\
        );

    \I__4299\ : InMux
    port map (
            O => \N__23895\,
            I => \N__23861\
        );

    \I__4298\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23861\
        );

    \I__4297\ : InMux
    port map (
            O => \N__23891\,
            I => \N__23858\
        );

    \I__4296\ : InMux
    port map (
            O => \N__23888\,
            I => \N__23854\
        );

    \I__4295\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23847\
        );

    \I__4294\ : InMux
    port map (
            O => \N__23886\,
            I => \N__23847\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__23881\,
            I => \N__23844\
        );

    \I__4292\ : InMux
    port map (
            O => \N__23880\,
            I => \N__23841\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23879\,
            I => \N__23838\
        );

    \I__4290\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23830\
        );

    \I__4289\ : InMux
    port map (
            O => \N__23877\,
            I => \N__23830\
        );

    \I__4288\ : InMux
    port map (
            O => \N__23876\,
            I => \N__23825\
        );

    \I__4287\ : InMux
    port map (
            O => \N__23875\,
            I => \N__23825\
        );

    \I__4286\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23822\
        );

    \I__4285\ : Span4Mux_s0_h
    port map (
            O => \N__23871\,
            I => \N__23817\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__23866\,
            I => \N__23817\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__23861\,
            I => \N__23812\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__23858\,
            I => \N__23812\
        );

    \I__4281\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23809\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__23854\,
            I => \N__23806\
        );

    \I__4279\ : InMux
    port map (
            O => \N__23853\,
            I => \N__23803\
        );

    \I__4278\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23800\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__23847\,
            I => \N__23793\
        );

    \I__4276\ : Span4Mux_v
    port map (
            O => \N__23844\,
            I => \N__23793\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__23841\,
            I => \N__23793\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__23838\,
            I => \N__23789\
        );

    \I__4273\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23782\
        );

    \I__4272\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23782\
        );

    \I__4271\ : InMux
    port map (
            O => \N__23835\,
            I => \N__23782\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23779\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__23825\,
            I => \N__23776\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__23822\,
            I => \N__23767\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__23817\,
            I => \N__23767\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__23812\,
            I => \N__23767\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__23809\,
            I => \N__23767\
        );

    \I__4264\ : Span4Mux_v
    port map (
            O => \N__23806\,
            I => \N__23758\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__23803\,
            I => \N__23758\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23758\
        );

    \I__4261\ : Span4Mux_h
    port map (
            O => \N__23793\,
            I => \N__23758\
        );

    \I__4260\ : InMux
    port map (
            O => \N__23792\,
            I => \N__23754\
        );

    \I__4259\ : Span4Mux_v
    port map (
            O => \N__23789\,
            I => \N__23751\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__23782\,
            I => \N__23748\
        );

    \I__4257\ : Span4Mux_h
    port map (
            O => \N__23779\,
            I => \N__23745\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__23776\,
            I => \N__23738\
        );

    \I__4255\ : Span4Mux_v
    port map (
            O => \N__23767\,
            I => \N__23738\
        );

    \I__4254\ : Span4Mux_v
    port map (
            O => \N__23758\,
            I => \N__23738\
        );

    \I__4253\ : InMux
    port map (
            O => \N__23757\,
            I => \N__23735\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__23754\,
            I => \RSMRSTn_fast_RNIGMH81\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__23751\,
            I => \RSMRSTn_fast_RNIGMH81\
        );

    \I__4250\ : Odrv12
    port map (
            O => \N__23748\,
            I => \RSMRSTn_fast_RNIGMH81\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__23745\,
            I => \RSMRSTn_fast_RNIGMH81\
        );

    \I__4248\ : Odrv4
    port map (
            O => \N__23738\,
            I => \RSMRSTn_fast_RNIGMH81\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__23735\,
            I => \RSMRSTn_fast_RNIGMH81\
        );

    \I__4246\ : InMux
    port map (
            O => \N__23722\,
            I => \N__23717\
        );

    \I__4245\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23711\
        );

    \I__4244\ : CascadeMux
    port map (
            O => \N__23720\,
            I => \N__23706\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23690\
        );

    \I__4242\ : InMux
    port map (
            O => \N__23716\,
            I => \N__23687\
        );

    \I__4241\ : InMux
    port map (
            O => \N__23715\,
            I => \N__23684\
        );

    \I__4240\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23681\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__23711\,
            I => \N__23678\
        );

    \I__4238\ : InMux
    port map (
            O => \N__23710\,
            I => \N__23673\
        );

    \I__4237\ : InMux
    port map (
            O => \N__23709\,
            I => \N__23673\
        );

    \I__4236\ : InMux
    port map (
            O => \N__23706\,
            I => \N__23664\
        );

    \I__4235\ : InMux
    port map (
            O => \N__23705\,
            I => \N__23664\
        );

    \I__4234\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23664\
        );

    \I__4233\ : InMux
    port map (
            O => \N__23703\,
            I => \N__23657\
        );

    \I__4232\ : InMux
    port map (
            O => \N__23702\,
            I => \N__23657\
        );

    \I__4231\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23657\
        );

    \I__4230\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23650\
        );

    \I__4229\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23650\
        );

    \I__4228\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23647\
        );

    \I__4227\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23640\
        );

    \I__4226\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23640\
        );

    \I__4225\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23640\
        );

    \I__4224\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23633\
        );

    \I__4223\ : InMux
    port map (
            O => \N__23693\,
            I => \N__23633\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__23690\,
            I => \N__23619\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__23687\,
            I => \N__23619\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__23684\,
            I => \N__23619\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__23681\,
            I => \N__23619\
        );

    \I__4218\ : Span4Mux_v
    port map (
            O => \N__23678\,
            I => \N__23619\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__23673\,
            I => \N__23619\
        );

    \I__4216\ : InMux
    port map (
            O => \N__23672\,
            I => \N__23612\
        );

    \I__4215\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23612\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__23664\,
            I => \N__23607\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__23657\,
            I => \N__23607\
        );

    \I__4212\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23602\
        );

    \I__4211\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23602\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23599\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__23647\,
            I => \N__23596\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23593\
        );

    \I__4207\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23588\
        );

    \I__4206\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23588\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__23633\,
            I => \N__23584\
        );

    \I__4204\ : InMux
    port map (
            O => \N__23632\,
            I => \N__23581\
        );

    \I__4203\ : Span4Mux_v
    port map (
            O => \N__23619\,
            I => \N__23578\
        );

    \I__4202\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23573\
        );

    \I__4201\ : InMux
    port map (
            O => \N__23617\,
            I => \N__23573\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__23612\,
            I => \N__23568\
        );

    \I__4199\ : Span12Mux_s11_v
    port map (
            O => \N__23607\,
            I => \N__23568\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__23602\,
            I => \N__23563\
        );

    \I__4197\ : Span4Mux_s3_h
    port map (
            O => \N__23599\,
            I => \N__23563\
        );

    \I__4196\ : Span4Mux_s3_h
    port map (
            O => \N__23596\,
            I => \N__23560\
        );

    \I__4195\ : Span4Mux_s3_h
    port map (
            O => \N__23593\,
            I => \N__23555\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__23588\,
            I => \N__23555\
        );

    \I__4193\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23552\
        );

    \I__4192\ : Odrv12
    port map (
            O => \N__23584\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__23581\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4190\ : Odrv4
    port map (
            O => \N__23578\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__23573\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4188\ : Odrv12
    port map (
            O => \N__23568\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4187\ : Odrv4
    port map (
            O => \N__23563\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4186\ : Odrv4
    port map (
            O => \N__23560\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4185\ : Odrv4
    port map (
            O => \N__23555\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__23552\,
            I => \func_state_RNI6BE8E_0_1\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__23533\,
            I => \N__23528\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__23532\,
            I => \N__23525\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__23531\,
            I => \N__23522\
        );

    \I__4180\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23514\
        );

    \I__4179\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23514\
        );

    \I__4178\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23511\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__23521\,
            I => \N__23506\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__23520\,
            I => \N__23503\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__23519\,
            I => \N__23500\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23496\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__23511\,
            I => \N__23493\
        );

    \I__4172\ : InMux
    port map (
            O => \N__23510\,
            I => \N__23490\
        );

    \I__4171\ : InMux
    port map (
            O => \N__23509\,
            I => \N__23487\
        );

    \I__4170\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23484\
        );

    \I__4169\ : InMux
    port map (
            O => \N__23503\,
            I => \N__23479\
        );

    \I__4168\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23476\
        );

    \I__4167\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23473\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__23496\,
            I => \N__23469\
        );

    \I__4165\ : Span4Mux_h
    port map (
            O => \N__23493\,
            I => \N__23462\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__23490\,
            I => \N__23462\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__23487\,
            I => \N__23462\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__23484\,
            I => \N__23459\
        );

    \I__4161\ : InMux
    port map (
            O => \N__23483\,
            I => \N__23456\
        );

    \I__4160\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23453\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23447\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__23476\,
            I => \N__23447\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__23473\,
            I => \N__23444\
        );

    \I__4156\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23441\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__23469\,
            I => \N__23430\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__23462\,
            I => \N__23430\
        );

    \I__4153\ : Span4Mux_v
    port map (
            O => \N__23459\,
            I => \N__23430\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__23456\,
            I => \N__23430\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__23453\,
            I => \N__23430\
        );

    \I__4150\ : InMux
    port map (
            O => \N__23452\,
            I => \N__23427\
        );

    \I__4149\ : Span4Mux_h
    port map (
            O => \N__23447\,
            I => \N__23423\
        );

    \I__4148\ : Span4Mux_h
    port map (
            O => \N__23444\,
            I => \N__23420\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23417\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__23430\,
            I => \N__23414\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__23427\,
            I => \N__23411\
        );

    \I__4144\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23408\
        );

    \I__4143\ : Odrv4
    port map (
            O => \N__23423\,
            I => b2v_inst11_dutycycle_1_0_iv_0_o3_out
        );

    \I__4142\ : Odrv4
    port map (
            O => \N__23420\,
            I => b2v_inst11_dutycycle_1_0_iv_0_o3_out
        );

    \I__4141\ : Odrv12
    port map (
            O => \N__23417\,
            I => b2v_inst11_dutycycle_1_0_iv_0_o3_out
        );

    \I__4140\ : Odrv4
    port map (
            O => \N__23414\,
            I => b2v_inst11_dutycycle_1_0_iv_0_o3_out
        );

    \I__4139\ : Odrv12
    port map (
            O => \N__23411\,
            I => b2v_inst11_dutycycle_1_0_iv_0_o3_out
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__23408\,
            I => b2v_inst11_dutycycle_1_0_iv_0_o3_out
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__4136\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23383\
        );

    \I__4135\ : InMux
    port map (
            O => \N__23391\,
            I => \N__23383\
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__23390\,
            I => \N__23377\
        );

    \I__4133\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23370\
        );

    \I__4132\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23370\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__23383\,
            I => \N__23367\
        );

    \I__4130\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23360\
        );

    \I__4129\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23360\
        );

    \I__4128\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23357\
        );

    \I__4127\ : InMux
    port map (
            O => \N__23377\,
            I => \N__23353\
        );

    \I__4126\ : InMux
    port map (
            O => \N__23376\,
            I => \N__23350\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__23375\,
            I => \N__23346\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__23370\,
            I => \N__23343\
        );

    \I__4123\ : Span4Mux_v
    port map (
            O => \N__23367\,
            I => \N__23340\
        );

    \I__4122\ : InMux
    port map (
            O => \N__23366\,
            I => \N__23335\
        );

    \I__4121\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23335\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__23360\,
            I => \N__23332\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__23357\,
            I => \N__23329\
        );

    \I__4118\ : InMux
    port map (
            O => \N__23356\,
            I => \N__23326\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23323\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__23350\,
            I => \N__23319\
        );

    \I__4115\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23316\
        );

    \I__4114\ : InMux
    port map (
            O => \N__23346\,
            I => \N__23313\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__23343\,
            I => \N__23310\
        );

    \I__4112\ : Span4Mux_h
    port map (
            O => \N__23340\,
            I => \N__23305\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__23335\,
            I => \N__23305\
        );

    \I__4110\ : Span4Mux_s3_h
    port map (
            O => \N__23332\,
            I => \N__23298\
        );

    \I__4109\ : Span4Mux_h
    port map (
            O => \N__23329\,
            I => \N__23298\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__23326\,
            I => \N__23298\
        );

    \I__4107\ : Span4Mux_s3_h
    port map (
            O => \N__23323\,
            I => \N__23295\
        );

    \I__4106\ : InMux
    port map (
            O => \N__23322\,
            I => \N__23292\
        );

    \I__4105\ : Odrv12
    port map (
            O => \N__23319\,
            I => \func_state_RNI_4_0\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__23316\,
            I => \func_state_RNI_4_0\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__23313\,
            I => \func_state_RNI_4_0\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__23310\,
            I => \func_state_RNI_4_0\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__23305\,
            I => \func_state_RNI_4_0\
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__23298\,
            I => \func_state_RNI_4_0\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__23295\,
            I => \func_state_RNI_4_0\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__23292\,
            I => \func_state_RNI_4_0\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__23275\,
            I => \N__23272\
        );

    \I__4096\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23266\
        );

    \I__4095\ : InMux
    port map (
            O => \N__23271\,
            I => \N__23266\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__23266\,
            I => \b2v_inst11.dutycycleZ0Z_13\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__23263\,
            I => \b2v_inst11.dutycycleZ0Z_5_cascade_\
        );

    \I__4092\ : InMux
    port map (
            O => \N__23260\,
            I => \N__23256\
        );

    \I__4091\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23253\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23248\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__23253\,
            I => \N__23248\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__23248\,
            I => \N__23245\
        );

    \I__4087\ : Odrv4
    port map (
            O => \N__23245\,
            I => \b2v_inst11.N_326_N\
        );

    \I__4086\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__4085\ : InMux
    port map (
            O => \N__23241\,
            I => \N__23236\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23226\
        );

    \I__4083\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23221\
        );

    \I__4082\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23221\
        );

    \I__4081\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23216\
        );

    \I__4080\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23216\
        );

    \I__4079\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23211\
        );

    \I__4078\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23211\
        );

    \I__4077\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23208\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__23226\,
            I => \N__23205\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__23221\,
            I => \N__23200\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__23216\,
            I => \N__23200\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23195\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__23208\,
            I => \N__23195\
        );

    \I__4071\ : Span4Mux_v
    port map (
            O => \N__23205\,
            I => \N__23192\
        );

    \I__4070\ : Span4Mux_h
    port map (
            O => \N__23200\,
            I => \N__23187\
        );

    \I__4069\ : Span4Mux_v
    port map (
            O => \N__23195\,
            I => \N__23187\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__23192\,
            I => \b2v_inst11.N_140_N\
        );

    \I__4067\ : Odrv4
    port map (
            O => \N__23187\,
            I => \b2v_inst11.N_140_N\
        );

    \I__4066\ : InMux
    port map (
            O => \N__23182\,
            I => \N__23176\
        );

    \I__4065\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23168\
        );

    \I__4064\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23168\
        );

    \I__4063\ : CascadeMux
    port map (
            O => \N__23179\,
            I => \N__23161\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23158\
        );

    \I__4061\ : InMux
    port map (
            O => \N__23175\,
            I => \N__23154\
        );

    \I__4060\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23149\
        );

    \I__4059\ : InMux
    port map (
            O => \N__23173\,
            I => \N__23149\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23146\
        );

    \I__4057\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23143\
        );

    \I__4056\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23136\
        );

    \I__4055\ : InMux
    port map (
            O => \N__23165\,
            I => \N__23136\
        );

    \I__4054\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23136\
        );

    \I__4053\ : InMux
    port map (
            O => \N__23161\,
            I => \N__23133\
        );

    \I__4052\ : Span4Mux_v
    port map (
            O => \N__23158\,
            I => \N__23129\
        );

    \I__4051\ : InMux
    port map (
            O => \N__23157\,
            I => \N__23126\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__23154\,
            I => \N__23116\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__23149\,
            I => \N__23116\
        );

    \I__4048\ : Span4Mux_v
    port map (
            O => \N__23146\,
            I => \N__23116\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__23143\,
            I => \N__23116\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__23136\,
            I => \N__23113\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__23133\,
            I => \N__23110\
        );

    \I__4044\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23107\
        );

    \I__4043\ : Span4Mux_h
    port map (
            O => \N__23129\,
            I => \N__23102\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__23102\
        );

    \I__4041\ : InMux
    port map (
            O => \N__23125\,
            I => \N__23099\
        );

    \I__4040\ : Span4Mux_h
    port map (
            O => \N__23116\,
            I => \N__23092\
        );

    \I__4039\ : Span4Mux_s3_h
    port map (
            O => \N__23113\,
            I => \N__23092\
        );

    \I__4038\ : Span4Mux_s3_h
    port map (
            O => \N__23110\,
            I => \N__23092\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__23107\,
            I => \b2v_inst11.N_425\
        );

    \I__4036\ : Odrv4
    port map (
            O => \N__23102\,
            I => \b2v_inst11.N_425\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__23099\,
            I => \b2v_inst11.N_425\
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__23092\,
            I => \b2v_inst11.N_425\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__23083\,
            I => \b2v_inst11.N_154_N_cascade_\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__23080\,
            I => \b2v_inst11.dutycycle_en_4_cascade_\
        );

    \I__4031\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23071\
        );

    \I__4030\ : InMux
    port map (
            O => \N__23076\,
            I => \N__23071\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__23071\,
            I => \b2v_inst11.dutycycle_e_1_8\
        );

    \I__4028\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23062\
        );

    \I__4027\ : InMux
    port map (
            O => \N__23067\,
            I => \N__23048\
        );

    \I__4026\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23038\
        );

    \I__4025\ : InMux
    port map (
            O => \N__23065\,
            I => \N__23038\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__23062\,
            I => \N__23035\
        );

    \I__4023\ : InMux
    port map (
            O => \N__23061\,
            I => \N__23032\
        );

    \I__4022\ : InMux
    port map (
            O => \N__23060\,
            I => \N__23027\
        );

    \I__4021\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23027\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__23058\,
            I => \N__23022\
        );

    \I__4019\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23019\
        );

    \I__4018\ : InMux
    port map (
            O => \N__23056\,
            I => \N__23012\
        );

    \I__4017\ : InMux
    port map (
            O => \N__23055\,
            I => \N__23012\
        );

    \I__4016\ : InMux
    port map (
            O => \N__23054\,
            I => \N__23012\
        );

    \I__4015\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23005\
        );

    \I__4014\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23005\
        );

    \I__4013\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23005\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__23048\,
            I => \N__23002\
        );

    \I__4011\ : InMux
    port map (
            O => \N__23047\,
            I => \N__22997\
        );

    \I__4010\ : InMux
    port map (
            O => \N__23046\,
            I => \N__22997\
        );

    \I__4009\ : InMux
    port map (
            O => \N__23045\,
            I => \N__22992\
        );

    \I__4008\ : InMux
    port map (
            O => \N__23044\,
            I => \N__22992\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__23043\,
            I => \N__22988\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__22983\
        );

    \I__4005\ : Span4Mux_s3_h
    port map (
            O => \N__23035\,
            I => \N__22976\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__23032\,
            I => \N__22976\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__23027\,
            I => \N__22976\
        );

    \I__4002\ : InMux
    port map (
            O => \N__23026\,
            I => \N__22971\
        );

    \I__4001\ : InMux
    port map (
            O => \N__23025\,
            I => \N__22971\
        );

    \I__4000\ : InMux
    port map (
            O => \N__23022\,
            I => \N__22968\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__23019\,
            I => \N__22961\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__23012\,
            I => \N__22961\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__23005\,
            I => \N__22961\
        );

    \I__3996\ : Span4Mux_h
    port map (
            O => \N__23002\,
            I => \N__22954\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__22997\,
            I => \N__22954\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__22992\,
            I => \N__22954\
        );

    \I__3993\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22947\
        );

    \I__3992\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22947\
        );

    \I__3991\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22947\
        );

    \I__3990\ : InMux
    port map (
            O => \N__22986\,
            I => \N__22944\
        );

    \I__3989\ : Span4Mux_v
    port map (
            O => \N__22983\,
            I => \N__22937\
        );

    \I__3988\ : Span4Mux_v
    port map (
            O => \N__22976\,
            I => \N__22937\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__22971\,
            I => \N__22937\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__22968\,
            I => \N__22930\
        );

    \I__3985\ : Span4Mux_h
    port map (
            O => \N__22961\,
            I => \N__22930\
        );

    \I__3984\ : Span4Mux_v
    port map (
            O => \N__22954\,
            I => \N__22930\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__22947\,
            I => \N__22925\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__22944\,
            I => \N__22925\
        );

    \I__3981\ : Span4Mux_h
    port map (
            O => \N__22937\,
            I => \N__22922\
        );

    \I__3980\ : Odrv4
    port map (
            O => \N__22930\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__3979\ : Odrv12
    port map (
            O => \N__22925\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__22922\,
            I => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\
        );

    \I__3977\ : InMux
    port map (
            O => \N__22915\,
            I => \N__22912\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__22912\,
            I => \b2v_inst11.dutycycle_en_4\
        );

    \I__3975\ : InMux
    port map (
            O => \N__22909\,
            I => \N__22903\
        );

    \I__3974\ : InMux
    port map (
            O => \N__22908\,
            I => \N__22903\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__22903\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22893\
        );

    \I__3970\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22890\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__22893\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__22890\,
            I => \b2v_inst11.dutycycleZ0Z_10\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__22885\,
            I => \N__22882\
        );

    \I__3966\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22873\
        );

    \I__3965\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22873\
        );

    \I__3964\ : InMux
    port map (
            O => \N__22880\,
            I => \N__22873\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__22873\,
            I => \b2v_inst11.dutycycleZ1Z_8\
        );

    \I__3962\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22867\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__22867\,
            I => \N__22864\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__22864\,
            I => \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__22861\,
            I => \N__22858\
        );

    \I__3958\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22852\
        );

    \I__3957\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22852\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__22852\,
            I => \b2v_inst11.dutycycle_RNI1KT13Z0Z_8\
        );

    \I__3955\ : InMux
    port map (
            O => \N__22849\,
            I => \N__22846\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__22846\,
            I => \b2v_inst11.dutycycle_RNI_1Z0Z_3\
        );

    \I__3953\ : CascadeMux
    port map (
            O => \N__22843\,
            I => \b2v_inst11.dutycycleZ0Z_8_cascade_\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__22840\,
            I => \b2v_inst11.N_153_N_cascade_\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__22837\,
            I => \b2v_inst11.N_156_N_cascade_\
        );

    \I__3950\ : InMux
    port map (
            O => \N__22834\,
            I => \N__22831\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__22831\,
            I => \b2v_inst11.dutycycle_e_1_9\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__22828\,
            I => \N__22825\
        );

    \I__3947\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22821\
        );

    \I__3946\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22818\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__22821\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__22818\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__22813\,
            I => \b2v_inst11.dutycycle_e_1_9_cascade_\
        );

    \I__3942\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22804\
        );

    \I__3941\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22804\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__22804\,
            I => \b2v_inst11.dutycycleZ1Z_9\
        );

    \I__3939\ : CascadeMux
    port map (
            O => \N__22801\,
            I => \N__22798\
        );

    \I__3938\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22792\
        );

    \I__3937\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22792\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__22792\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\
        );

    \I__3935\ : InMux
    port map (
            O => \N__22789\,
            I => \N__22783\
        );

    \I__3934\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22783\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__22783\,
            I => \b2v_inst11.dutycycle_en_10\
        );

    \I__3932\ : InMux
    port map (
            O => \N__22780\,
            I => \N__22777\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__22777\,
            I => \b2v_inst5.count_rst_10\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__22774\,
            I => \b2v_inst5.countZ0Z_8_cascade_\
        );

    \I__3929\ : InMux
    port map (
            O => \N__22771\,
            I => \N__22765\
        );

    \I__3928\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22765\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__22765\,
            I => \b2v_inst5.count_1_4\
        );

    \I__3926\ : CascadeMux
    port map (
            O => \N__22762\,
            I => \b2v_inst5.un12_clk_100khz_7_cascade_\
        );

    \I__3925\ : CascadeMux
    port map (
            O => \N__22759\,
            I => \b2v_inst11.N_8_1_cascade_\
        );

    \I__3924\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22753\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__22753\,
            I => \N__22750\
        );

    \I__3922\ : Span4Mux_v
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__22747\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_8\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__22744\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_\
        );

    \I__3919\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22738\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__22738\,
            I => \N__22734\
        );

    \I__3917\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22731\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__22734\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__22731\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\
        );

    \I__3914\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__22723\,
            I => \N__22720\
        );

    \I__3912\ : Odrv4
    port map (
            O => \N__22720\,
            I => \b2v_inst11.dutycycle_en_11\
        );

    \I__3911\ : CascadeMux
    port map (
            O => \N__22717\,
            I => \N__22714\
        );

    \I__3910\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22711\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22707\
        );

    \I__3908\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22704\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__22707\,
            I => \N__22701\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__22704\,
            I => \b2v_inst11.dutycycleZ0Z_14\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__22701\,
            I => \b2v_inst11.dutycycleZ0Z_14\
        );

    \I__3904\ : CascadeMux
    port map (
            O => \N__22696\,
            I => \b2v_inst11.dutycycleZ0Z_12_cascade_\
        );

    \I__3903\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22690\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__22690\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_11\
        );

    \I__3901\ : InMux
    port map (
            O => \N__22687\,
            I => \N__22683\
        );

    \I__3900\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22680\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22677\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__22680\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_9\
        );

    \I__3897\ : Odrv4
    port map (
            O => \N__22677\,
            I => \b2v_inst11.dutycycle_RNI_4Z0Z_9\
        );

    \I__3896\ : InMux
    port map (
            O => \N__22672\,
            I => \N__22668\
        );

    \I__3895\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22665\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__22668\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__22665\,
            I => \b2v_inst11.mult1_un124_sum_cry_3_s\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__22660\,
            I => \N__22657\
        );

    \I__3891\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22654\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__22654\,
            I => \N__22651\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__22651\,
            I => \b2v_inst11.mult1_un131_sum_axb_4_l_fx\
        );

    \I__3888\ : InMux
    port map (
            O => \N__22648\,
            I => \N__22645\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__22645\,
            I => \b2v_inst11.g0_13_1\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__22642\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_9_cascade_\
        );

    \I__3885\ : InMux
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__22636\,
            I => \N__22633\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__22633\,
            I => \N__22630\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__22630\,
            I => \b2v_inst200.count_RNIC03N_6Z0Z_0\
        );

    \I__3881\ : InMux
    port map (
            O => \N__22627\,
            I => \N__22624\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22620\
        );

    \I__3879\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22617\
        );

    \I__3878\ : Span4Mux_v
    port map (
            O => \N__22620\,
            I => \N__22614\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__22617\,
            I => \N__22611\
        );

    \I__3876\ : Span4Mux_v
    port map (
            O => \N__22614\,
            I => \N__22608\
        );

    \I__3875\ : Span12Mux_s5_h
    port map (
            O => \N__22611\,
            I => \N__22605\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__22608\,
            I => \N_411\
        );

    \I__3873\ : Odrv12
    port map (
            O => \N__22605\,
            I => \N_411\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__3871\ : InMux
    port map (
            O => \N__22597\,
            I => \N__22590\
        );

    \I__3870\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22590\
        );

    \I__3869\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22587\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22582\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__22587\,
            I => \N__22582\
        );

    \I__3866\ : Span4Mux_h
    port map (
            O => \N__22582\,
            I => \N__22579\
        );

    \I__3865\ : Span4Mux_v
    port map (
            O => \N__22579\,
            I => \N__22576\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__22576\,
            I => \N__22573\
        );

    \I__3863\ : Odrv4
    port map (
            O => \N__22573\,
            I => \b2v_inst200.m11_0_a3_0\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \b2v_inst5.count_rst_10_cascade_\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__22567\,
            I => \b2v_inst5.un2_count_1_axb_4_cascade_\
        );

    \I__3860\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22561\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__22561\,
            I => \b2v_inst5.count_1_8\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__22558\,
            I => \N__22555\
        );

    \I__3857\ : InMux
    port map (
            O => \N__22555\,
            I => \N__22552\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__22552\,
            I => \b2v_inst11.mult1_un124_sum_cry_4_s\
        );

    \I__3855\ : InMux
    port map (
            O => \N__22549\,
            I => \b2v_inst11.mult1_un124_sum_cry_3\
        );

    \I__3854\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22543\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__22543\,
            I => \b2v_inst11.mult1_un124_sum_cry_5_s\
        );

    \I__3852\ : InMux
    port map (
            O => \N__22540\,
            I => \b2v_inst11.mult1_un124_sum_cry_4\
        );

    \I__3851\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22531\
        );

    \I__3850\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22531\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__22531\,
            I => \b2v_inst11.mult1_un124_sum_cry_6_s\
        );

    \I__3848\ : InMux
    port map (
            O => \N__22528\,
            I => \b2v_inst11.mult1_un124_sum_cry_5\
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__3846\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__22519\,
            I => \b2v_inst11.mult1_un131_sum_axb_8\
        );

    \I__3844\ : InMux
    port map (
            O => \N__22516\,
            I => \b2v_inst11.mult1_un124_sum_cry_6\
        );

    \I__3843\ : InMux
    port map (
            O => \N__22513\,
            I => \b2v_inst11.mult1_un124_sum_cry_7\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__22510\,
            I => \b2v_inst11.mult1_un124_sum_s_8_cascade_\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__22507\,
            I => \N__22504\
        );

    \I__3840\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22501\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__22501\,
            I => \b2v_inst11.mult1_un124_sum_i_0_8\
        );

    \I__3838\ : InMux
    port map (
            O => \N__22498\,
            I => \N__22493\
        );

    \I__3837\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22490\
        );

    \I__3836\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22487\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__22493\,
            I => \N__22484\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__22490\,
            I => \N__22480\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__22487\,
            I => \N__22477\
        );

    \I__3832\ : Sp12to4
    port map (
            O => \N__22484\,
            I => \N__22474\
        );

    \I__3831\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22471\
        );

    \I__3830\ : Span4Mux_h
    port map (
            O => \N__22480\,
            I => \N__22468\
        );

    \I__3829\ : Span4Mux_h
    port map (
            O => \N__22477\,
            I => \N__22465\
        );

    \I__3828\ : Odrv12
    port map (
            O => \N__22474\,
            I => \b2v_inst11.N_382\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__22471\,
            I => \b2v_inst11.N_382\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__22468\,
            I => \b2v_inst11.N_382\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__22465\,
            I => \b2v_inst11.N_382\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__3823\ : InMux
    port map (
            O => \N__22453\,
            I => \N__22450\
        );

    \I__3822\ : LocalMux
    port map (
            O => \N__22450\,
            I => \N__22447\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__22447\,
            I => \b2v_inst11.N_302\
        );

    \I__3820\ : InMux
    port map (
            O => \N__22444\,
            I => \b2v_inst11.mult1_un131_sum_cry_2\
        );

    \I__3819\ : InMux
    port map (
            O => \N__22441\,
            I => \b2v_inst11.mult1_un131_sum_cry_3\
        );

    \I__3818\ : InMux
    port map (
            O => \N__22438\,
            I => \b2v_inst11.mult1_un131_sum_cry_4\
        );

    \I__3817\ : InMux
    port map (
            O => \N__22435\,
            I => \b2v_inst11.mult1_un131_sum_cry_5\
        );

    \I__3816\ : InMux
    port map (
            O => \N__22432\,
            I => \b2v_inst11.mult1_un131_sum_cry_6\
        );

    \I__3815\ : InMux
    port map (
            O => \N__22429\,
            I => \b2v_inst11.mult1_un131_sum_cry_7\
        );

    \I__3814\ : CascadeMux
    port map (
            O => \N__22426\,
            I => \N__22423\
        );

    \I__3813\ : InMux
    port map (
            O => \N__22423\,
            I => \N__22420\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__22420\,
            I => \b2v_inst11.mult1_un131_sum_axb_7_l_fx\
        );

    \I__3811\ : InMux
    port map (
            O => \N__22417\,
            I => \b2v_inst11.mult1_un124_sum_cry_2\
        );

    \I__3810\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22411\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__22411\,
            I => \b2v_inst36.DSW_PWROK_0\
        );

    \I__3808\ : InMux
    port map (
            O => \N__22408\,
            I => \N__22405\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__22405\,
            I => \b2v_inst36.curr_state_0_0\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \b2v_inst36.curr_state_7_0_cascade_\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__22399\,
            I => \N__22394\
        );

    \I__3804\ : InMux
    port map (
            O => \N__22398\,
            I => \N__22390\
        );

    \I__3803\ : InMux
    port map (
            O => \N__22397\,
            I => \N__22383\
        );

    \I__3802\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22383\
        );

    \I__3801\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22383\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__22390\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__22383\,
            I => \b2v_inst36.curr_stateZ0Z_0\
        );

    \I__3798\ : CascadeMux
    port map (
            O => \N__22378\,
            I => \b2v_inst36.curr_stateZ0Z_0_cascade_\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__22375\,
            I => \b2v_inst36.N_2939_i_cascade_\
        );

    \I__3796\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22369\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__22369\,
            I => \b2v_inst36.count_2_4\
        );

    \I__3794\ : InMux
    port map (
            O => \N__22366\,
            I => \N__22363\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__22363\,
            I => \b2v_inst36.count_2_9\
        );

    \I__3792\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__22357\,
            I => \b2v_inst36.count_2_12\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__22354\,
            I => \b2v_inst36.curr_state_RNI8TT2Z0Z_0_cascade_\
        );

    \I__3789\ : IoInMux
    port map (
            O => \N__22351\,
            I => \N__22348\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__22348\,
            I => \N__22345\
        );

    \I__3787\ : IoSpan4Mux
    port map (
            O => \N__22345\,
            I => \N__22342\
        );

    \I__3786\ : Span4Mux_s2_h
    port map (
            O => \N__22342\,
            I => \N__22339\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__22339\,
            I => \N__22336\
        );

    \I__3784\ : Odrv4
    port map (
            O => \N__22336\,
            I => \DSW_PWROK_c\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__22333\,
            I => \b2v_inst200.curr_stateZ0Z_1_cascade_\
        );

    \I__3782\ : InMux
    port map (
            O => \N__22330\,
            I => \N__22326\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__22329\,
            I => \N__22319\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22314\
        );

    \I__3779\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22296\
        );

    \I__3778\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22296\
        );

    \I__3777\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22296\
        );

    \I__3776\ : InMux
    port map (
            O => \N__22322\,
            I => \N__22296\
        );

    \I__3775\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22296\
        );

    \I__3774\ : InMux
    port map (
            O => \N__22318\,
            I => \N__22296\
        );

    \I__3773\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22293\
        );

    \I__3772\ : Span12Mux_s7_v
    port map (
            O => \N__22314\,
            I => \N__22290\
        );

    \I__3771\ : InMux
    port map (
            O => \N__22313\,
            I => \N__22287\
        );

    \I__3770\ : InMux
    port map (
            O => \N__22312\,
            I => \N__22278\
        );

    \I__3769\ : InMux
    port map (
            O => \N__22311\,
            I => \N__22278\
        );

    \I__3768\ : InMux
    port map (
            O => \N__22310\,
            I => \N__22278\
        );

    \I__3767\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22278\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22273\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22273\
        );

    \I__3764\ : Odrv12
    port map (
            O => \N__22290\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__22287\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__22278\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__22273\,
            I => \b2v_inst200.count_RNI_0_0\
        );

    \I__3760\ : InMux
    port map (
            O => \N__22264\,
            I => \N__22261\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__22261\,
            I => \N__22258\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__22258\,
            I => \N__22255\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__22255\,
            I => \GPIO_FPGA_SoC_1_c\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__22252\,
            I => \N_411_cascade_\
        );

    \I__3755\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22246\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__22246\,
            I => \b2v_inst200.m6_i_0\
        );

    \I__3753\ : CascadeMux
    port map (
            O => \N__22243\,
            I => \b2v_inst200.m6_i_0_cascade_\
        );

    \I__3752\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22237\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__22237\,
            I => \b2v_inst200.curr_state_3_0\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__22234\,
            I => \b2v_inst200.N_58_cascade_\
        );

    \I__3749\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22220\
        );

    \I__3748\ : InMux
    port map (
            O => \N__22230\,
            I => \N__22220\
        );

    \I__3747\ : InMux
    port map (
            O => \N__22229\,
            I => \N__22220\
        );

    \I__3746\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22215\
        );

    \I__3745\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22215\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__22220\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__22215\,
            I => \b2v_inst200.curr_stateZ0Z_0\
        );

    \I__3742\ : CascadeMux
    port map (
            O => \N__22210\,
            I => \b2v_inst200.curr_stateZ0Z_0_cascade_\
        );

    \I__3741\ : InMux
    port map (
            O => \N__22207\,
            I => \N__22201\
        );

    \I__3740\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22201\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__22201\,
            I => \N_412\
        );

    \I__3738\ : CascadeMux
    port map (
            O => \N__22198\,
            I => \N_412_cascade_\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__22195\,
            I => \N__22187\
        );

    \I__3736\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22181\
        );

    \I__3735\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22181\
        );

    \I__3734\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22176\
        );

    \I__3733\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22176\
        );

    \I__3732\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22169\
        );

    \I__3731\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22169\
        );

    \I__3730\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22169\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__22181\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__22176\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__22169\,
            I => \b2v_inst200.curr_stateZ0Z_1\
        );

    \I__3726\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22159\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__22159\,
            I => \b2v_inst200.curr_state_3_1\
        );

    \I__3724\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22153\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__22153\,
            I => \b2v_inst36.count_2_6\
        );

    \I__3722\ : InMux
    port map (
            O => \N__22150\,
            I => \N__22147\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__22147\,
            I => \b2v_inst11.count_0_9\
        );

    \I__3720\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__22141\,
            I => \b2v_inst11.count_0_10\
        );

    \I__3718\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__22135\,
            I => \b2v_inst11.count_0_11\
        );

    \I__3716\ : InMux
    port map (
            O => \N__22132\,
            I => \N__22129\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__22129\,
            I => \b2v_inst11.count_0_2\
        );

    \I__3714\ : CascadeMux
    port map (
            O => \N__22126\,
            I => \b2v_inst200.N_56_cascade_\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__22123\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1_cascade_\
        );

    \I__3712\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22116\
        );

    \I__3711\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22110\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__22116\,
            I => \N__22107\
        );

    \I__3709\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22104\
        );

    \I__3708\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22099\
        );

    \I__3707\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22099\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__22110\,
            I => \N__22090\
        );

    \I__3705\ : Span4Mux_v
    port map (
            O => \N__22107\,
            I => \N__22087\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__22104\,
            I => \N__22084\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__22099\,
            I => \N__22081\
        );

    \I__3702\ : InMux
    port map (
            O => \N__22098\,
            I => \N__22074\
        );

    \I__3701\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22074\
        );

    \I__3700\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22074\
        );

    \I__3699\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22067\
        );

    \I__3698\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22067\
        );

    \I__3697\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22067\
        );

    \I__3696\ : Span4Mux_s2_v
    port map (
            O => \N__22090\,
            I => \N__22060\
        );

    \I__3695\ : Span4Mux_v
    port map (
            O => \N__22087\,
            I => \N__22060\
        );

    \I__3694\ : Span4Mux_v
    port map (
            O => \N__22084\,
            I => \N__22055\
        );

    \I__3693\ : Span4Mux_h
    port map (
            O => \N__22081\,
            I => \N__22055\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__22050\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22050\
        );

    \I__3690\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22045\
        );

    \I__3689\ : InMux
    port map (
            O => \N__22065\,
            I => \N__22045\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__22060\,
            I => \b2v_inst5_RSMRSTn_latmux\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__22055\,
            I => \b2v_inst5_RSMRSTn_latmux\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__22050\,
            I => \b2v_inst5_RSMRSTn_latmux\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__22045\,
            I => \b2v_inst5_RSMRSTn_latmux\
        );

    \I__3684\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22032\
        );

    \I__3683\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22028\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__22032\,
            I => \N__22025\
        );

    \I__3681\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22022\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22018\
        );

    \I__3679\ : Span4Mux_h
    port map (
            O => \N__22025\,
            I => \N__22013\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__22022\,
            I => \N__22013\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__22021\,
            I => \N__22010\
        );

    \I__3676\ : Span12Mux_s5_h
    port map (
            O => \N__22018\,
            I => \N__22006\
        );

    \I__3675\ : Span4Mux_v
    port map (
            O => \N__22013\,
            I => \N__22003\
        );

    \I__3674\ : InMux
    port map (
            O => \N__22010\,
            I => \N__21998\
        );

    \I__3673\ : InMux
    port map (
            O => \N__22009\,
            I => \N__21998\
        );

    \I__3672\ : Odrv12
    port map (
            O => \N__22006\,
            I => \b2v_inst5_RSMRSTn_fast\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__22003\,
            I => \b2v_inst5_RSMRSTn_fast\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__21998\,
            I => \b2v_inst5_RSMRSTn_fast\
        );

    \I__3669\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21988\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21983\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21987\,
            I => \N__21980\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__21986\,
            I => \N__21974\
        );

    \I__3665\ : Span4Mux_s2_v
    port map (
            O => \N__21983\,
            I => \N__21969\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21969\
        );

    \I__3663\ : InMux
    port map (
            O => \N__21979\,
            I => \N__21966\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21978\,
            I => \N__21959\
        );

    \I__3661\ : InMux
    port map (
            O => \N__21977\,
            I => \N__21959\
        );

    \I__3660\ : InMux
    port map (
            O => \N__21974\,
            I => \N__21959\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__21969\,
            I => \N__21956\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__21966\,
            I => \N__21951\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__21959\,
            I => \N__21951\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__21956\,
            I => \RSMRSTn_0\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__21951\,
            I => \RSMRSTn_0\
        );

    \I__3654\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21939\
        );

    \I__3653\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21939\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21944\,
            I => \N__21936\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__21939\,
            I => \N__21933\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__21936\,
            I => \b2v_inst5.N_2897_i\
        );

    \I__3649\ : Odrv4
    port map (
            O => \N__21933\,
            I => \b2v_inst5.N_2897_i\
        );

    \I__3648\ : InMux
    port map (
            O => \N__21928\,
            I => \N__21915\
        );

    \I__3647\ : InMux
    port map (
            O => \N__21927\,
            I => \N__21915\
        );

    \I__3646\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21915\
        );

    \I__3645\ : InMux
    port map (
            O => \N__21925\,
            I => \N__21915\
        );

    \I__3644\ : InMux
    port map (
            O => \N__21924\,
            I => \N__21912\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21909\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__21912\,
            I => \b2v_inst5.curr_stateZ0Z_0\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__21909\,
            I => \b2v_inst5.curr_stateZ0Z_0\
        );

    \I__3640\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21889\
        );

    \I__3639\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21889\
        );

    \I__3638\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21889\
        );

    \I__3637\ : InMux
    port map (
            O => \N__21901\,
            I => \N__21889\
        );

    \I__3636\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21889\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__21889\,
            I => \b2v_inst5.curr_state_RNIZ0Z_1\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__21886\,
            I => \b2v_inst5.N_51_cascade_\
        );

    \I__3633\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__21880\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_0\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__21877\,
            I => \N__21871\
        );

    \I__3630\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21858\
        );

    \I__3629\ : InMux
    port map (
            O => \N__21875\,
            I => \N__21858\
        );

    \I__3628\ : InMux
    port map (
            O => \N__21874\,
            I => \N__21858\
        );

    \I__3627\ : InMux
    port map (
            O => \N__21871\,
            I => \N__21858\
        );

    \I__3626\ : InMux
    port map (
            O => \N__21870\,
            I => \N__21858\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__21869\,
            I => \N__21854\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__21858\,
            I => \N__21850\
        );

    \I__3623\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21843\
        );

    \I__3622\ : InMux
    port map (
            O => \N__21854\,
            I => \N__21843\
        );

    \I__3621\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21843\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__21850\,
            I => \N__21840\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__21843\,
            I => \N__21837\
        );

    \I__3618\ : Odrv4
    port map (
            O => \N__21840\,
            I => \b2v_inst11.N_19_i\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__21837\,
            I => \b2v_inst11.N_19_i\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__3615\ : InMux
    port map (
            O => \N__21829\,
            I => \N__21826\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__21826\,
            I => \b2v_inst11.N_5572_0\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__3612\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21814\
        );

    \I__3611\ : InMux
    port map (
            O => \N__21819\,
            I => \N__21814\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21809\
        );

    \I__3609\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21806\
        );

    \I__3608\ : InMux
    port map (
            O => \N__21812\,
            I => \N__21803\
        );

    \I__3607\ : Span4Mux_v
    port map (
            O => \N__21809\,
            I => \N__21798\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__21806\,
            I => \N__21798\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__21803\,
            I => \N__21795\
        );

    \I__3604\ : Odrv4
    port map (
            O => \N__21798\,
            I => \b2v_inst11.N_172\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__21795\,
            I => \b2v_inst11.N_172\
        );

    \I__3602\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__21787\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_1\
        );

    \I__3600\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__21781\,
            I => \b2v_inst11.dutycycle_eena\
        );

    \I__3598\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21772\
        );

    \I__3597\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21772\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__21772\,
            I => \b2v_inst11.dutycycleZ1Z_0\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__21769\,
            I => \N__21766\
        );

    \I__3594\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21762\
        );

    \I__3593\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21759\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__21762\,
            I => \b2v_inst11.dutycycle_1_0_0\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__21759\,
            I => \b2v_inst11.dutycycle_1_0_0\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__21754\,
            I => \b2v_inst11.dutycycle_eena_cascade_\
        );

    \I__3589\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21745\
        );

    \I__3588\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21745\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__21745\,
            I => \b2v_inst11.N_117_f0_1\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__21742\,
            I => \b2v_inst11.dutycycle_eena_0_cascade_\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__21739\,
            I => \b2v_inst11.dutycycle_cascade_\
        );

    \I__3584\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21730\
        );

    \I__3583\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21730\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__21730\,
            I => \b2v_inst11.dutycycle_1_0_1\
        );

    \I__3581\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__21724\,
            I => \b2v_inst11.dutycycle_eena_0\
        );

    \I__3579\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21715\
        );

    \I__3578\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21715\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__21715\,
            I => \b2v_inst11.dutycycleZ1Z_1\
        );

    \I__3576\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21706\
        );

    \I__3575\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21706\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__21706\,
            I => \b2v_inst11.dutycycle_0_6\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__3572\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21694\
        );

    \I__3571\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21694\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__21694\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQZ0Z6\
        );

    \I__3569\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21685\
        );

    \I__3568\ : InMux
    port map (
            O => \N__21690\,
            I => \N__21685\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__21679\,
            I => \b2v_inst11.dutycycle_e_1_6\
        );

    \I__3564\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21669\
        );

    \I__3562\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21666\
        );

    \I__3561\ : Span4Mux_v
    port map (
            O => \N__21669\,
            I => \N__21662\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__21666\,
            I => \N__21659\
        );

    \I__3559\ : InMux
    port map (
            O => \N__21665\,
            I => \N__21656\
        );

    \I__3558\ : Span4Mux_h
    port map (
            O => \N__21662\,
            I => \N__21651\
        );

    \I__3557\ : Span4Mux_v
    port map (
            O => \N__21659\,
            I => \N__21651\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__21656\,
            I => \b2v_inst11.func_state_RNI_5Z0Z_1\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__21651\,
            I => \b2v_inst11.func_state_RNI_5Z0Z_1\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__21646\,
            I => \b2v_inst11.N_186_cascade_\
        );

    \I__3553\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__3551\ : Span4Mux_h
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__3550\ : Odrv4
    port map (
            O => \N__21634\,
            I => \b2v_inst11.N_426_0\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__21631\,
            I => \b2v_inst11_g0_i_m2_i_a6_1_1_cascade_\
        );

    \I__3548\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21625\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__21622\,
            I => \N__21619\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__21616\,
            I => \SLP_S3n_ibuf_RNI9HQHZ0Z3\
        );

    \I__3543\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21607\
        );

    \I__3542\ : InMux
    port map (
            O => \N__21612\,
            I => \N__21607\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__3540\ : Span4Mux_v
    port map (
            O => \N__21604\,
            I => \N__21599\
        );

    \I__3539\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21594\
        );

    \I__3538\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21594\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__21599\,
            I => \b2v_inst11.dutycycle_RNI_9Z0Z_1\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__21594\,
            I => \b2v_inst11.dutycycle_RNI_9Z0Z_1\
        );

    \I__3535\ : InMux
    port map (
            O => \N__21589\,
            I => \N__21586\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__21586\,
            I => \b2v_inst11.N_165_0\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__21583\,
            I => \b2v_inst11.g0_i_m2_i_0_1_cascade_\
        );

    \I__3532\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N_15_i_0_a4_1_0\
        );

    \I__3530\ : InMux
    port map (
            O => \N__21574\,
            I => \b2v_inst11.un1_dutycycle_94_cry_12\
        );

    \I__3529\ : InMux
    port map (
            O => \N__21571\,
            I => \b2v_inst11.un1_dutycycle_94_cry_13\
        );

    \I__3528\ : InMux
    port map (
            O => \N__21568\,
            I => \b2v_inst11.un1_dutycycle_94_cry_14\
        );

    \I__3527\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21562\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21559\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__21559\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\
        );

    \I__3524\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21553\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__21553\,
            I => \b2v_inst11.dutycycle_RNIP7P13Z0Z_4\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__21550\,
            I => \N__21546\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__21549\,
            I => \N__21542\
        );

    \I__3520\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21537\
        );

    \I__3519\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21537\
        );

    \I__3518\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21534\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__21537\,
            I => \b2v_inst11.dutycycleZ1Z_4\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__21534\,
            I => \b2v_inst11.dutycycleZ1Z_4\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__21529\,
            I => \b2v_inst11.dutycycle_RNIP7P13Z0Z_4_cascade_\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__21526\,
            I => \b2v_inst11.dutycycleZ0Z_7_cascade_\
        );

    \I__3513\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21517\
        );

    \I__3512\ : InMux
    port map (
            O => \N__21522\,
            I => \N__21517\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__21517\,
            I => \b2v_inst11.dutycycle_e_1_4\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__21514\,
            I => \b2v_inst11.N_158_N_cascade_\
        );

    \I__3509\ : InMux
    port map (
            O => \N__21511\,
            I => \b2v_inst11.un1_dutycycle_94_cry_3\
        );

    \I__3508\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__21502\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19\
        );

    \I__3505\ : InMux
    port map (
            O => \N__21499\,
            I => \b2v_inst11.un1_dutycycle_94_cry_4_cZ0\
        );

    \I__3504\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__3502\ : Span4Mux_h
    port map (
            O => \N__21490\,
            I => \N__21487\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__21487\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29\
        );

    \I__3500\ : InMux
    port map (
            O => \N__21484\,
            I => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__3499\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21478\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__3497\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__21472\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\
        );

    \I__3495\ : InMux
    port map (
            O => \N__21469\,
            I => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__3494\ : InMux
    port map (
            O => \N__21466\,
            I => \bfn_6_10_0_\
        );

    \I__3493\ : InMux
    port map (
            O => \N__21463\,
            I => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\
        );

    \I__3492\ : InMux
    port map (
            O => \N__21460\,
            I => \b2v_inst11.un1_dutycycle_94_cry_9\
        );

    \I__3491\ : InMux
    port map (
            O => \N__21457\,
            I => \N__21451\
        );

    \I__3490\ : InMux
    port map (
            O => \N__21456\,
            I => \N__21451\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__21451\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5\
        );

    \I__3488\ : InMux
    port map (
            O => \N__21448\,
            I => \b2v_inst11.un1_dutycycle_94_cry_10_cZ0\
        );

    \I__3487\ : InMux
    port map (
            O => \N__21445\,
            I => \b2v_inst11.un1_dutycycle_94_cry_11\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__21442\,
            I => \b2v_inst11.un1_dutycycle_53_30_1_0_cascade_\
        );

    \I__3485\ : CascadeMux
    port map (
            O => \N__21439\,
            I => \N__21436\
        );

    \I__3484\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21433\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__21433\,
            I => \b2v_inst11.dutycycle_RNI_2Z0Z_9\
        );

    \I__3482\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21427\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__21427\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_8\
        );

    \I__3480\ : CascadeMux
    port map (
            O => \N__21424\,
            I => \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_\
        );

    \I__3479\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21414\
        );

    \I__3478\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21414\
        );

    \I__3477\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21410\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__21414\,
            I => \N__21407\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__21413\,
            I => \N__21403\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21399\
        );

    \I__3473\ : Span4Mux_v
    port map (
            O => \N__21407\,
            I => \N__21396\
        );

    \I__3472\ : InMux
    port map (
            O => \N__21406\,
            I => \N__21391\
        );

    \I__3471\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21391\
        );

    \I__3470\ : InMux
    port map (
            O => \N__21402\,
            I => \N__21388\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__21399\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_11\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__21396\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_11\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__21391\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_11\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__21388\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_11\
        );

    \I__3465\ : InMux
    port map (
            O => \N__21379\,
            I => \N__21375\
        );

    \I__3464\ : InMux
    port map (
            O => \N__21378\,
            I => \N__21372\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__21375\,
            I => \N__21369\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__21372\,
            I => \N__21366\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__21369\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_1\
        );

    \I__3460\ : Odrv4
    port map (
            O => \N__21366\,
            I => \b2v_inst11.dutycycle_RNI_7Z0Z_1\
        );

    \I__3459\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21358\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__21358\,
            I => \N__21355\
        );

    \I__3457\ : Span4Mux_v
    port map (
            O => \N__21355\,
            I => \N__21352\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__21352\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\
        );

    \I__3455\ : InMux
    port map (
            O => \N__21349\,
            I => \b2v_inst11.un1_dutycycle_94_cry_0\
        );

    \I__3454\ : InMux
    port map (
            O => \N__21346\,
            I => \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__3453\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21340\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__21340\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\
        );

    \I__3451\ : InMux
    port map (
            O => \N__21337\,
            I => \b2v_inst11.un1_dutycycle_94_cry_2\
        );

    \I__3450\ : InMux
    port map (
            O => \N__21334\,
            I => \N__21331\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__21331\,
            I => \b2v_inst11.un2_count_clk_17_0_a2_1_3\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__21328\,
            I => \b2v_inst11.un2_count_clk_17_0_a2_1_2_cascade_\
        );

    \I__3447\ : InMux
    port map (
            O => \N__21325\,
            I => \N__21318\
        );

    \I__3446\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21318\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__21323\,
            I => \N__21315\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__21318\,
            I => \N__21312\
        );

    \I__3443\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21309\
        );

    \I__3442\ : Span4Mux_v
    port map (
            O => \N__21312\,
            I => \N__21304\
        );

    \I__3441\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21304\
        );

    \I__3440\ : Odrv4
    port map (
            O => \N__21304\,
            I => \b2v_inst11.N_363\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__21301\,
            I => \N__21298\
        );

    \I__3438\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21294\
        );

    \I__3437\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21291\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21288\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__21291\,
            I => \b2v_inst11.N_360\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__21288\,
            I => \b2v_inst11.N_360\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__21283\,
            I => \b2v_inst11.N_363_cascade_\
        );

    \I__3432\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21277\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__21277\,
            I => \b2v_inst11.N_365\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__21274\,
            I => \b2v_inst11.N_365_cascade_\
        );

    \I__3429\ : InMux
    port map (
            O => \N__21271\,
            I => \N__21268\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__21268\,
            I => \N__21265\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__21265\,
            I => \b2v_inst11.N_293\
        );

    \I__3426\ : InMux
    port map (
            O => \N__21262\,
            I => \b2v_inst11.mult1_un152_sum_cry_2_c\
        );

    \I__3425\ : InMux
    port map (
            O => \N__21259\,
            I => \b2v_inst11.mult1_un152_sum_cry_3_c\
        );

    \I__3424\ : InMux
    port map (
            O => \N__21256\,
            I => \b2v_inst11.mult1_un152_sum_cry_4_c\
        );

    \I__3423\ : InMux
    port map (
            O => \N__21253\,
            I => \b2v_inst11.mult1_un152_sum_cry_5_c\
        );

    \I__3422\ : InMux
    port map (
            O => \N__21250\,
            I => \b2v_inst11.mult1_un152_sum_cry_6_c\
        );

    \I__3421\ : InMux
    port map (
            O => \N__21247\,
            I => \b2v_inst11.mult1_un152_sum_cry_7\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__21244\,
            I => \N__21239\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__21243\,
            I => \N__21236\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__21242\,
            I => \N__21233\
        );

    \I__3417\ : InMux
    port map (
            O => \N__21239\,
            I => \N__21230\
        );

    \I__3416\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21225\
        );

    \I__3415\ : InMux
    port map (
            O => \N__21233\,
            I => \N__21225\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__21230\,
            I => \b2v_inst11.mult1_un145_sum_i_0_8\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__21225\,
            I => \b2v_inst11.mult1_un145_sum_i_0_8\
        );

    \I__3412\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21217\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__21217\,
            I => \N__21214\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__21214\,
            I => \N__21211\
        );

    \I__3409\ : Span4Mux_v
    port map (
            O => \N__21211\,
            I => \N__21208\
        );

    \I__3408\ : Span4Mux_h
    port map (
            O => \N__21208\,
            I => \N__21205\
        );

    \I__3407\ : Odrv4
    port map (
            O => \N__21205\,
            I => \VDDQ_OK_c\
        );

    \I__3406\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21196\
        );

    \I__3405\ : InMux
    port map (
            O => \N__21201\,
            I => \N__21193\
        );

    \I__3404\ : InMux
    port map (
            O => \N__21200\,
            I => \N__21190\
        );

    \I__3403\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21187\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21184\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__21193\,
            I => \N__21181\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__21190\,
            I => \N__21178\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21174\
        );

    \I__3398\ : Span4Mux_v
    port map (
            O => \N__21184\,
            I => \N__21169\
        );

    \I__3397\ : Span4Mux_v
    port map (
            O => \N__21181\,
            I => \N__21169\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__21178\,
            I => \N__21166\
        );

    \I__3395\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21161\
        );

    \I__3394\ : Span4Mux_v
    port map (
            O => \N__21174\,
            I => \N__21154\
        );

    \I__3393\ : Span4Mux_v
    port map (
            O => \N__21169\,
            I => \N__21154\
        );

    \I__3392\ : Span4Mux_v
    port map (
            O => \N__21166\,
            I => \N__21154\
        );

    \I__3391\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21149\
        );

    \I__3390\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21149\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__21161\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__3388\ : Odrv4
    port map (
            O => \N__21154\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__21149\,
            I => \VCCST_EN_i_0_o3_0\
        );

    \I__3386\ : InMux
    port map (
            O => \N__21142\,
            I => \N__21127\
        );

    \I__3385\ : InMux
    port map (
            O => \N__21141\,
            I => \N__21127\
        );

    \I__3384\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21127\
        );

    \I__3383\ : InMux
    port map (
            O => \N__21139\,
            I => \N__21127\
        );

    \I__3382\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21127\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__21127\,
            I => \N__21124\
        );

    \I__3380\ : Span12Mux_s6_v
    port map (
            O => \N__21124\,
            I => \N__21121\
        );

    \I__3379\ : Odrv12
    port map (
            O => \N__21121\,
            I => \b2v_inst16.N_208_0\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__21118\,
            I => \N__21115\
        );

    \I__3377\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21112\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__21112\,
            I => \N__21109\
        );

    \I__3375\ : Span4Mux_v
    port map (
            O => \N__21109\,
            I => \N__21105\
        );

    \I__3374\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21102\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__21105\,
            I => \b2v_inst11.N_354\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__21102\,
            I => \b2v_inst11.N_354\
        );

    \I__3371\ : InMux
    port map (
            O => \N__21097\,
            I => \N__21091\
        );

    \I__3370\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21091\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__21091\,
            I => \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__21088\,
            I => \N__21085\
        );

    \I__3367\ : InMux
    port map (
            O => \N__21085\,
            I => \N__21082\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__21082\,
            I => \b2v_inst200.count_3_11\
        );

    \I__3365\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21076\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__21076\,
            I => \b2v_inst200.countZ0Z_11\
        );

    \I__3363\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21069\
        );

    \I__3362\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21066\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__21069\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__21066\,
            I => \b2v_inst200.countZ0Z_17\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__21061\,
            I => \b2v_inst200.countZ0Z_11_cascade_\
        );

    \I__3358\ : InMux
    port map (
            O => \N__21058\,
            I => \N__21054\
        );

    \I__3357\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21051\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__21054\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__21051\,
            I => \b2v_inst200.countZ0Z_16\
        );

    \I__3354\ : InMux
    port map (
            O => \N__21046\,
            I => \N__21043\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__21043\,
            I => \N__21040\
        );

    \I__3352\ : Odrv4
    port map (
            O => \N__21040\,
            I => \b2v_inst200.un25_clk_100khz_9\
        );

    \I__3351\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21034\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__21031\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__21031\,
            I => \N__21028\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__21028\,
            I => \b2v_inst200.un25_clk_100khz_12\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__21025\,
            I => \b2v_inst200.un25_clk_100khz_13_cascade_\
        );

    \I__3346\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21019\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__21019\,
            I => \b2v_inst200.un25_clk_100khz_14\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__21016\,
            I => \b2v_inst200.count_RNIC03N_6Z0Z_0_cascade_\
        );

    \I__3343\ : InMux
    port map (
            O => \N__21013\,
            I => \N__21007\
        );

    \I__3342\ : InMux
    port map (
            O => \N__21012\,
            I => \N__21007\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__21007\,
            I => \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0\
        );

    \I__3340\ : InMux
    port map (
            O => \N__21004\,
            I => \N__21001\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__21001\,
            I => \b2v_inst200.count_3_10\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__20998\,
            I => \b2v_inst200.count_RNI_0_0_cascade_\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__20995\,
            I => \N__20991\
        );

    \I__3336\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20988\
        );

    \I__3335\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20985\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__20988\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__20985\,
            I => \b2v_inst200.countZ0Z_10\
        );

    \I__3332\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20977\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__20977\,
            I => \N__20974\
        );

    \I__3330\ : Span4Mux_h
    port map (
            O => \N__20974\,
            I => \N__20970\
        );

    \I__3329\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20967\
        );

    \I__3328\ : Odrv4
    port map (
            O => \N__20970\,
            I => \b2v_inst16.count_rst_1\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__20967\,
            I => \b2v_inst16.count_rst_1\
        );

    \I__3326\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20959\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__20959\,
            I => \N__20956\
        );

    \I__3324\ : Span4Mux_s3_h
    port map (
            O => \N__20956\,
            I => \N__20953\
        );

    \I__3323\ : Odrv4
    port map (
            O => \N__20953\,
            I => \b2v_inst16.count_4_12\
        );

    \I__3322\ : CEMux
    port map (
            O => \N__20950\,
            I => \N__20946\
        );

    \I__3321\ : CEMux
    port map (
            O => \N__20949\,
            I => \N__20929\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20925\
        );

    \I__3319\ : CEMux
    port map (
            O => \N__20945\,
            I => \N__20922\
        );

    \I__3318\ : CEMux
    port map (
            O => \N__20944\,
            I => \N__20919\
        );

    \I__3317\ : CEMux
    port map (
            O => \N__20943\,
            I => \N__20916\
        );

    \I__3316\ : CEMux
    port map (
            O => \N__20942\,
            I => \N__20907\
        );

    \I__3315\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20902\
        );

    \I__3314\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20902\
        );

    \I__3313\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20897\
        );

    \I__3312\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20897\
        );

    \I__3311\ : InMux
    port map (
            O => \N__20937\,
            I => \N__20890\
        );

    \I__3310\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20890\
        );

    \I__3309\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20890\
        );

    \I__3308\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20883\
        );

    \I__3307\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20883\
        );

    \I__3306\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20883\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__20929\,
            I => \N__20879\
        );

    \I__3304\ : CEMux
    port map (
            O => \N__20928\,
            I => \N__20876\
        );

    \I__3303\ : Span4Mux_v
    port map (
            O => \N__20925\,
            I => \N__20873\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20870\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__20919\,
            I => \N__20867\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__20916\,
            I => \N__20864\
        );

    \I__3299\ : InMux
    port map (
            O => \N__20915\,
            I => \N__20859\
        );

    \I__3298\ : CEMux
    port map (
            O => \N__20914\,
            I => \N__20859\
        );

    \I__3297\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20856\
        );

    \I__3296\ : InMux
    port map (
            O => \N__20912\,
            I => \N__20849\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20911\,
            I => \N__20849\
        );

    \I__3294\ : InMux
    port map (
            O => \N__20910\,
            I => \N__20849\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__20907\,
            I => \N__20838\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__20902\,
            I => \N__20838\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__20897\,
            I => \N__20838\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__20890\,
            I => \N__20838\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__20883\,
            I => \N__20838\
        );

    \I__3288\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20835\
        );

    \I__3287\ : Span4Mux_s1_v
    port map (
            O => \N__20879\,
            I => \N__20832\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__20876\,
            I => \N__20829\
        );

    \I__3285\ : Span4Mux_h
    port map (
            O => \N__20873\,
            I => \N__20820\
        );

    \I__3284\ : Span4Mux_v
    port map (
            O => \N__20870\,
            I => \N__20820\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__20867\,
            I => \N__20820\
        );

    \I__3282\ : Span4Mux_s1_h
    port map (
            O => \N__20864\,
            I => \N__20820\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__20859\,
            I => \N__20809\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__20856\,
            I => \N__20809\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__20849\,
            I => \N__20809\
        );

    \I__3278\ : Span4Mux_s1_v
    port map (
            O => \N__20838\,
            I => \N__20809\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20809\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__20832\,
            I => \b2v_inst16.count_en\
        );

    \I__3275\ : Odrv12
    port map (
            O => \N__20829\,
            I => \b2v_inst16.count_en\
        );

    \I__3274\ : Odrv4
    port map (
            O => \N__20820\,
            I => \b2v_inst16.count_en\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__20809\,
            I => \b2v_inst16.count_en\
        );

    \I__3272\ : SRMux
    port map (
            O => \N__20800\,
            I => \N__20793\
        );

    \I__3271\ : SRMux
    port map (
            O => \N__20799\,
            I => \N__20790\
        );

    \I__3270\ : SRMux
    port map (
            O => \N__20798\,
            I => \N__20786\
        );

    \I__3269\ : SRMux
    port map (
            O => \N__20797\,
            I => \N__20782\
        );

    \I__3268\ : SRMux
    port map (
            O => \N__20796\,
            I => \N__20779\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__20793\,
            I => \N__20776\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__20790\,
            I => \N__20773\
        );

    \I__3265\ : SRMux
    port map (
            O => \N__20789\,
            I => \N__20770\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__20786\,
            I => \N__20767\
        );

    \I__3263\ : SRMux
    port map (
            O => \N__20785\,
            I => \N__20764\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__20782\,
            I => \N__20760\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__20779\,
            I => \N__20757\
        );

    \I__3260\ : Span4Mux_h
    port map (
            O => \N__20776\,
            I => \N__20750\
        );

    \I__3259\ : Span4Mux_s3_v
    port map (
            O => \N__20773\,
            I => \N__20750\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__20770\,
            I => \N__20750\
        );

    \I__3257\ : Span4Mux_h
    port map (
            O => \N__20767\,
            I => \N__20745\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20745\
        );

    \I__3255\ : SRMux
    port map (
            O => \N__20763\,
            I => \N__20742\
        );

    \I__3254\ : Span4Mux_s2_v
    port map (
            O => \N__20760\,
            I => \N__20739\
        );

    \I__3253\ : Span4Mux_h
    port map (
            O => \N__20757\,
            I => \N__20736\
        );

    \I__3252\ : Span4Mux_h
    port map (
            O => \N__20750\,
            I => \N__20733\
        );

    \I__3251\ : Span4Mux_v
    port map (
            O => \N__20745\,
            I => \N__20728\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20728\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__20739\,
            I => \N__20725\
        );

    \I__3248\ : Span4Mux_s0_h
    port map (
            O => \N__20736\,
            I => \N__20722\
        );

    \I__3247\ : Span4Mux_s0_h
    port map (
            O => \N__20733\,
            I => \N__20719\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__20728\,
            I => \N__20716\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__20725\,
            I => \b2v_inst16.N_2987_i\
        );

    \I__3244\ : Odrv4
    port map (
            O => \N__20722\,
            I => \b2v_inst16.N_2987_i\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__20719\,
            I => \b2v_inst16.N_2987_i\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__20716\,
            I => \b2v_inst16.N_2987_i\
        );

    \I__3241\ : InMux
    port map (
            O => \N__20707\,
            I => \N__20703\
        );

    \I__3240\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20700\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__20703\,
            I => \N__20688\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__20700\,
            I => \N__20688\
        );

    \I__3237\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20685\
        );

    \I__3236\ : InMux
    port map (
            O => \N__20698\,
            I => \N__20682\
        );

    \I__3235\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20675\
        );

    \I__3234\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20675\
        );

    \I__3233\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20675\
        );

    \I__3232\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20670\
        );

    \I__3231\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20670\
        );

    \I__3230\ : Span4Mux_v
    port map (
            O => \N__20688\,
            I => \N__20659\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__20685\,
            I => \N__20659\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20659\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__20675\,
            I => \N__20659\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__20670\,
            I => \N__20659\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__20659\,
            I => \N__20656\
        );

    \I__3224\ : Odrv4
    port map (
            O => \N__20656\,
            I => \b2v_inst11.N_366\
        );

    \I__3223\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20650\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__20650\,
            I => \N__20647\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__20647\,
            I => \b2v_inst200.count_3_13\
        );

    \I__3220\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20640\
        );

    \I__3219\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20637\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__20640\,
            I => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__20637\,
            I => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\
        );

    \I__3216\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20629\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__20629\,
            I => \b2v_inst200.countZ0Z_13\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__20626\,
            I => \b2v_inst200.countZ0Z_13_cascade_\
        );

    \I__3213\ : InMux
    port map (
            O => \N__20623\,
            I => \N__20619\
        );

    \I__3212\ : InMux
    port map (
            O => \N__20622\,
            I => \N__20616\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__20619\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__20616\,
            I => \b2v_inst200.countZ0Z_0\
        );

    \I__3209\ : InMux
    port map (
            O => \N__20611\,
            I => \N__20607\
        );

    \I__3208\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20604\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20601\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__20604\,
            I => \N__20598\
        );

    \I__3205\ : Span4Mux_h
    port map (
            O => \N__20601\,
            I => \N__20593\
        );

    \I__3204\ : Span4Mux_s1_v
    port map (
            O => \N__20598\,
            I => \N__20593\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__20593\,
            I => \b2v_inst200.countZ0Z_7\
        );

    \I__3202\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20586\
        );

    \I__3201\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20583\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20578\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__20583\,
            I => \N__20578\
        );

    \I__3198\ : Span4Mux_s1_v
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__3197\ : Odrv4
    port map (
            O => \N__20575\,
            I => \b2v_inst200.countZ0Z_5\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__20572\,
            I => \b2v_inst200.un25_clk_100khz_10_cascade_\
        );

    \I__3195\ : InMux
    port map (
            O => \N__20569\,
            I => \N__20566\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__20566\,
            I => \b2v_inst200.un25_clk_100khz_3\
        );

    \I__3193\ : InMux
    port map (
            O => \N__20563\,
            I => \N__20559\
        );

    \I__3192\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20556\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__20559\,
            I => \b2v_inst200.countZ0Z_15\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__20556\,
            I => \b2v_inst200.countZ0Z_15\
        );

    \I__3189\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20545\
        );

    \I__3188\ : InMux
    port map (
            O => \N__20550\,
            I => \N__20545\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__20545\,
            I => \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\
        );

    \I__3186\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20539\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__20539\,
            I => \b2v_inst200.count_3_15\
        );

    \I__3184\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20530\
        );

    \I__3183\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20530\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__20530\,
            I => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\
        );

    \I__3181\ : InMux
    port map (
            O => \N__20527\,
            I => \N__20524\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__20524\,
            I => \b2v_inst200.count_3_14\
        );

    \I__3179\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20517\
        );

    \I__3178\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20514\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__20517\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__20514\,
            I => \b2v_inst200.countZ0Z_14\
        );

    \I__3175\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20506\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20503\
        );

    \I__3173\ : Span4Mux_v
    port map (
            O => \N__20503\,
            I => \N__20500\
        );

    \I__3172\ : Odrv4
    port map (
            O => \N__20500\,
            I => \b2v_inst200.count_0_16\
        );

    \I__3171\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20493\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__20496\,
            I => \N__20490\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__20493\,
            I => \N__20487\
        );

    \I__3168\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20484\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__20487\,
            I => \b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__20484\,
            I => \b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79\
        );

    \I__3165\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__20476\,
            I => \b2v_inst200.countZ0Z_6\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__20473\,
            I => \b2v_inst200.countZ0Z_6_cascade_\
        );

    \I__3162\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20466\
        );

    \I__3161\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20463\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__20466\,
            I => \b2v_inst200.countZ0Z_8\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__20463\,
            I => \b2v_inst200.countZ0Z_8\
        );

    \I__3158\ : InMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__3157\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20452\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__20452\,
            I => \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\
        );

    \I__3155\ : CascadeMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__3154\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__20443\,
            I => \b2v_inst200.count_3_6\
        );

    \I__3152\ : InMux
    port map (
            O => \N__20440\,
            I => \N__20434\
        );

    \I__3151\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20434\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__20434\,
            I => \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0\
        );

    \I__3149\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20428\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__20428\,
            I => \b2v_inst200.count_3_8\
        );

    \I__3147\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20422\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__20422\,
            I => \b2v_inst200.count_1_0\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__20419\,
            I => \b2v_inst200.countZ0Z_0_cascade_\
        );

    \I__3144\ : InMux
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__20413\,
            I => \b2v_inst200.count_3_0\
        );

    \I__3142\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20406\
        );

    \I__3141\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20403\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__20406\,
            I => \N__20400\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20397\
        );

    \I__3138\ : Odrv12
    port map (
            O => \N__20400\,
            I => \b2v_inst200.countZ0Z_12\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__20397\,
            I => \b2v_inst200.countZ0Z_12\
        );

    \I__3136\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__20389\,
            I => \N__20385\
        );

    \I__3134\ : InMux
    port map (
            O => \N__20388\,
            I => \N__20382\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__20385\,
            I => \N__20379\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__20382\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__3131\ : Odrv4
    port map (
            O => \N__20379\,
            I => \b2v_inst20.counterZ0Z_7\
        );

    \I__3130\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__20371\,
            I => \N__20367\
        );

    \I__3128\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20363\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__20367\,
            I => \N__20360\
        );

    \I__3126\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20357\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__20363\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__20360\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__20357\,
            I => \b2v_inst20.counterZ0Z_5\
        );

    \I__3122\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20347\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__20347\,
            I => \N__20343\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__20346\,
            I => \N__20339\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__20343\,
            I => \N__20336\
        );

    \I__3118\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20331\
        );

    \I__3117\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20331\
        );

    \I__3116\ : Odrv4
    port map (
            O => \N__20336\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__20331\,
            I => \b2v_inst20.counterZ0Z_6\
        );

    \I__3114\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20323\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__20323\,
            I => \N__20319\
        );

    \I__3112\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20315\
        );

    \I__3111\ : Span4Mux_s3_h
    port map (
            O => \N__20319\,
            I => \N__20312\
        );

    \I__3110\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20309\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__20315\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__20312\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__20309\,
            I => \b2v_inst20.counterZ0Z_1\
        );

    \I__3106\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20299\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20296\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__20296\,
            I => \b2v_inst20.un4_counter_1_and\
        );

    \I__3103\ : InMux
    port map (
            O => \N__20293\,
            I => \N__20290\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__20290\,
            I => \N__20284\
        );

    \I__3101\ : InMux
    port map (
            O => \N__20289\,
            I => \N__20281\
        );

    \I__3100\ : InMux
    port map (
            O => \N__20288\,
            I => \N__20278\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__20287\,
            I => \N__20273\
        );

    \I__3098\ : Span4Mux_v
    port map (
            O => \N__20284\,
            I => \N__20270\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__20281\,
            I => \N__20267\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20264\
        );

    \I__3095\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20261\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20256\
        );

    \I__3093\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20253\
        );

    \I__3092\ : Span4Mux_h
    port map (
            O => \N__20270\,
            I => \N__20248\
        );

    \I__3091\ : Span4Mux_h
    port map (
            O => \N__20267\,
            I => \N__20248\
        );

    \I__3090\ : Span12Mux_s7_h
    port map (
            O => \N__20264\,
            I => \N__20243\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__20261\,
            I => \N__20243\
        );

    \I__3088\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20236\
        );

    \I__3087\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20236\
        );

    \I__3086\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20236\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__20253\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__3084\ : Odrv4
    port map (
            O => \N__20248\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__3083\ : Odrv12
    port map (
            O => \N__20243\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__20236\,
            I => \SYNTHESIZED_WIRE_1keep_3_fast\
        );

    \I__3081\ : IoInMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__3079\ : Span12Mux_s4_h
    port map (
            O => \N__20221\,
            I => \N__20218\
        );

    \I__3078\ : Odrv12
    port map (
            O => \N__20218\,
            I => \HDA_SDO_ATP_c\
        );

    \I__3077\ : InMux
    port map (
            O => \N__20215\,
            I => \N__20212\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__20212\,
            I => \b2v_inst200.N_205\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__20209\,
            I => \b2v_inst200.N_205_cascade_\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__20206\,
            I => \G_2734_cascade_\
        );

    \I__3073\ : InMux
    port map (
            O => \N__20203\,
            I => \N__20197\
        );

    \I__3072\ : InMux
    port map (
            O => \N__20202\,
            I => \N__20197\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__20197\,
            I => \b2v_inst200.curr_stateZ0Z_2\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__20194\,
            I => \b2v_inst200.curr_stateZ0Z_2_cascade_\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__20191\,
            I => \N__20188\
        );

    \I__3068\ : InMux
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__20185\,
            I => \b2v_inst200.HDA_SDO_ATP_0\
        );

    \I__3066\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20179\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__20179\,
            I => \G_2734\
        );

    \I__3064\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20173\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__20173\,
            I => \b2v_inst200.curr_state_0_2\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__20170\,
            I => \N_73_mux_i_i_a7_4_0_cascade_\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__20167\,
            I => \N__20164\
        );

    \I__3060\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20161\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__20161\,
            I => \b2v_inst11.N_73_mux_i_i_1\
        );

    \I__3058\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20154\
        );

    \I__3057\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20151\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__20154\,
            I => \b2v_inst11.N_73_mux_i_i_2\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__20151\,
            I => \b2v_inst11.N_73_mux_i_i_2\
        );

    \I__3054\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20142\
        );

    \I__3053\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20139\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__20142\,
            I => \N__20134\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20134\
        );

    \I__3050\ : Span4Mux_v
    port map (
            O => \N__20134\,
            I => \N__20131\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__20131\,
            I => \N_15\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__20128\,
            I => \b2v_inst11.N_73_mux_i_i_1_cascade_\
        );

    \I__3047\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20113\
        );

    \I__3046\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20113\
        );

    \I__3045\ : InMux
    port map (
            O => \N__20123\,
            I => \N__20113\
        );

    \I__3044\ : InMux
    port map (
            O => \N__20122\,
            I => \N__20113\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__20113\,
            I => \b2v_inst11.dutycycle_0_5\
        );

    \I__3042\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20107\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__20107\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__20104\,
            I => \RSMRSTn_fast_RNIGMH81_cascade_\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__20101\,
            I => \N__20098\
        );

    \I__3038\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20095\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__20095\,
            I => \N__20091\
        );

    \I__3036\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20088\
        );

    \I__3035\ : Odrv12
    port map (
            O => \N__20091\,
            I => \N_7_2\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N_7_2\
        );

    \I__3033\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20078\
        );

    \I__3032\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20073\
        );

    \I__3031\ : InMux
    port map (
            O => \N__20081\,
            I => \N__20073\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__20078\,
            I => \N__20070\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__20073\,
            I => \N_10_0\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__20070\,
            I => \N_10_0\
        );

    \I__3027\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20062\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__20062\,
            I => \b2v_inst20.tmp_1_rep1_RNI07FZ0Z73\
        );

    \I__3025\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20056\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__20056\,
            I => \N__20053\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__20053\,
            I => \N__20050\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__20050\,
            I => \N__20047\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__20047\,
            I => \b2v_inst20.counter_1_cry_5_THRU_CO\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__20044\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_5_cascade_\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__20041\,
            I => \N__20035\
        );

    \I__3018\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20028\
        );

    \I__3017\ : InMux
    port map (
            O => \N__20039\,
            I => \N__20028\
        );

    \I__3016\ : InMux
    port map (
            O => \N__20038\,
            I => \N__20028\
        );

    \I__3015\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20025\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__20028\,
            I => \N__20022\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__20016\
        );

    \I__3012\ : Span4Mux_h
    port map (
            O => \N__20022\,
            I => \N__20016\
        );

    \I__3011\ : InMux
    port map (
            O => \N__20021\,
            I => \N__20013\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__20016\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_1\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__20013\,
            I => \b2v_inst11.dutycycle_RNI_3Z0Z_1\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__20008\,
            I => \b2v_inst11.N_73_mux_i_i_o7_1_cascade_\
        );

    \I__3007\ : InMux
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__20002\,
            I => \b2v_inst11.dutycycle_RNIUNGA5Z0Z_5\
        );

    \I__3005\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19996\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__19996\,
            I => \b2v_inst11.N_73_mux_i_i_0\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__19993\,
            I => \b2v_inst11.N_73_mux_i_i_a7_1_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19983\
        );

    \I__3001\ : InMux
    port map (
            O => \N__19989\,
            I => \N__19983\
        );

    \I__3000\ : InMux
    port map (
            O => \N__19988\,
            I => \N__19980\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__19983\,
            I => \N__19977\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__19980\,
            I => \N__19972\
        );

    \I__2997\ : Span4Mux_h
    port map (
            O => \N__19977\,
            I => \N__19972\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__19972\,
            I => \N__19969\
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__19969\,
            I => g0_0_0
        );

    \I__2994\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19959\
        );

    \I__2993\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19959\
        );

    \I__2992\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19956\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__19959\,
            I => \N_5_0\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__19956\,
            I => \N_5_0\
        );

    \I__2989\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19944\
        );

    \I__2987\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19941\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__19944\,
            I => \N__19936\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__19941\,
            I => \N__19936\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__19936\,
            I => b2v_inst11_un1_dutycycle_172_m3_amcf1
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__19933\,
            I => \N_73_mux_i_i_a7_4_0_1_cascade_\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__19930\,
            I => \b2v_inst5.N_2897_i_cascade_\
        );

    \I__2981\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19924\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__19924\,
            I => \b2v_inst5.curr_state_0_0\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__19921\,
            I => \b2v_inst5.m4_0_cascade_\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__19918\,
            I => \b2v_inst11.g2_0_1_cascade_\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__19915\,
            I => \dutycycle_RNISSAOS1_0_5_cascade_\
        );

    \I__2976\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__19909\,
            I => \b2v_inst11.N_301\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \b2v_inst11.N_382_cascade_\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__19903\,
            I => \b2v_inst11.g0_2_0_cascade_\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__19900\,
            I => \N__19897\
        );

    \I__2971\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19893\
        );

    \I__2970\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19890\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__19893\,
            I => \N__19885\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__19890\,
            I => \N__19885\
        );

    \I__2967\ : Span4Mux_h
    port map (
            O => \N__19885\,
            I => \N__19882\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__19882\,
            I => \b2v_inst11.N_430\
        );

    \I__2965\ : InMux
    port map (
            O => \N__19879\,
            I => \N__19876\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__19876\,
            I => \b2v_inst11.func_state_RNIRF2E4Z0Z_0\
        );

    \I__2963\ : IoInMux
    port map (
            O => \N__19873\,
            I => \N__19870\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19867\
        );

    \I__2961\ : IoSpan4Mux
    port map (
            O => \N__19867\,
            I => \N__19864\
        );

    \I__2960\ : Span4Mux_s2_h
    port map (
            O => \N__19864\,
            I => \N__19861\
        );

    \I__2959\ : Odrv4
    port map (
            O => \N__19861\,
            I => \VCCST_EN_i_0_i\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__19858\,
            I => \N__19855\
        );

    \I__2957\ : InMux
    port map (
            O => \N__19855\,
            I => \N__19852\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__19852\,
            I => \b2v_inst11.un1_clk_100khz_2_i_o3_sx\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19849\,
            I => \N__19844\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__19848\,
            I => \N__19836\
        );

    \I__2953\ : CascadeMux
    port map (
            O => \N__19847\,
            I => \N__19833\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19830\
        );

    \I__2951\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19827\
        );

    \I__2950\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19822\
        );

    \I__2949\ : InMux
    port map (
            O => \N__19841\,
            I => \N__19822\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__19840\,
            I => \N__19819\
        );

    \I__2947\ : InMux
    port map (
            O => \N__19839\,
            I => \N__19816\
        );

    \I__2946\ : InMux
    port map (
            O => \N__19836\,
            I => \N__19808\
        );

    \I__2945\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19808\
        );

    \I__2944\ : Span4Mux_s2_h
    port map (
            O => \N__19830\,
            I => \N__19803\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__19827\,
            I => \N__19803\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__19822\,
            I => \N__19800\
        );

    \I__2941\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19797\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__19816\,
            I => \N__19794\
        );

    \I__2939\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19787\
        );

    \I__2938\ : InMux
    port map (
            O => \N__19814\,
            I => \N__19787\
        );

    \I__2937\ : InMux
    port map (
            O => \N__19813\,
            I => \N__19787\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__19808\,
            I => \N__19784\
        );

    \I__2935\ : Span4Mux_v
    port map (
            O => \N__19803\,
            I => \N__19781\
        );

    \I__2934\ : Span4Mux_s3_h
    port map (
            O => \N__19800\,
            I => \N__19778\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__19797\,
            I => \N__19775\
        );

    \I__2932\ : Odrv12
    port map (
            O => \N__19794\,
            I => \b2v_inst11.func_state\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__19787\,
            I => \b2v_inst11.func_state\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__19784\,
            I => \b2v_inst11.func_state\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__19781\,
            I => \b2v_inst11.func_state\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__19778\,
            I => \b2v_inst11.func_state\
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__19775\,
            I => \b2v_inst11.func_state\
        );

    \I__2926\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19757\
        );

    \I__2925\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19751\
        );

    \I__2924\ : InMux
    port map (
            O => \N__19760\,
            I => \N__19751\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__19757\,
            I => \N__19748\
        );

    \I__2922\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19745\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__19751\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__19748\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__19745\,
            I => \b2v_inst11.func_state_RNI_0Z0Z_0\
        );

    \I__2918\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19735\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__19735\,
            I => \b2v_inst11.N_305\
        );

    \I__2916\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19723\
        );

    \I__2914\ : InMux
    port map (
            O => \N__19728\,
            I => \N__19720\
        );

    \I__2913\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19715\
        );

    \I__2912\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19715\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__19723\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_6\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__19720\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_6\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__19715\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_6\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__19708\,
            I => \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__19705\,
            I => \b2v_inst11.i2_mux_cascade_\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__19702\,
            I => \b2v_inst11.N_307_cascade_\
        );

    \I__2905\ : InMux
    port map (
            O => \N__19699\,
            I => \N__19696\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__19696\,
            I => \b2v_inst11.N_234_N\
        );

    \I__2903\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19690\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__19690\,
            I => \N__19687\
        );

    \I__2901\ : Odrv4
    port map (
            O => \N__19687\,
            I => \b2v_inst11.N_308\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \b2v_inst11.N_234_N_cascade_\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__19681\,
            I => \b2v_inst11.func_state_RNI9R6T4Z0Z_1_cascade_\
        );

    \I__2898\ : InMux
    port map (
            O => \N__19678\,
            I => \N__19675\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__19675\,
            I => \b2v_inst11.func_state_RNI9R6T4Z0Z_1\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__19672\,
            I => \N__19669\
        );

    \I__2895\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19663\
        );

    \I__2894\ : InMux
    port map (
            O => \N__19668\,
            I => \N__19663\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__19663\,
            I => \b2v_inst11.dutycycleZ1Z_11\
        );

    \I__2892\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19657\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__19657\,
            I => \N__19654\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__19654\,
            I => \b2v_inst11.N_159\
        );

    \I__2889\ : InMux
    port map (
            O => \N__19651\,
            I => \N__19648\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__19648\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__19645\,
            I => \b2v_inst11.N_155_N_cascade_\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__19642\,
            I => \b2v_inst11.dutycycle_en_11_cascade_\
        );

    \I__2885\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19636\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__19636\,
            I => \b2v_inst11.g2_0\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__19633\,
            I => \b2v_inst11.dutycycle_eena_8_cascade_\
        );

    \I__2882\ : InMux
    port map (
            O => \N__19630\,
            I => \N__19627\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__19627\,
            I => \b2v_inst11.dutycycle_rst_7\
        );

    \I__2880\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19618\
        );

    \I__2879\ : InMux
    port map (
            O => \N__19623\,
            I => \N__19618\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__19618\,
            I => \b2v_inst11.dutycycle_0_3\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__19615\,
            I => \b2v_inst11.dutycycle_rst_7_cascade_\
        );

    \I__2876\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19609\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__19609\,
            I => \b2v_inst11.dutycycle_eena_8\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__19606\,
            I => \b2v_inst11.dutycycleZ0Z_3_cascade_\
        );

    \I__2873\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19600\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__19600\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0\
        );

    \I__2871\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19594\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__19594\,
            I => \N__19591\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__19591\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_0_ccf1\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__19588\,
            I => \N__19585\
        );

    \I__2867\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__19582\,
            I => \b2v_inst11.un1_clk_100khz_43_and_i_0_c\
        );

    \I__2865\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19573\
        );

    \I__2864\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19573\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__19573\,
            I => \N__19570\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__19570\,
            I => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\
        );

    \I__2861\ : InMux
    port map (
            O => \N__19567\,
            I => \N__19564\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__19564\,
            I => \N__19560\
        );

    \I__2859\ : InMux
    port map (
            O => \N__19563\,
            I => \N__19557\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__19560\,
            I => \N__19554\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__19557\,
            I => \b2v_inst11.count_off_1_6\
        );

    \I__2856\ : Odrv4
    port map (
            O => \N__19554\,
            I => \b2v_inst11.count_off_1_6\
        );

    \I__2855\ : InMux
    port map (
            O => \N__19549\,
            I => \N__19543\
        );

    \I__2854\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19543\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__19543\,
            I => \N__19540\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__19540\,
            I => \b2v_inst11.count_offZ0Z_7\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__19537\,
            I => \N__19527\
        );

    \I__2850\ : CEMux
    port map (
            O => \N__19536\,
            I => \N__19522\
        );

    \I__2849\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19510\
        );

    \I__2848\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19510\
        );

    \I__2847\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19503\
        );

    \I__2846\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19503\
        );

    \I__2845\ : InMux
    port map (
            O => \N__19531\,
            I => \N__19503\
        );

    \I__2844\ : InMux
    port map (
            O => \N__19530\,
            I => \N__19496\
        );

    \I__2843\ : InMux
    port map (
            O => \N__19527\,
            I => \N__19496\
        );

    \I__2842\ : CEMux
    port map (
            O => \N__19526\,
            I => \N__19496\
        );

    \I__2841\ : CEMux
    port map (
            O => \N__19525\,
            I => \N__19491\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__19522\,
            I => \N__19481\
        );

    \I__2839\ : CEMux
    port map (
            O => \N__19521\,
            I => \N__19476\
        );

    \I__2838\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19476\
        );

    \I__2837\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19465\
        );

    \I__2836\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19465\
        );

    \I__2835\ : CEMux
    port map (
            O => \N__19517\,
            I => \N__19465\
        );

    \I__2834\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19465\
        );

    \I__2833\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19465\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__19510\,
            I => \N__19462\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__19503\,
            I => \N__19459\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19455\
        );

    \I__2829\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19450\
        );

    \I__2828\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19450\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19447\
        );

    \I__2826\ : InMux
    port map (
            O => \N__19490\,
            I => \N__19438\
        );

    \I__2825\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19438\
        );

    \I__2824\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19438\
        );

    \I__2823\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19438\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__19486\,
            I => \N__19435\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__19485\,
            I => \N__19432\
        );

    \I__2820\ : CEMux
    port map (
            O => \N__19484\,
            I => \N__19428\
        );

    \I__2819\ : Span4Mux_s3_v
    port map (
            O => \N__19481\,
            I => \N__19421\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__19476\,
            I => \N__19421\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__19465\,
            I => \N__19421\
        );

    \I__2816\ : Span4Mux_h
    port map (
            O => \N__19462\,
            I => \N__19416\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__19459\,
            I => \N__19416\
        );

    \I__2814\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19413\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__19455\,
            I => \N__19410\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__19450\,
            I => \N__19407\
        );

    \I__2811\ : Span4Mux_s3_v
    port map (
            O => \N__19447\,
            I => \N__19402\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__19438\,
            I => \N__19402\
        );

    \I__2809\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19395\
        );

    \I__2808\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19395\
        );

    \I__2807\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19395\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__19428\,
            I => \N__19392\
        );

    \I__2805\ : Span4Mux_v
    port map (
            O => \N__19421\,
            I => \N__19389\
        );

    \I__2804\ : Span4Mux_v
    port map (
            O => \N__19416\,
            I => \N__19384\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__19413\,
            I => \N__19384\
        );

    \I__2802\ : Span4Mux_h
    port map (
            O => \N__19410\,
            I => \N__19379\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__19407\,
            I => \N__19379\
        );

    \I__2800\ : Span4Mux_h
    port map (
            O => \N__19402\,
            I => \N__19374\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__19395\,
            I => \N__19374\
        );

    \I__2798\ : Odrv12
    port map (
            O => \N__19392\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__19389\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2796\ : Odrv4
    port map (
            O => \N__19384\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2795\ : Odrv4
    port map (
            O => \N__19379\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__19374\,
            I => \b2v_inst11.count_off_enZ0\
        );

    \I__2793\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19357\
        );

    \I__2792\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19357\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__19354\,
            I => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__19351\,
            I => \N__19344\
        );

    \I__2788\ : InMux
    port map (
            O => \N__19350\,
            I => \N__19310\
        );

    \I__2787\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19310\
        );

    \I__2786\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19310\
        );

    \I__2785\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19305\
        );

    \I__2784\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19305\
        );

    \I__2783\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19302\
        );

    \I__2782\ : InMux
    port map (
            O => \N__19342\,
            I => \N__19293\
        );

    \I__2781\ : InMux
    port map (
            O => \N__19341\,
            I => \N__19293\
        );

    \I__2780\ : InMux
    port map (
            O => \N__19340\,
            I => \N__19293\
        );

    \I__2779\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19293\
        );

    \I__2778\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19286\
        );

    \I__2777\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19286\
        );

    \I__2776\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19286\
        );

    \I__2775\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19273\
        );

    \I__2774\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19273\
        );

    \I__2773\ : InMux
    port map (
            O => \N__19333\,
            I => \N__19273\
        );

    \I__2772\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19273\
        );

    \I__2771\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19273\
        );

    \I__2770\ : InMux
    port map (
            O => \N__19330\,
            I => \N__19273\
        );

    \I__2769\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19260\
        );

    \I__2768\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19260\
        );

    \I__2767\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19260\
        );

    \I__2766\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19260\
        );

    \I__2765\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19260\
        );

    \I__2764\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19260\
        );

    \I__2763\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19245\
        );

    \I__2762\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19245\
        );

    \I__2761\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19245\
        );

    \I__2760\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19245\
        );

    \I__2759\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19245\
        );

    \I__2758\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19245\
        );

    \I__2757\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19245\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__19310\,
            I => \N__19240\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__19305\,
            I => \N__19240\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__19302\,
            I => \N__19229\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__19293\,
            I => \N__19229\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__19286\,
            I => \N__19229\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__19273\,
            I => \N__19229\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__19260\,
            I => \N__19229\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__19245\,
            I => \N__19224\
        );

    \I__2748\ : Span4Mux_h
    port map (
            O => \N__19240\,
            I => \N__19224\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__19229\,
            I => \N__19221\
        );

    \I__2746\ : Odrv4
    port map (
            O => \N__19224\,
            I => \b2v_inst11.N_125\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__19221\,
            I => \b2v_inst11.N_125\
        );

    \I__2744\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19212\
        );

    \I__2743\ : InMux
    port map (
            O => \N__19215\,
            I => \N__19209\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__19212\,
            I => \N__19206\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__19209\,
            I => \N__19203\
        );

    \I__2740\ : Span4Mux_s2_v
    port map (
            O => \N__19206\,
            I => \N__19198\
        );

    \I__2739\ : Span4Mux_s2_v
    port map (
            O => \N__19203\,
            I => \N__19198\
        );

    \I__2738\ : Odrv4
    port map (
            O => \N__19198\,
            I => \b2v_inst11.count_off_1_7\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__19195\,
            I => \N__19192\
        );

    \I__2736\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__19189\,
            I => \b2v_inst11.g0_3_0\
        );

    \I__2734\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19182\
        );

    \I__2733\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19179\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__19182\,
            I => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__19179\,
            I => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\
        );

    \I__2730\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19168\
        );

    \I__2729\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19168\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__19168\,
            I => \b2v_inst11.count_offZ0Z_2\
        );

    \I__2727\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19161\
        );

    \I__2726\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19158\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__19161\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__19158\,
            I => \b2v_inst11.count_offZ0Z_5\
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__19153\,
            I => \N__19150\
        );

    \I__2722\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19146\
        );

    \I__2721\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19142\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__19146\,
            I => \N__19139\
        );

    \I__2719\ : InMux
    port map (
            O => \N__19145\,
            I => \N__19136\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19133\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__19139\,
            I => \N__19126\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__19136\,
            I => \N__19126\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__19133\,
            I => \N__19126\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__19126\,
            I => \b2v_inst11.count_offZ0Z_1\
        );

    \I__2713\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19120\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__19120\,
            I => \b2v_inst11.un34_clk_100khz_0\
        );

    \I__2711\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19114\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__19114\,
            I => \b2v_inst11.un34_clk_100khz_2\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__19111\,
            I => \b2v_inst11.un34_clk_100khz_1_cascade_\
        );

    \I__2708\ : InMux
    port map (
            O => \N__19108\,
            I => \N__19105\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19102\
        );

    \I__2706\ : Odrv4
    port map (
            O => \N__19102\,
            I => \b2v_inst11.un34_clk_100khz_3\
        );

    \I__2705\ : InMux
    port map (
            O => \N__19099\,
            I => \N__19096\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__19096\,
            I => \b2v_inst11.un34_clk_100khz_12\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__19093\,
            I => \N__19089\
        );

    \I__2702\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19084\
        );

    \I__2701\ : InMux
    port map (
            O => \N__19089\,
            I => \N__19084\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__19084\,
            I => \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__19081\,
            I => \N__19078\
        );

    \I__2698\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19075\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__19075\,
            I => \b2v_inst11.count_off_0_5\
        );

    \I__2696\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19069\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__19069\,
            I => \N__19066\
        );

    \I__2694\ : Span4Mux_s2_h
    port map (
            O => \N__19066\,
            I => \N__19062\
        );

    \I__2693\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19059\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__19062\,
            I => \N__19056\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__19059\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__2690\ : Odrv4
    port map (
            O => \N__19056\,
            I => \b2v_inst11.count_offZ0Z_6\
        );

    \I__2689\ : InMux
    port map (
            O => \N__19051\,
            I => \N__19045\
        );

    \I__2688\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19045\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__19045\,
            I => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\
        );

    \I__2686\ : InMux
    port map (
            O => \N__19042\,
            I => \N__19039\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__19039\,
            I => \b2v_inst11.count_off_1_9\
        );

    \I__2684\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19032\
        );

    \I__2683\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19029\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__19032\,
            I => \b2v_inst11.count_offZ0Z_9\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__19029\,
            I => \b2v_inst11.count_offZ0Z_9\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__19024\,
            I => \b2v_inst11.count_off_1_9_cascade_\
        );

    \I__2679\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19018\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__19018\,
            I => \b2v_inst11.un3_count_off_1_axb_9\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__19015\,
            I => \b2v_inst11.count_off_1_3_cascade_\
        );

    \I__2676\ : InMux
    port map (
            O => \N__19012\,
            I => \N__19009\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__19009\,
            I => \b2v_inst11.un3_count_off_1_axb_3\
        );

    \I__2674\ : InMux
    port map (
            O => \N__19006\,
            I => \N__19003\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__19003\,
            I => \b2v_inst11.count_offZ0Z_4\
        );

    \I__2672\ : InMux
    port map (
            O => \N__19000\,
            I => \N__18997\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__18997\,
            I => \b2v_inst11.count_off_1_3\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__18994\,
            I => \b2v_inst11.count_offZ0Z_4_cascade_\
        );

    \I__2669\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18985\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18985\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__18985\,
            I => \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18976\
        );

    \I__2665\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18976\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__18976\,
            I => \b2v_inst11.count_offZ0Z_3\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__18973\,
            I => \N__18970\
        );

    \I__2662\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18964\
        );

    \I__2661\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18964\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__18964\,
            I => \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__18961\,
            I => \N__18958\
        );

    \I__2658\ : InMux
    port map (
            O => \N__18958\,
            I => \N__18955\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__18955\,
            I => \b2v_inst11.count_off_0_4\
        );

    \I__2656\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18949\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__18949\,
            I => \b2v_inst11.count_off_0_14\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__18946\,
            I => \N__18943\
        );

    \I__2653\ : InMux
    port map (
            O => \N__18943\,
            I => \N__18937\
        );

    \I__2652\ : InMux
    port map (
            O => \N__18942\,
            I => \N__18937\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__18937\,
            I => \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\
        );

    \I__2650\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18930\
        );

    \I__2649\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18927\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__18930\,
            I => \b2v_inst11.count_offZ0Z_14\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__18927\,
            I => \b2v_inst11.count_offZ0Z_14\
        );

    \I__2646\ : InMux
    port map (
            O => \N__18922\,
            I => \N__18916\
        );

    \I__2645\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18916\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__18916\,
            I => \b2v_inst11.count_off_1_2\
        );

    \I__2643\ : InMux
    port map (
            O => \N__18913\,
            I => \N__18910\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__18910\,
            I => \b2v_inst11.un3_count_off_1_axb_2\
        );

    \I__2641\ : InMux
    port map (
            O => \N__18907\,
            I => \b2v_inst200.un2_count_1_cry_10\
        );

    \I__2640\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18900\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18897\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__18900\,
            I => \N__18894\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__18897\,
            I => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__18894\,
            I => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\
        );

    \I__2635\ : InMux
    port map (
            O => \N__18889\,
            I => \b2v_inst200.un2_count_1_cry_11\
        );

    \I__2634\ : InMux
    port map (
            O => \N__18886\,
            I => \b2v_inst200.un2_count_1_cry_12\
        );

    \I__2633\ : InMux
    port map (
            O => \N__18883\,
            I => \b2v_inst200.un2_count_1_cry_13\
        );

    \I__2632\ : InMux
    port map (
            O => \N__18880\,
            I => \b2v_inst200.un2_count_1_cry_14\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18877\,
            I => \bfn_5_3_0_\
        );

    \I__2630\ : InMux
    port map (
            O => \N__18874\,
            I => \b2v_inst200.un2_count_1_cry_16\
        );

    \I__2629\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18868\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__18868\,
            I => \b2v_inst200.count_0_17\
        );

    \I__2627\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18861\
        );

    \I__2626\ : InMux
    port map (
            O => \N__18864\,
            I => \N__18858\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__18861\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__18858\,
            I => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\
        );

    \I__2623\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18849\
        );

    \I__2622\ : InMux
    port map (
            O => \N__18852\,
            I => \N__18846\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__18849\,
            I => \b2v_inst200.countZ0Z_3\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__18846\,
            I => \b2v_inst200.countZ0Z_3\
        );

    \I__2619\ : InMux
    port map (
            O => \N__18841\,
            I => \N__18835\
        );

    \I__2618\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18835\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__18835\,
            I => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\
        );

    \I__2616\ : InMux
    port map (
            O => \N__18832\,
            I => \b2v_inst200.un2_count_1_cry_2\
        );

    \I__2615\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18825\
        );

    \I__2614\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18822\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__18825\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__18822\,
            I => \b2v_inst200.countZ0Z_4\
        );

    \I__2611\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18813\
        );

    \I__2610\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18810\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__18813\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__18810\,
            I => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\
        );

    \I__2607\ : InMux
    port map (
            O => \N__18805\,
            I => \b2v_inst200.un2_count_1_cry_3\
        );

    \I__2606\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18799\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__18799\,
            I => \N__18795\
        );

    \I__2604\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18792\
        );

    \I__2603\ : Span4Mux_v
    port map (
            O => \N__18795\,
            I => \N__18789\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__18792\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__18789\,
            I => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\
        );

    \I__2600\ : InMux
    port map (
            O => \N__18784\,
            I => \b2v_inst200.un2_count_1_cry_4\
        );

    \I__2599\ : InMux
    port map (
            O => \N__18781\,
            I => \b2v_inst200.un2_count_1_cry_5_cZ0\
        );

    \I__2598\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__18775\,
            I => \N__18771\
        );

    \I__2596\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18768\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__18771\,
            I => \N__18765\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__18768\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__18765\,
            I => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\
        );

    \I__2592\ : InMux
    port map (
            O => \N__18760\,
            I => \b2v_inst200.un2_count_1_cry_6\
        );

    \I__2591\ : InMux
    port map (
            O => \N__18757\,
            I => \bfn_5_2_0_\
        );

    \I__2590\ : InMux
    port map (
            O => \N__18754\,
            I => \b2v_inst200.un2_count_1_cry_8\
        );

    \I__2589\ : InMux
    port map (
            O => \N__18751\,
            I => \b2v_inst200.un2_count_1_cry_9\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__18748\,
            I => \N__18745\
        );

    \I__2587\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18742\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__18742\,
            I => \N__18737\
        );

    \I__2585\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18731\
        );

    \I__2584\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18731\
        );

    \I__2583\ : Span4Mux_s3_h
    port map (
            O => \N__18737\,
            I => \N__18728\
        );

    \I__2582\ : InMux
    port map (
            O => \N__18736\,
            I => \N__18725\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__18731\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__2580\ : Odrv4
    port map (
            O => \N__18728\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__18725\,
            I => \b2v_inst20.counterZ0Z_0\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__18718\,
            I => \N__18714\
        );

    \I__2577\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18709\
        );

    \I__2576\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18709\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__2574\ : Span4Mux_s2_h
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__18703\,
            I => \N__18700\
        );

    \I__2572\ : Span4Mux_v
    port map (
            O => \N__18700\,
            I => \N__18696\
        );

    \I__2571\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18693\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__18696\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__18693\,
            I => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\
        );

    \I__2568\ : InMux
    port map (
            O => \N__18688\,
            I => \N__18685\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__18682\,
            I => \N__18679\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__18679\,
            I => \b2v_inst20.counter_1_cry_3_THRU_CO\
        );

    \I__2564\ : InMux
    port map (
            O => \N__18676\,
            I => \N__18673\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__18673\,
            I => \N__18669\
        );

    \I__2562\ : InMux
    port map (
            O => \N__18672\,
            I => \N__18665\
        );

    \I__2561\ : Span4Mux_v
    port map (
            O => \N__18669\,
            I => \N__18662\
        );

    \I__2560\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18659\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__18665\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__18662\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__18659\,
            I => \b2v_inst20.counterZ0Z_4\
        );

    \I__2556\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18649\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__18649\,
            I => \N__18646\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__18646\,
            I => \N__18643\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__18643\,
            I => \b2v_inst20.counter_1_cry_4_THRU_CO\
        );

    \I__2552\ : IoInMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__18637\,
            I => \N__18632\
        );

    \I__2550\ : IoInMux
    port map (
            O => \N__18636\,
            I => \N__18629\
        );

    \I__2549\ : IoInMux
    port map (
            O => \N__18635\,
            I => \N__18626\
        );

    \I__2548\ : IoSpan4Mux
    port map (
            O => \N__18632\,
            I => \N__18621\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__18629\,
            I => \N__18621\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__18626\,
            I => \N__18618\
        );

    \I__2545\ : IoSpan4Mux
    port map (
            O => \N__18621\,
            I => \N__18615\
        );

    \I__2544\ : Span12Mux_s0_v
    port map (
            O => \N__18618\,
            I => \N__18612\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__18615\,
            I => \delayed_vccin_vccinaux_ok_RNI8L1J7_0\
        );

    \I__2542\ : Odrv12
    port map (
            O => \N__18612\,
            I => \delayed_vccin_vccinaux_ok_RNI8L1J7_0\
        );

    \I__2541\ : InMux
    port map (
            O => \N__18607\,
            I => \N__18604\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__2539\ : Span4Mux_s3_v
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__18598\,
            I => \b2v_inst20.counter_1_cry_1_THRU_CO\
        );

    \I__2537\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18592\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__18592\,
            I => \N__18588\
        );

    \I__2535\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18584\
        );

    \I__2534\ : Span4Mux_s3_h
    port map (
            O => \N__18588\,
            I => \N__18581\
        );

    \I__2533\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18578\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__18584\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__18581\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__18578\,
            I => \b2v_inst20.counterZ0Z_2\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__18571\,
            I => \N__18568\
        );

    \I__2528\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18564\
        );

    \I__2527\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18561\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__18564\,
            I => \b2v_inst200.countZ0Z_1\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__18561\,
            I => \b2v_inst200.countZ0Z_1\
        );

    \I__2524\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18550\
        );

    \I__2523\ : InMux
    port map (
            O => \N__18555\,
            I => \N__18550\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__18550\,
            I => \b2v_inst200.count_RNIC03N_5Z0Z_0\
        );

    \I__2521\ : InMux
    port map (
            O => \N__18547\,
            I => \b2v_inst200.un2_count_1_cry_1_cy\
        );

    \I__2520\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18540\
        );

    \I__2519\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18537\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__18540\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__18537\,
            I => \b2v_inst200.countZ0Z_2\
        );

    \I__2516\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18526\
        );

    \I__2515\ : InMux
    port map (
            O => \N__18531\,
            I => \N__18526\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__18526\,
            I => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\
        );

    \I__2513\ : InMux
    port map (
            O => \N__18523\,
            I => \b2v_inst200.un2_count_1_cry_1\
        );

    \I__2512\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18517\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18514\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__18514\,
            I => \b2v_inst20.un4_counter_0_and\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__18511\,
            I => \b2v_inst11.N_381_cascade_\
        );

    \I__2508\ : InMux
    port map (
            O => \N__18508\,
            I => \N__18505\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__18505\,
            I => \N__18502\
        );

    \I__2506\ : Odrv12
    port map (
            O => \N__18502\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__18499\,
            I => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_\
        );

    \I__2504\ : InMux
    port map (
            O => \N__18496\,
            I => \N__18493\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__18493\,
            I => \N__18490\
        );

    \I__2502\ : Span12Mux_s3_h
    port map (
            O => \N__18490\,
            I => \N__18487\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__18487\,
            I => \b2v_inst11.N_381_0\
        );

    \I__2500\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18481\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__2498\ : Span4Mux_s2_v
    port map (
            O => \N__18478\,
            I => \N__18475\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__18475\,
            I => \N__18472\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__18469\,
            I => \N_15_i_0_a4_0_1\
        );

    \I__2494\ : InMux
    port map (
            O => \N__18466\,
            I => \N__18463\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__18463\,
            I => \N__18460\
        );

    \I__2492\ : Span4Mux_s3_v
    port map (
            O => \N__18460\,
            I => \N__18457\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__18457\,
            I => \b2v_inst20.counter_1_cry_2_THRU_CO\
        );

    \I__2490\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18451\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__18451\,
            I => \N__18447\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__18450\,
            I => \N__18443\
        );

    \I__2487\ : Span4Mux_s3_h
    port map (
            O => \N__18447\,
            I => \N__18440\
        );

    \I__2486\ : InMux
    port map (
            O => \N__18446\,
            I => \N__18435\
        );

    \I__2485\ : InMux
    port map (
            O => \N__18443\,
            I => \N__18435\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__18440\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__18435\,
            I => \b2v_inst20.counterZ0Z_3\
        );

    \I__2482\ : InMux
    port map (
            O => \N__18430\,
            I => \N__18425\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__18429\,
            I => \N__18422\
        );

    \I__2480\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18419\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__18425\,
            I => \N__18416\
        );

    \I__2478\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18413\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__18419\,
            I => \N__18410\
        );

    \I__2476\ : Span4Mux_s3_h
    port map (
            O => \N__18416\,
            I => \N__18407\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18404\
        );

    \I__2474\ : Span4Mux_s3_h
    port map (
            O => \N__18410\,
            I => \N__18401\
        );

    \I__2473\ : Span4Mux_v
    port map (
            O => \N__18407\,
            I => \N__18396\
        );

    \I__2472\ : Span4Mux_s3_h
    port map (
            O => \N__18404\,
            I => \N__18396\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__18401\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__2470\ : Odrv4
    port map (
            O => \N__18396\,
            I => \b2v_inst11.count_clkZ0Z_8\
        );

    \I__2469\ : InMux
    port map (
            O => \N__18391\,
            I => \N__18388\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__18388\,
            I => \N__18385\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__18385\,
            I => \N__18381\
        );

    \I__2466\ : InMux
    port map (
            O => \N__18384\,
            I => \N__18378\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__18381\,
            I => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__18378\,
            I => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\
        );

    \I__2463\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18370\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18367\
        );

    \I__2461\ : Span4Mux_h
    port map (
            O => \N__18367\,
            I => \N__18364\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__18364\,
            I => \b2v_inst11.count_clk_0_2\
        );

    \I__2459\ : InMux
    port map (
            O => \N__18361\,
            I => \N__18357\
        );

    \I__2458\ : InMux
    port map (
            O => \N__18360\,
            I => \N__18353\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__18357\,
            I => \N__18350\
        );

    \I__2456\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18347\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__18353\,
            I => \N__18344\
        );

    \I__2454\ : Span4Mux_h
    port map (
            O => \N__18350\,
            I => \N__18341\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__18347\,
            I => \N__18338\
        );

    \I__2452\ : Span4Mux_s3_h
    port map (
            O => \N__18344\,
            I => \N__18335\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__18341\,
            I => \N__18332\
        );

    \I__2450\ : Span4Mux_s3_h
    port map (
            O => \N__18338\,
            I => \N__18329\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__18335\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__18332\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__18329\,
            I => \b2v_inst11.count_clkZ0Z_2\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__18322\,
            I => \N__18317\
        );

    \I__2445\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18313\
        );

    \I__2444\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18308\
        );

    \I__2443\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18308\
        );

    \I__2442\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18305\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__18313\,
            I => \N__18302\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18299\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__18305\,
            I => \N__18296\
        );

    \I__2438\ : Span4Mux_s3_h
    port map (
            O => \N__18302\,
            I => \N__18293\
        );

    \I__2437\ : Span4Mux_s3_h
    port map (
            O => \N__18299\,
            I => \N__18288\
        );

    \I__2436\ : Span4Mux_s3_h
    port map (
            O => \N__18296\,
            I => \N__18288\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__18293\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__18288\,
            I => \b2v_inst11.count_clkZ0Z_5\
        );

    \I__2433\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18280\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__18280\,
            I => \N__18276\
        );

    \I__2431\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18273\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__18276\,
            I => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__18273\,
            I => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\
        );

    \I__2428\ : InMux
    port map (
            O => \N__18268\,
            I => \N__18265\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__18265\,
            I => \N__18262\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__18262\,
            I => \b2v_inst11.count_clk_0_9\
        );

    \I__2425\ : InMux
    port map (
            O => \N__18259\,
            I => \N__18249\
        );

    \I__2424\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18249\
        );

    \I__2423\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18249\
        );

    \I__2422\ : InMux
    port map (
            O => \N__18256\,
            I => \N__18246\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__18249\,
            I => \N__18243\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__18246\,
            I => \N__18240\
        );

    \I__2419\ : Span4Mux_s3_h
    port map (
            O => \N__18243\,
            I => \N__18237\
        );

    \I__2418\ : Odrv4
    port map (
            O => \N__18240\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__18237\,
            I => \b2v_inst11.count_clkZ0Z_9\
        );

    \I__2416\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18228\
        );

    \I__2415\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18225\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__18228\,
            I => \N__18220\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__18225\,
            I => \N__18220\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__18217\,
            I => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\
        );

    \I__2410\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18211\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__18211\,
            I => \b2v_inst11.count_clk_0_3\
        );

    \I__2408\ : InMux
    port map (
            O => \N__18208\,
            I => \N__18204\
        );

    \I__2407\ : InMux
    port map (
            O => \N__18207\,
            I => \N__18201\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__18204\,
            I => \N__18198\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__18201\,
            I => \N__18195\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__18198\,
            I => \N__18192\
        );

    \I__2403\ : Span4Mux_h
    port map (
            O => \N__18195\,
            I => \N__18189\
        );

    \I__2402\ : Odrv4
    port map (
            O => \N__18192\,
            I => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__18189\,
            I => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\
        );

    \I__2400\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18181\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__18181\,
            I => \b2v_inst11.count_clk_0_5\
        );

    \I__2398\ : InMux
    port map (
            O => \N__18178\,
            I => \N__18174\
        );

    \I__2397\ : InMux
    port map (
            O => \N__18177\,
            I => \N__18171\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__18174\,
            I => \N__18168\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__18171\,
            I => \N__18165\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__18168\,
            I => \N__18162\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__18165\,
            I => \N__18159\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__18162\,
            I => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__18159\,
            I => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\
        );

    \I__2390\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18151\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__18151\,
            I => \b2v_inst11.count_clk_0_6\
        );

    \I__2388\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18144\
        );

    \I__2387\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18141\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__18144\,
            I => \N__18138\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__18138\,
            I => \N__18132\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__18135\,
            I => \N__18129\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__18132\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__18129\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\
        );

    \I__2380\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__18121\,
            I => \b2v_inst11.count_clk_0_8\
        );

    \I__2378\ : CEMux
    port map (
            O => \N__18118\,
            I => \N__18115\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__18115\,
            I => \N__18108\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \N__18103\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__18113\,
            I => \N__18099\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \N__18096\
        );

    \I__2373\ : CEMux
    port map (
            O => \N__18111\,
            I => \N__18092\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__18108\,
            I => \N__18088\
        );

    \I__2371\ : CEMux
    port map (
            O => \N__18107\,
            I => \N__18085\
        );

    \I__2370\ : InMux
    port map (
            O => \N__18106\,
            I => \N__18069\
        );

    \I__2369\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18069\
        );

    \I__2368\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18069\
        );

    \I__2367\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18069\
        );

    \I__2366\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18069\
        );

    \I__2365\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18069\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18065\
        );

    \I__2363\ : CEMux
    port map (
            O => \N__18091\,
            I => \N__18062\
        );

    \I__2362\ : Span4Mux_h
    port map (
            O => \N__18088\,
            I => \N__18057\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__18085\,
            I => \N__18057\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__18084\,
            I => \N__18051\
        );

    \I__2359\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18043\
        );

    \I__2358\ : CEMux
    port map (
            O => \N__18082\,
            I => \N__18043\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__18069\,
            I => \N__18040\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__18068\,
            I => \N__18037\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__18065\,
            I => \N__18034\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__18062\,
            I => \N__18031\
        );

    \I__2353\ : Span4Mux_s1_h
    port map (
            O => \N__18057\,
            I => \N__18028\
        );

    \I__2352\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18021\
        );

    \I__2351\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18021\
        );

    \I__2350\ : InMux
    port map (
            O => \N__18054\,
            I => \N__18021\
        );

    \I__2349\ : InMux
    port map (
            O => \N__18051\,
            I => \N__18018\
        );

    \I__2348\ : InMux
    port map (
            O => \N__18050\,
            I => \N__18011\
        );

    \I__2347\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18011\
        );

    \I__2346\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18011\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__18043\,
            I => \N__18006\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__18040\,
            I => \N__18006\
        );

    \I__2343\ : InMux
    port map (
            O => \N__18037\,
            I => \N__18003\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__18034\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__18031\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__18028\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__18021\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__18018\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__18011\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__18006\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__18003\,
            I => \b2v_inst11.count_clk_en\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__17986\,
            I => \N__17983\
        );

    \I__2333\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17980\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__17980\,
            I => \N__17977\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__17977\,
            I => \N__17974\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__17974\,
            I => \func_state_RNIVS8U1_4_1\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \N__17968\
        );

    \I__2328\ : InMux
    port map (
            O => \N__17968\,
            I => \N__17962\
        );

    \I__2327\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17962\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__17962\,
            I => \b2v_inst11.func_stateZ0Z_1\
        );

    \I__2325\ : InMux
    port map (
            O => \N__17959\,
            I => \N__17956\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__17956\,
            I => \N__17952\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \N__17949\
        );

    \I__2322\ : Span4Mux_s3_h
    port map (
            O => \N__17952\,
            I => \N__17943\
        );

    \I__2321\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17938\
        );

    \I__2320\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17938\
        );

    \I__2319\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17933\
        );

    \I__2318\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17933\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__17943\,
            I => \b2v_inst11.count_clk_enZ0Z_0\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__17938\,
            I => \b2v_inst11.count_clk_enZ0Z_0\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__17933\,
            I => \b2v_inst11.count_clk_enZ0Z_0\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__17926\,
            I => \VCCST_EN_i_0_o3_0_cascade_\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17923\,
            I => \N__17917\
        );

    \I__2312\ : InMux
    port map (
            O => \N__17922\,
            I => \N__17917\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__17917\,
            I => \b2v_inst11.func_state_1_m2_1\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__17914\,
            I => \func_state_RNI6BE8E_0_1_cascade_\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17908\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__17908\,
            I => \b2v_inst11.count_0_7\
        );

    \I__2307\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17900\
        );

    \I__2306\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17897\
        );

    \I__2305\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17894\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__17900\,
            I => \N__17891\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__17897\,
            I => \N__17886\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__17894\,
            I => \N__17886\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__17891\,
            I => \N__17883\
        );

    \I__2300\ : Span4Mux_s3_h
    port map (
            O => \N__17886\,
            I => \N__17880\
        );

    \I__2299\ : Odrv4
    port map (
            O => \N__17883\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__17880\,
            I => \b2v_inst11.count_clkZ0Z_3\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17871\
        );

    \I__2296\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17867\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17864\
        );

    \I__2294\ : InMux
    port map (
            O => \N__17870\,
            I => \N__17861\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__17867\,
            I => \N__17856\
        );

    \I__2292\ : Span4Mux_s2_h
    port map (
            O => \N__17864\,
            I => \N__17856\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17853\
        );

    \I__2290\ : Span4Mux_v
    port map (
            O => \N__17856\,
            I => \N__17850\
        );

    \I__2289\ : Span4Mux_s3_h
    port map (
            O => \N__17853\,
            I => \N__17847\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__17850\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__17847\,
            I => \b2v_inst11.count_clkZ0Z_6\
        );

    \I__2286\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17838\
        );

    \I__2285\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17835\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17831\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__17835\,
            I => \N__17828\
        );

    \I__2282\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17825\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__17831\,
            I => \N__17822\
        );

    \I__2280\ : Span12Mux_s7_v
    port map (
            O => \N__17828\,
            I => \N__17819\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__17825\,
            I => \N__17816\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__17822\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__2277\ : Odrv12
    port map (
            O => \N__17819\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__2276\ : Odrv12
    port map (
            O => \N__17816\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__17809\,
            I => \b2v_inst11.func_state_1_m2_am_1_1_cascade_\
        );

    \I__2274\ : InMux
    port map (
            O => \N__17806\,
            I => \N__17803\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__17803\,
            I => \N__17800\
        );

    \I__2272\ : Span4Mux_h
    port map (
            O => \N__17800\,
            I => \N__17794\
        );

    \I__2271\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17787\
        );

    \I__2270\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17787\
        );

    \I__2269\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17787\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__17794\,
            I => \b2v_inst11.count_off_RNIZ0Z_9\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__17787\,
            I => \b2v_inst11.count_off_RNIZ0Z_9\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__17782\,
            I => \b2v_inst11.func_state_RNIR5S85Z0Z_1_cascade_\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__17779\,
            I => \b2v_inst11.func_state_cascade_\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__17776\,
            I => \N__17772\
        );

    \I__2263\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17767\
        );

    \I__2262\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17767\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__17767\,
            I => \b2v_inst11.func_stateZ0Z_0\
        );

    \I__2260\ : InMux
    port map (
            O => \N__17764\,
            I => \N__17758\
        );

    \I__2259\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17758\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__17758\,
            I => \N__17755\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__17755\,
            I => \b2v_inst11.N_160_i\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__17752\,
            I => \N__17747\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__17751\,
            I => \N__17742\
        );

    \I__2254\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17737\
        );

    \I__2253\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17731\
        );

    \I__2252\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17731\
        );

    \I__2251\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17728\
        );

    \I__2250\ : InMux
    port map (
            O => \N__17742\,
            I => \N__17720\
        );

    \I__2249\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17720\
        );

    \I__2248\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17720\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__17737\,
            I => \N__17717\
        );

    \I__2246\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17714\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__17731\,
            I => \N__17711\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__17728\,
            I => \N__17708\
        );

    \I__2243\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17705\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__17720\,
            I => \N__17702\
        );

    \I__2241\ : Span12Mux_s10_v
    port map (
            O => \N__17717\,
            I => \N__17699\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__17714\,
            I => \N__17696\
        );

    \I__2239\ : Span4Mux_s3_h
    port map (
            O => \N__17711\,
            I => \N__17693\
        );

    \I__2238\ : Span4Mux_s3_h
    port map (
            O => \N__17708\,
            I => \N__17690\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__17705\,
            I => \N__17685\
        );

    \I__2236\ : Span4Mux_s3_h
    port map (
            O => \N__17702\,
            I => \N__17685\
        );

    \I__2235\ : Odrv12
    port map (
            O => \N__17699\,
            I => \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\
        );

    \I__2234\ : Odrv12
    port map (
            O => \N__17696\,
            I => \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__17693\,
            I => \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__17690\,
            I => \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__17685\,
            I => \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\
        );

    \I__2230\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17671\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17668\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__17668\,
            I => \b2v_inst11.func_state_1_m0_0_1_0\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__17665\,
            I => \b2v_inst11.func_state_1_m2_1_0_cascade_\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__17662\,
            I => \N__17658\
        );

    \I__2225\ : InMux
    port map (
            O => \N__17661\,
            I => \N__17650\
        );

    \I__2224\ : InMux
    port map (
            O => \N__17658\,
            I => \N__17650\
        );

    \I__2223\ : InMux
    port map (
            O => \N__17657\,
            I => \N__17650\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__17650\,
            I => \b2v_inst11.N_76\
        );

    \I__2221\ : InMux
    port map (
            O => \N__17647\,
            I => \N__17641\
        );

    \I__2220\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17641\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__17641\,
            I => \b2v_inst11.func_state_1_m2_0\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_\
        );

    \I__2217\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17632\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17629\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__17629\,
            I => \N__17626\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__17626\,
            I => \b2v_inst11.N_337\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__17623\,
            I => \b2v_inst11.func_state_1_m2s2_i_0_cascade_\
        );

    \I__2212\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17614\
        );

    \I__2210\ : Span4Mux_h
    port map (
            O => \N__17614\,
            I => \N__17611\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__17611\,
            I => \b2v_inst11.N_338\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__17608\,
            I => \b2v_inst11.dutycycle_RNI_5Z0Z_6_cascade_\
        );

    \I__2207\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17602\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__2205\ : Odrv4
    port map (
            O => \N__17599\,
            I => \b2v_inst11.N_231_N\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__17596\,
            I => \b2v_inst11.N_306_cascade_\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__17593\,
            I => \b2v_inst11.N_354_cascade_\
        );

    \I__2202\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__2200\ : Odrv4
    port map (
            O => \N__17584\,
            I => b2v_inst11_g0_i_m2_i_a6_3_2
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__17581\,
            I => \b2v_inst11.N_159_cascade_\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__17578\,
            I => \b2v_inst11.func_state_1_m0_0_1_1_0_cascade_\
        );

    \I__2197\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17572\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17569\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__17569\,
            I => \N__17566\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__17566\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_313_N\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__17563\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_sx_cascade_\
        );

    \I__2192\ : InMux
    port map (
            O => \N__17560\,
            I => \N__17557\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__17557\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1\
        );

    \I__2190\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17549\
        );

    \I__2189\ : InMux
    port map (
            O => \N__17553\,
            I => \N__17544\
        );

    \I__2188\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17544\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__17549\,
            I => \b2v_inst11.dutycycleZ1Z_7\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__17544\,
            I => \b2v_inst11.dutycycleZ1Z_7\
        );

    \I__2185\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17535\
        );

    \I__2184\ : InMux
    port map (
            O => \N__17538\,
            I => \N__17532\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__17535\,
            I => \N__17527\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__17532\,
            I => \N__17527\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__17527\,
            I => \b2v_inst11.dutycycle_RNI24DD8Z0Z_7\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__17524\,
            I => \b2v_inst11.dutycycle_RNIVGS13Z0Z_7_cascade_\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__17521\,
            I => \b2v_inst11.N_160_i_cascade_\
        );

    \I__2178\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17515\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__17515\,
            I => \N__17512\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__17512\,
            I => \b2v_inst11.g1_0_sx\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__17509\,
            I => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_0_cascade_\
        );

    \I__2174\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17503\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__17503\,
            I => \N__17500\
        );

    \I__2172\ : Span4Mux_v
    port map (
            O => \N__17500\,
            I => \N__17497\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__17497\,
            I => \b2v_inst11.func_state_RNI608H1_0Z0Z_1\
        );

    \I__2170\ : InMux
    port map (
            O => \N__17494\,
            I => \N__17488\
        );

    \I__2169\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17488\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17485\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__17485\,
            I => \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__17482\,
            I => \N__17479\
        );

    \I__2165\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17476\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__17476\,
            I => \b2v_inst11.count_off_0_12\
        );

    \I__2163\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17469\
        );

    \I__2162\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17466\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__17469\,
            I => \b2v_inst11.count_offZ0Z_12\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__17466\,
            I => \b2v_inst11.count_offZ0Z_12\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__17461\,
            I => \N__17458\
        );

    \I__2158\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17455\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__17455\,
            I => \N__17451\
        );

    \I__2156\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17448\
        );

    \I__2155\ : Span4Mux_h
    port map (
            O => \N__17451\,
            I => \N__17445\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__17448\,
            I => \N__17442\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__17445\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__2152\ : Odrv4
    port map (
            O => \N__17442\,
            I => \b2v_inst11.count_offZ0Z_10\
        );

    \I__2151\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17434\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__17434\,
            I => \b2v_inst11.un34_clk_100khz_5\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__17431\,
            I => \b2v_inst11.un34_clk_100khz_4_cascade_\
        );

    \I__2148\ : InMux
    port map (
            O => \N__17428\,
            I => \N__17425\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__17425\,
            I => \N__17422\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__17422\,
            I => \b2v_inst11.un34_clk_100khz_11\
        );

    \I__2145\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__2144\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17413\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__17413\,
            I => \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\
        );

    \I__2142\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17404\
        );

    \I__2141\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17404\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__17404\,
            I => \b2v_inst11.count_offZ0Z_11\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \b2v_inst11.g4_cascade_\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__17398\,
            I => \b2v_inst11.g0_17_N_3L3_1_cascade_\
        );

    \I__2137\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17392\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__17392\,
            I => \b2v_inst11.dutycycle_RNIVGS13Z0Z_7\
        );

    \I__2135\ : InMux
    port map (
            O => \N__17389\,
            I => \b2v_inst11.un3_count_off_1_cry_11\
        );

    \I__2134\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17383\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__17383\,
            I => \N__17380\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__17380\,
            I => \b2v_inst11.count_offZ0Z_13\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \N__17374\
        );

    \I__2130\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17370\
        );

    \I__2129\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17367\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__17370\,
            I => \N__17364\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__17367\,
            I => \N__17361\
        );

    \I__2126\ : Odrv12
    port map (
            O => \N__17364\,
            I => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__17361\,
            I => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\
        );

    \I__2124\ : InMux
    port map (
            O => \N__17356\,
            I => \b2v_inst11.un3_count_off_1_cry_12\
        );

    \I__2123\ : InMux
    port map (
            O => \N__17353\,
            I => \b2v_inst11.un3_count_off_1_cry_13\
        );

    \I__2122\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17347\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__17347\,
            I => \N__17343\
        );

    \I__2120\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17340\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__17343\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__17340\,
            I => \b2v_inst11.count_offZ0Z_15\
        );

    \I__2117\ : InMux
    port map (
            O => \N__17335\,
            I => \b2v_inst11.un3_count_off_1_cry_14\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__17332\,
            I => \N__17329\
        );

    \I__2115\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17323\
        );

    \I__2114\ : InMux
    port map (
            O => \N__17328\,
            I => \N__17323\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__17323\,
            I => \N__17320\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__17320\,
            I => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\
        );

    \I__2111\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17314\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__17314\,
            I => \b2v_inst11.un3_count_off_1_axb_11\
        );

    \I__2109\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17308\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__17308\,
            I => \b2v_inst11.count_off_1_11\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__17305\,
            I => \b2v_inst11.count_off_1_11_cascade_\
        );

    \I__2106\ : InMux
    port map (
            O => \N__17302\,
            I => \b2v_inst11.un3_count_off_1_cry_3\
        );

    \I__2105\ : InMux
    port map (
            O => \N__17299\,
            I => \b2v_inst11.un3_count_off_1_cry_4\
        );

    \I__2104\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17293\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__17293\,
            I => \N__17290\
        );

    \I__2102\ : Span4Mux_h
    port map (
            O => \N__17290\,
            I => \N__17287\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__17287\,
            I => \N__17284\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__17284\,
            I => \b2v_inst11.un3_count_off_1_axb_6\
        );

    \I__2099\ : InMux
    port map (
            O => \N__17281\,
            I => \b2v_inst11.un3_count_off_1_cry_5\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__17278\,
            I => \N__17275\
        );

    \I__2097\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17272\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__17272\,
            I => \b2v_inst11.un3_count_off_1_axb_7\
        );

    \I__2095\ : InMux
    port map (
            O => \N__17269\,
            I => \b2v_inst11.un3_count_off_1_cry_6\
        );

    \I__2094\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17263\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__17263\,
            I => \b2v_inst11.count_offZ0Z_8\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__17260\,
            I => \N__17257\
        );

    \I__2091\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17251\
        );

    \I__2090\ : InMux
    port map (
            O => \N__17256\,
            I => \N__17251\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__17251\,
            I => \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\
        );

    \I__2088\ : InMux
    port map (
            O => \N__17248\,
            I => \b2v_inst11.un3_count_off_1_cry_7\
        );

    \I__2087\ : InMux
    port map (
            O => \N__17245\,
            I => \bfn_4_5_0_\
        );

    \I__2086\ : InMux
    port map (
            O => \N__17242\,
            I => \N__17238\
        );

    \I__2085\ : InMux
    port map (
            O => \N__17241\,
            I => \N__17235\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__17238\,
            I => \N__17230\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__17235\,
            I => \N__17230\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__17230\,
            I => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\
        );

    \I__2081\ : InMux
    port map (
            O => \N__17227\,
            I => \b2v_inst11.un3_count_off_1_cry_9\
        );

    \I__2080\ : InMux
    port map (
            O => \N__17224\,
            I => \b2v_inst11.un3_count_off_1_cry_10\
        );

    \I__2079\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17218\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__17218\,
            I => \b2v_inst11.count_off_0_15\
        );

    \I__2077\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17212\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__17212\,
            I => \N__17209\
        );

    \I__2075\ : Span4Mux_h
    port map (
            O => \N__17209\,
            I => \N__17206\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__17206\,
            I => \b2v_inst11.count_off_0_13\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__17203\,
            I => \b2v_inst11.count_offZ0Z_13_cascade_\
        );

    \I__2072\ : InMux
    port map (
            O => \N__17200\,
            I => \N__17197\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__17197\,
            I => \b2v_inst11.count_off_0_8\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__17194\,
            I => \b2v_inst11.count_offZ0Z_8_cascade_\
        );

    \I__2069\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17187\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__17190\,
            I => \N__17184\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__17187\,
            I => \N__17181\
        );

    \I__2066\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17178\
        );

    \I__2065\ : Span4Mux_v
    port map (
            O => \N__17181\,
            I => \N__17175\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__17178\,
            I => \N__17172\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__17175\,
            I => \N__17165\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__17172\,
            I => \N__17165\
        );

    \I__2061\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17160\
        );

    \I__2060\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17160\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__17165\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__17160\,
            I => \b2v_inst11.count_offZ0Z_0\
        );

    \I__2057\ : InMux
    port map (
            O => \N__17155\,
            I => \b2v_inst11.un3_count_off_1_cry_1\
        );

    \I__2056\ : InMux
    port map (
            O => \N__17152\,
            I => \b2v_inst11.un3_count_off_1_cry_2\
        );

    \I__2055\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17146\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__17146\,
            I => \b2v_inst200.count_3_3\
        );

    \I__2053\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17140\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__17140\,
            I => \N__17137\
        );

    \I__2051\ : Odrv12
    port map (
            O => \N__17137\,
            I => \b2v_inst200.count_3_12\
        );

    \I__2050\ : InMux
    port map (
            O => \N__17134\,
            I => \N__17131\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__17131\,
            I => \b2v_inst200.count_3_4\
        );

    \I__2048\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__2046\ : Odrv12
    port map (
            O => \N__17122\,
            I => \b2v_inst200.count_3_5\
        );

    \I__2045\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__17116\,
            I => \N__17113\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__17113\,
            I => \b2v_inst200.count_3_7\
        );

    \I__2042\ : InMux
    port map (
            O => \N__17110\,
            I => \bfn_2_16_0_\
        );

    \I__2041\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17103\
        );

    \I__2040\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__17103\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__17100\,
            I => \b2v_inst20.counterZ0Z_31\
        );

    \I__2037\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17091\
        );

    \I__2036\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17088\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__17091\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__17088\,
            I => \b2v_inst20.counterZ0Z_29\
        );

    \I__2033\ : CascadeMux
    port map (
            O => \N__17083\,
            I => \N__17079\
        );

    \I__2032\ : InMux
    port map (
            O => \N__17082\,
            I => \N__17076\
        );

    \I__2031\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17073\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__17076\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__17073\,
            I => \b2v_inst20.counterZ0Z_30\
        );

    \I__2028\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17064\
        );

    \I__2027\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17061\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__17064\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__17061\,
            I => \b2v_inst20.counterZ0Z_28\
        );

    \I__2024\ : InMux
    port map (
            O => \N__17056\,
            I => \N__17053\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__17053\,
            I => \b2v_inst20.un4_counter_7_and\
        );

    \I__2022\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17046\
        );

    \I__2021\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17043\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__17046\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__17043\,
            I => \b2v_inst20.counterZ0Z_27\
        );

    \I__2018\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17034\
        );

    \I__2017\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17031\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__17034\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__17031\,
            I => \b2v_inst20.counterZ0Z_25\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__17026\,
            I => \N__17022\
        );

    \I__2013\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17019\
        );

    \I__2012\ : InMux
    port map (
            O => \N__17022\,
            I => \N__17016\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__17019\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__17016\,
            I => \b2v_inst20.counterZ0Z_26\
        );

    \I__2009\ : InMux
    port map (
            O => \N__17011\,
            I => \N__17007\
        );

    \I__2008\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17004\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__17007\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__17004\,
            I => \b2v_inst20.counterZ0Z_24\
        );

    \I__2005\ : InMux
    port map (
            O => \N__16999\,
            I => \N__16996\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__16996\,
            I => \b2v_inst20.un4_counter_6_and\
        );

    \I__2003\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16990\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__16990\,
            I => \b2v_inst200.count_3_1\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16984\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__16984\,
            I => \b2v_inst200.count_3_2\
        );

    \I__1999\ : InMux
    port map (
            O => \N__16981\,
            I => \N__16978\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__16978\,
            I => \N__16975\
        );

    \I__1997\ : IoSpan4Mux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__1996\ : IoSpan4Mux
    port map (
            O => \N__16972\,
            I => \N__16969\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__16969\,
            I => \VPP_OK_c\
        );

    \I__1994\ : IoInMux
    port map (
            O => \N__16966\,
            I => \N__16963\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__16963\,
            I => \N__16960\
        );

    \I__1992\ : Odrv12
    port map (
            O => \N__16960\,
            I => \VDDQ_EN_c\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__16957\,
            I => \N__16954\
        );

    \I__1990\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16951\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__16951\,
            I => \b2v_inst20.un4_counter_2_and\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__16948\,
            I => \N__16945\
        );

    \I__1987\ : InMux
    port map (
            O => \N__16945\,
            I => \N__16942\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__16942\,
            I => \b2v_inst20.un4_counter_3_and\
        );

    \I__1985\ : InMux
    port map (
            O => \N__16939\,
            I => \N__16936\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__16936\,
            I => \b2v_inst20.un4_counter_4_and\
        );

    \I__1983\ : InMux
    port map (
            O => \N__16933\,
            I => \N__16930\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__16930\,
            I => \b2v_inst20.un4_counter_5_and\
        );

    \I__1981\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16923\
        );

    \I__1980\ : InMux
    port map (
            O => \N__16926\,
            I => \N__16920\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__16923\,
            I => \N__16917\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__16920\,
            I => \N__16914\
        );

    \I__1977\ : Span4Mux_s1_h
    port map (
            O => \N__16917\,
            I => \N__16911\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__16914\,
            I => \b2v_inst11.count_clk_1_14\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__16911\,
            I => \b2v_inst11.count_clk_1_14\
        );

    \I__1974\ : InMux
    port map (
            O => \N__16906\,
            I => \b2v_inst11.un1_count_clk_2_cry_13\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16903\,
            I => \N__16900\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__16900\,
            I => \N__16896\
        );

    \I__1971\ : InMux
    port map (
            O => \N__16899\,
            I => \N__16893\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__16896\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__16893\,
            I => \b2v_inst11.count_clkZ0Z_15\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__16888\,
            I => \N__16881\
        );

    \I__1967\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16862\
        );

    \I__1966\ : InMux
    port map (
            O => \N__16886\,
            I => \N__16859\
        );

    \I__1965\ : InMux
    port map (
            O => \N__16885\,
            I => \N__16852\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16852\
        );

    \I__1963\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16852\
        );

    \I__1962\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16845\
        );

    \I__1961\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16845\
        );

    \I__1960\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16845\
        );

    \I__1959\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16838\
        );

    \I__1958\ : InMux
    port map (
            O => \N__16876\,
            I => \N__16838\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16838\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16874\,
            I => \N__16831\
        );

    \I__1955\ : InMux
    port map (
            O => \N__16873\,
            I => \N__16831\
        );

    \I__1954\ : InMux
    port map (
            O => \N__16872\,
            I => \N__16831\
        );

    \I__1953\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16816\
        );

    \I__1952\ : InMux
    port map (
            O => \N__16870\,
            I => \N__16816\
        );

    \I__1951\ : InMux
    port map (
            O => \N__16869\,
            I => \N__16816\
        );

    \I__1950\ : InMux
    port map (
            O => \N__16868\,
            I => \N__16816\
        );

    \I__1949\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16816\
        );

    \I__1948\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16816\
        );

    \I__1947\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16816\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__16862\,
            I => \N__16809\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__16859\,
            I => \N__16809\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__16852\,
            I => \N__16809\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__16845\,
            I => \b2v_inst11.func_state_RNICGI84_0_0\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__16838\,
            I => \b2v_inst11.func_state_RNICGI84_0_0\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__16831\,
            I => \b2v_inst11.func_state_RNICGI84_0_0\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__16816\,
            I => \b2v_inst11.func_state_RNICGI84_0_0\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__16809\,
            I => \b2v_inst11.func_state_RNICGI84_0_0\
        );

    \I__1938\ : InMux
    port map (
            O => \N__16798\,
            I => \b2v_inst11.un1_count_clk_2_cry_14\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__16795\,
            I => \N__16791\
        );

    \I__1936\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16786\
        );

    \I__1935\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16786\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__16786\,
            I => \N__16783\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__16783\,
            I => \b2v_inst11.count_clk_1_15\
        );

    \I__1932\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16776\
        );

    \I__1931\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16773\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__16776\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__16773\,
            I => \b2v_inst20.counterZ0Z_11\
        );

    \I__1928\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16764\
        );

    \I__1927\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16761\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__16764\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__16761\,
            I => \b2v_inst20.counterZ0Z_9\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__16756\,
            I => \N__16752\
        );

    \I__1923\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16749\
        );

    \I__1922\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16746\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__16749\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__16746\,
            I => \b2v_inst20.counterZ0Z_10\
        );

    \I__1919\ : InMux
    port map (
            O => \N__16741\,
            I => \N__16737\
        );

    \I__1918\ : InMux
    port map (
            O => \N__16740\,
            I => \N__16734\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__16737\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__16734\,
            I => \b2v_inst20.counterZ0Z_8\
        );

    \I__1915\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16725\
        );

    \I__1914\ : InMux
    port map (
            O => \N__16728\,
            I => \N__16722\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__16725\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__16722\,
            I => \b2v_inst20.counterZ0Z_15\
        );

    \I__1911\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16713\
        );

    \I__1910\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16710\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__16713\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__16710\,
            I => \b2v_inst20.counterZ0Z_14\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__16705\,
            I => \N__16701\
        );

    \I__1906\ : InMux
    port map (
            O => \N__16704\,
            I => \N__16698\
        );

    \I__1905\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16695\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__16698\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__16695\,
            I => \b2v_inst20.counterZ0Z_13\
        );

    \I__1902\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16686\
        );

    \I__1901\ : InMux
    port map (
            O => \N__16689\,
            I => \N__16683\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__16686\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__16683\,
            I => \b2v_inst20.counterZ0Z_12\
        );

    \I__1898\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16674\
        );

    \I__1897\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16671\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__16674\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__16671\,
            I => \b2v_inst20.counterZ0Z_19\
        );

    \I__1894\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16662\
        );

    \I__1893\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16659\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__16662\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__16659\,
            I => \b2v_inst20.counterZ0Z_17\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__16654\,
            I => \N__16650\
        );

    \I__1889\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16647\
        );

    \I__1888\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16644\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__16647\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__16644\,
            I => \b2v_inst20.counterZ0Z_18\
        );

    \I__1885\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16635\
        );

    \I__1884\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16632\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__16635\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__16632\,
            I => \b2v_inst20.counterZ0Z_16\
        );

    \I__1881\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16623\
        );

    \I__1880\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16620\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__16623\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__16620\,
            I => \b2v_inst20.counterZ0Z_23\
        );

    \I__1877\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16611\
        );

    \I__1876\ : InMux
    port map (
            O => \N__16614\,
            I => \N__16608\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__16611\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__16608\,
            I => \b2v_inst20.counterZ0Z_21\
        );

    \I__1873\ : CascadeMux
    port map (
            O => \N__16603\,
            I => \N__16599\
        );

    \I__1872\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16596\
        );

    \I__1871\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16593\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__16596\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__16593\,
            I => \b2v_inst20.counterZ0Z_22\
        );

    \I__1868\ : InMux
    port map (
            O => \N__16588\,
            I => \N__16584\
        );

    \I__1867\ : InMux
    port map (
            O => \N__16587\,
            I => \N__16581\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__16584\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__16581\,
            I => \b2v_inst20.counterZ0Z_20\
        );

    \I__1864\ : InMux
    port map (
            O => \N__16576\,
            I => \b2v_inst11.un1_count_clk_2_cry_5\
        );

    \I__1863\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16569\
        );

    \I__1862\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16563\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16560\
        );

    \I__1860\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16555\
        );

    \I__1859\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16555\
        );

    \I__1858\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16552\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__16563\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__16560\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__16555\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__16552\,
            I => \b2v_inst11.count_clkZ0Z_7\
        );

    \I__1853\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16537\
        );

    \I__1852\ : InMux
    port map (
            O => \N__16542\,
            I => \N__16537\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__16537\,
            I => \N__16534\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__16534\,
            I => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\
        );

    \I__1849\ : InMux
    port map (
            O => \N__16531\,
            I => \b2v_inst11.un1_count_clk_2_cry_6\
        );

    \I__1848\ : InMux
    port map (
            O => \N__16528\,
            I => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\
        );

    \I__1847\ : InMux
    port map (
            O => \N__16525\,
            I => \bfn_2_13_0_\
        );

    \I__1846\ : InMux
    port map (
            O => \N__16522\,
            I => \N__16519\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__16519\,
            I => \b2v_inst11.count_clkZ0Z_10\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__16516\,
            I => \N__16513\
        );

    \I__1843\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16507\
        );

    \I__1842\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16507\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__16507\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\
        );

    \I__1840\ : InMux
    port map (
            O => \N__16504\,
            I => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\
        );

    \I__1839\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16497\
        );

    \I__1838\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16494\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__16497\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__16494\,
            I => \b2v_inst11.count_clkZ0Z_11\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__16489\,
            I => \N__16486\
        );

    \I__1834\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16480\
        );

    \I__1833\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16480\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__16480\,
            I => \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0\
        );

    \I__1831\ : InMux
    port map (
            O => \N__16477\,
            I => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\
        );

    \I__1830\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16470\
        );

    \I__1829\ : InMux
    port map (
            O => \N__16473\,
            I => \N__16467\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__16470\,
            I => \b2v_inst11.count_clkZ0Z_12\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__16467\,
            I => \b2v_inst11.count_clkZ0Z_12\
        );

    \I__1826\ : InMux
    port map (
            O => \N__16462\,
            I => \N__16456\
        );

    \I__1825\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16456\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__16456\,
            I => \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0\
        );

    \I__1823\ : InMux
    port map (
            O => \N__16453\,
            I => \b2v_inst11.un1_count_clk_2_cry_11\
        );

    \I__1822\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16446\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__16449\,
            I => \N__16442\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16439\
        );

    \I__1819\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16434\
        );

    \I__1818\ : InMux
    port map (
            O => \N__16442\,
            I => \N__16434\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__16439\,
            I => \b2v_inst11.count_clkZ0Z_13\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__16434\,
            I => \b2v_inst11.count_clkZ0Z_13\
        );

    \I__1815\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16423\
        );

    \I__1814\ : InMux
    port map (
            O => \N__16428\,
            I => \N__16423\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__16423\,
            I => \N__16420\
        );

    \I__1812\ : Span4Mux_s1_h
    port map (
            O => \N__16420\,
            I => \N__16417\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__16417\,
            I => \b2v_inst11.count_clk_1_13\
        );

    \I__1810\ : InMux
    port map (
            O => \N__16414\,
            I => \b2v_inst11.un1_count_clk_2_cry_12\
        );

    \I__1809\ : InMux
    port map (
            O => \N__16411\,
            I => \N__16408\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__16408\,
            I => \N__16403\
        );

    \I__1807\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16398\
        );

    \I__1806\ : InMux
    port map (
            O => \N__16406\,
            I => \N__16398\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__16403\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__16398\,
            I => \b2v_inst11.count_clkZ0Z_14\
        );

    \I__1803\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16390\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__16390\,
            I => \b2v_inst11.count_clk_0_14\
        );

    \I__1801\ : InMux
    port map (
            O => \N__16387\,
            I => \N__16384\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__16384\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_2\
        );

    \I__1799\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16378\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__16378\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_3\
        );

    \I__1797\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16371\
        );

    \I__1796\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16365\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__16371\,
            I => \N__16362\
        );

    \I__1794\ : InMux
    port map (
            O => \N__16370\,
            I => \N__16359\
        );

    \I__1793\ : InMux
    port map (
            O => \N__16369\,
            I => \N__16356\
        );

    \I__1792\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16353\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__16365\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__16362\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__16359\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__16356\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__16353\,
            I => \b2v_inst11.count_clkZ0Z_1\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__16342\,
            I => \N__16338\
        );

    \I__1785\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16331\
        );

    \I__1784\ : InMux
    port map (
            O => \N__16338\,
            I => \N__16327\
        );

    \I__1783\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16324\
        );

    \I__1782\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16317\
        );

    \I__1781\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16317\
        );

    \I__1780\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16317\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16314\
        );

    \I__1778\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16311\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__16327\,
            I => \N__16308\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__16324\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__16317\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__16314\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__16311\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__16308\,
            I => \b2v_inst11.count_clkZ0Z_0\
        );

    \I__1771\ : InMux
    port map (
            O => \N__16297\,
            I => \b2v_inst11.un1_count_clk_2_cry_1\
        );

    \I__1770\ : InMux
    port map (
            O => \N__16294\,
            I => \b2v_inst11.un1_count_clk_2_cry_2\
        );

    \I__1769\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16288\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__16288\,
            I => \N__16283\
        );

    \I__1767\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16278\
        );

    \I__1766\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16278\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__16283\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__16278\,
            I => \b2v_inst11.count_clkZ0Z_4\
        );

    \I__1763\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16270\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__16270\,
            I => \N__16267\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__16267\,
            I => \N__16263\
        );

    \I__1760\ : InMux
    port map (
            O => \N__16266\,
            I => \N__16260\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__16263\,
            I => \N__16255\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__16260\,
            I => \N__16255\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__16255\,
            I => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\
        );

    \I__1756\ : InMux
    port map (
            O => \N__16252\,
            I => \b2v_inst11.un1_count_clk_2_cry_3\
        );

    \I__1755\ : InMux
    port map (
            O => \N__16249\,
            I => \b2v_inst11.un1_count_clk_2_cry_4\
        );

    \I__1754\ : InMux
    port map (
            O => \N__16246\,
            I => \N__16243\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__16243\,
            I => \b2v_inst11.count_clk_0_0\
        );

    \I__1752\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16237\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__16237\,
            I => \b2v_inst11.count_clk_0_7\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__16234\,
            I => \b2v_inst11.N_168_cascade_\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__16231\,
            I => \b2v_inst11.func_state_RNICGI84_0_0_cascade_\
        );

    \I__1748\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16225\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__16225\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_0\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__16222\,
            I => \N__16219\
        );

    \I__1745\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__16216\,
            I => \b2v_inst11.func_state_RNIVS8U1_0Z0Z_0\
        );

    \I__1743\ : InMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__16207\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1\
        );

    \I__1740\ : InMux
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__16201\,
            I => \N__16198\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__16198\,
            I => \b2v_inst11.N_340\
        );

    \I__1737\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16192\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__16192\,
            I => \b2v_inst11.func_state_1_ss0_i_0_o3_1\
        );

    \I__1735\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16184\
        );

    \I__1734\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16179\
        );

    \I__1733\ : InMux
    port map (
            O => \N__16187\,
            I => \N__16179\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__16184\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__16179\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_1\
        );

    \I__1730\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16171\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__16171\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__16168\,
            I => \b2v_inst11.count_off_RNIZ0Z_9_cascade_\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__16165\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_1_cascade_\
        );

    \I__1726\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16159\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__16159\,
            I => \b2v_inst11.un1_func_state25_4_i_a3_0_1\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__16156\,
            I => \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__16153\,
            I => \b2v_inst11.count_clkZ0Z_1_cascade_\
        );

    \I__1722\ : InMux
    port map (
            O => \N__16150\,
            I => \N__16147\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__16147\,
            I => \b2v_inst11.count_clk_0_1\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__16144\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__16141\,
            I => \N__16138\
        );

    \I__1718\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16135\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__16135\,
            I => \N__16131\
        );

    \I__1716\ : InMux
    port map (
            O => \N__16134\,
            I => \N__16128\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__16131\,
            I => \b2v_inst11.count_clk_RNIVS8U1Z0Z_13\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__16128\,
            I => \b2v_inst11.count_clk_RNIVS8U1Z0Z_13\
        );

    \I__1713\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16120\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__16120\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_329_N\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__16117\,
            I => \b2v_inst11.un1_func_state25_6_0_1_cascade_\
        );

    \I__1710\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16110\
        );

    \I__1709\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16107\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__16110\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_0\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__16107\,
            I => \b2v_inst11.func_state_RNI_1Z0Z_0\
        );

    \I__1706\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16099\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__16099\,
            I => \N__16096\
        );

    \I__1704\ : Span4Mux_s1_h
    port map (
            O => \N__16096\,
            I => \N__16093\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__16093\,
            I => \N_236_0\
        );

    \I__1702\ : InMux
    port map (
            O => \N__16090\,
            I => \N__16087\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__16087\,
            I => \b2v_inst11.g1_0_0_1\
        );

    \I__1700\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16081\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__16081\,
            I => \b2v_inst11.un1_func_state25_6_0_o_N_331_N\
        );

    \I__1698\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16075\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__16075\,
            I => \N__16072\
        );

    \I__1696\ : Odrv4
    port map (
            O => \N__16072\,
            I => \b2v_inst11.count_clk_en_1\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__16069\,
            I => \N__16066\
        );

    \I__1694\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__16063\,
            I => \b2v_inst11.N_328\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__16060\,
            I => \b2v_inst16.N_268_cascade_\
        );

    \I__1691\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16046\
        );

    \I__1690\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16046\
        );

    \I__1689\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16046\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__16054\,
            I => \N__16040\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__16053\,
            I => \N__16031\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__16046\,
            I => \N__16020\
        );

    \I__1685\ : InMux
    port map (
            O => \N__16045\,
            I => \N__16009\
        );

    \I__1684\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16009\
        );

    \I__1683\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16009\
        );

    \I__1682\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16009\
        );

    \I__1681\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16009\
        );

    \I__1680\ : InMux
    port map (
            O => \N__16038\,
            I => \N__16004\
        );

    \I__1679\ : InMux
    port map (
            O => \N__16037\,
            I => \N__16004\
        );

    \I__1678\ : InMux
    port map (
            O => \N__16036\,
            I => \N__15999\
        );

    \I__1677\ : InMux
    port map (
            O => \N__16035\,
            I => \N__15999\
        );

    \I__1676\ : InMux
    port map (
            O => \N__16034\,
            I => \N__15992\
        );

    \I__1675\ : InMux
    port map (
            O => \N__16031\,
            I => \N__15992\
        );

    \I__1674\ : InMux
    port map (
            O => \N__16030\,
            I => \N__15992\
        );

    \I__1673\ : InMux
    port map (
            O => \N__16029\,
            I => \N__15985\
        );

    \I__1672\ : InMux
    port map (
            O => \N__16028\,
            I => \N__15985\
        );

    \I__1671\ : InMux
    port map (
            O => \N__16027\,
            I => \N__15985\
        );

    \I__1670\ : InMux
    port map (
            O => \N__16026\,
            I => \N__15977\
        );

    \I__1669\ : InMux
    port map (
            O => \N__16025\,
            I => \N__15977\
        );

    \I__1668\ : InMux
    port map (
            O => \N__16024\,
            I => \N__15970\
        );

    \I__1667\ : InMux
    port map (
            O => \N__16023\,
            I => \N__15970\
        );

    \I__1666\ : Span4Mux_v
    port map (
            O => \N__16020\,
            I => \N__15965\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__16009\,
            I => \N__15965\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__16004\,
            I => \N__15956\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__15999\,
            I => \N__15956\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__15992\,
            I => \N__15956\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__15985\,
            I => \N__15956\
        );

    \I__1660\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15949\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15949\
        );

    \I__1658\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15949\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__15977\,
            I => \N__15946\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15976\,
            I => \N__15941\
        );

    \I__1655\ : InMux
    port map (
            O => \N__15975\,
            I => \N__15941\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__15970\,
            I => \N__15932\
        );

    \I__1653\ : Span4Mux_s2_v
    port map (
            O => \N__15965\,
            I => \N__15932\
        );

    \I__1652\ : Span4Mux_s2_v
    port map (
            O => \N__15956\,
            I => \N__15932\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15932\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__15946\,
            I => \b2v_inst16.N_26\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15941\,
            I => \b2v_inst16.N_26\
        );

    \I__1648\ : Odrv4
    port map (
            O => \N__15932\,
            I => \b2v_inst16.N_26\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__15925\,
            I => \b2v_inst11.un1_func_state25_6_0_a3_0_0_cascade_\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__15922\,
            I => \b2v_inst11.func_state_RNINPGR_2Z0Z_1_cascade_\
        );

    \I__1645\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15916\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__15916\,
            I => \b2v_inst11.g0_20_1\
        );

    \I__1643\ : InMux
    port map (
            O => \N__15913\,
            I => \N__15910\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__15910\,
            I => \b2v_inst11.count_off_0_10\
        );

    \I__1641\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15904\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__15904\,
            I => \b2v_inst16.N_1440\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__15901\,
            I => \b2v_inst16.curr_state_RNI3B692Z0Z_0_cascade_\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__15898\,
            I => \N__15891\
        );

    \I__1637\ : InMux
    port map (
            O => \N__15897\,
            I => \N__15878\
        );

    \I__1636\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15873\
        );

    \I__1635\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15873\
        );

    \I__1634\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15870\
        );

    \I__1633\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15859\
        );

    \I__1632\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15859\
        );

    \I__1631\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15859\
        );

    \I__1630\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15859\
        );

    \I__1629\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15859\
        );

    \I__1628\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15856\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15845\
        );

    \I__1626\ : InMux
    port map (
            O => \N__15884\,
            I => \N__15845\
        );

    \I__1625\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15845\
        );

    \I__1624\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15845\
        );

    \I__1623\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15845\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__15878\,
            I => \N__15838\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__15873\,
            I => \N__15838\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__15870\,
            I => \N__15838\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__15859\,
            I => \b2v_inst16.N_416\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__15856\,
            I => \b2v_inst16.N_416\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__15845\,
            I => \b2v_inst16.N_416\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__15838\,
            I => \b2v_inst16.N_416\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__15829\,
            I => \b2v_inst16.curr_state_7_0_1_cascade_\
        );

    \I__1614\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15823\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__15823\,
            I => \b2v_inst16.curr_state_2_1\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__15820\,
            I => \b2v_inst16.curr_stateZ0Z_1_cascade_\
        );

    \I__1611\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15814\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__15814\,
            I => \b2v_inst16.curr_state_2_0\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__15811\,
            I => \N__15804\
        );

    \I__1608\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15795\
        );

    \I__1607\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15795\
        );

    \I__1606\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15795\
        );

    \I__1605\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15790\
        );

    \I__1604\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15790\
        );

    \I__1603\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15785\
        );

    \I__1602\ : InMux
    port map (
            O => \N__15802\,
            I => \N__15785\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__15795\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__15790\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__15785\,
            I => \b2v_inst16.curr_stateZ0Z_1\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__15778\,
            I => \N__15774\
        );

    \I__1597\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15769\
        );

    \I__1596\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15762\
        );

    \I__1595\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15762\
        );

    \I__1594\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15762\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__15769\,
            I => \b2v_inst16.curr_state_RNI3B692Z0Z_0\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__15762\,
            I => \b2v_inst16.curr_state_RNI3B692Z0Z_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15754\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__15754\,
            I => \b2v_inst16.N_268\
        );

    \I__1589\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15748\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15745\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__15745\,
            I => \b2v_inst16.count_4_i_a3_8_0\
        );

    \I__1586\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15739\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__15739\,
            I => \b2v_inst16.count_4_i_a3_10_0\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__15736\,
            I => \b2v_inst16.count_4_i_a3_7_0_cascade_\
        );

    \I__1583\ : InMux
    port map (
            O => \N__15733\,
            I => \N__15730\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__15730\,
            I => \b2v_inst16.count_4_i_a3_9_0\
        );

    \I__1581\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__1580\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15721\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__15721\,
            I => \N__15718\
        );

    \I__1578\ : Span4Mux_s0_v
    port map (
            O => \N__15718\,
            I => \N__15715\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__15715\,
            I => \b2v_inst16.N_414\
        );

    \I__1576\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15702\
        );

    \I__1575\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15702\
        );

    \I__1574\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15702\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__15709\,
            I => \N__15699\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__15702\,
            I => \N__15695\
        );

    \I__1571\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15692\
        );

    \I__1570\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15689\
        );

    \I__1569\ : Span4Mux_v
    port map (
            O => \N__15695\,
            I => \N__15684\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15684\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__15689\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__15684\,
            I => \b2v_inst16.countZ0Z_0\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__15679\,
            I => \b2v_inst16.N_414_cascade_\
        );

    \I__1564\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15673\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__15673\,
            I => \N__15670\
        );

    \I__1562\ : Odrv12
    port map (
            O => \N__15670\,
            I => \b2v_inst16.count_4_0\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__15667\,
            I => \b2v_inst11.count_offZ0Z_0_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15661\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__15661\,
            I => \b2v_inst11.count_off_RNIZ0Z_1\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__15658\,
            I => \b2v_inst11.count_off_RNIZ0Z_1_cascade_\
        );

    \I__1557\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15652\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__15652\,
            I => \b2v_inst11.count_off_0_1\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \N__15646\
        );

    \I__1554\ : InMux
    port map (
            O => \N__15646\,
            I => \N__15643\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__15643\,
            I => \b2v_inst11.count_off_0_0\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__15640\,
            I => \b2v_inst16.count_rst_9_cascade_\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__15637\,
            I => \N__15634\
        );

    \I__1550\ : InMux
    port map (
            O => \N__15634\,
            I => \N__15627\
        );

    \I__1549\ : InMux
    port map (
            O => \N__15633\,
            I => \N__15627\
        );

    \I__1548\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15624\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__15627\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__15624\,
            I => \b2v_inst16.countZ0Z_4\
        );

    \I__1545\ : InMux
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__1544\ : InMux
    port map (
            O => \N__15618\,
            I => \N__15613\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__15613\,
            I => \b2v_inst16.un4_count_1_cry_3_THRU_CO\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__15610\,
            I => \b2v_inst16.countZ0Z_4_cascade_\
        );

    \I__1541\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15604\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__15604\,
            I => \b2v_inst16.count_4_4\
        );

    \I__1539\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15595\
        );

    \I__1538\ : InMux
    port map (
            O => \N__15600\,
            I => \N__15595\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__15595\,
            I => \b2v_inst16.count_rst_2\
        );

    \I__1536\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15589\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__15589\,
            I => \b2v_inst16.count_4_13\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__15586\,
            I => \b2v_inst16.un4_count_1_axb_1_cascade_\
        );

    \I__1533\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15579\
        );

    \I__1532\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15576\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__15579\,
            I => \b2v_inst16.un4_count_1_axb_1\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__15576\,
            I => \b2v_inst16.un4_count_1_axb_1\
        );

    \I__1529\ : InMux
    port map (
            O => \N__15571\,
            I => \N__15568\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__15568\,
            I => \N__15565\
        );

    \I__1527\ : Span4Mux_s2_h
    port map (
            O => \N__15565\,
            I => \N__15561\
        );

    \I__1526\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15558\
        );

    \I__1525\ : Odrv4
    port map (
            O => \N__15561\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__15558\,
            I => \b2v_inst16.countZ0Z_6\
        );

    \I__1523\ : InMux
    port map (
            O => \N__15553\,
            I => \N__15549\
        );

    \I__1522\ : InMux
    port map (
            O => \N__15552\,
            I => \N__15546\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__15549\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__15546\,
            I => \b2v_inst16.countZ0Z_12\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__15541\,
            I => \N__15537\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__15540\,
            I => \N__15534\
        );

    \I__1517\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15531\
        );

    \I__1516\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15528\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__15531\,
            I => \N__15523\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__15528\,
            I => \N__15523\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__15523\,
            I => \b2v_inst16.countZ0Z_10\
        );

    \I__1512\ : InMux
    port map (
            O => \N__15520\,
            I => \N__15516\
        );

    \I__1511\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15513\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__15516\,
            I => \N__15510\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__15513\,
            I => \N__15507\
        );

    \I__1508\ : Odrv4
    port map (
            O => \N__15510\,
            I => \b2v_inst16.countZ0Z_2\
        );

    \I__1507\ : Odrv12
    port map (
            O => \N__15507\,
            I => \b2v_inst16.countZ0Z_2\
        );

    \I__1506\ : InMux
    port map (
            O => \N__15502\,
            I => \N__15498\
        );

    \I__1505\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15495\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__15498\,
            I => \b2v_inst16.count_4_1\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__15495\,
            I => \b2v_inst16.count_4_1\
        );

    \I__1502\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__1501\ : InMux
    port map (
            O => \N__15489\,
            I => \N__15484\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__15484\,
            I => \b2v_inst16.count_rst_6\
        );

    \I__1499\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15478\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__15478\,
            I => \N__15474\
        );

    \I__1497\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15471\
        );

    \I__1496\ : Span12Mux_s1_h
    port map (
            O => \N__15474\,
            I => \N__15466\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__15471\,
            I => \N__15466\
        );

    \I__1494\ : Odrv12
    port map (
            O => \N__15466\,
            I => \b2v_inst16.countZ0Z_15\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__15463\,
            I => \b2v_inst16.countZ0Z_1_cascade_\
        );

    \I__1492\ : InMux
    port map (
            O => \N__15460\,
            I => \N__15457\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__15457\,
            I => \N__15453\
        );

    \I__1490\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15449\
        );

    \I__1489\ : Span4Mux_v
    port map (
            O => \N__15453\,
            I => \N__15446\
        );

    \I__1488\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15443\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__15449\,
            I => \N__15440\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__15446\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__15443\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1484\ : Odrv12
    port map (
            O => \N__15440\,
            I => \b2v_inst16.countZ0Z_11\
        );

    \I__1483\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15427\
        );

    \I__1482\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15427\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__15427\,
            I => \N__15424\
        );

    \I__1480\ : Span4Mux_s1_v
    port map (
            O => \N__15424\,
            I => \N__15421\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__15421\,
            I => \b2v_inst16.count_rst_4\
        );

    \I__1478\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15415\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__15415\,
            I => \b2v_inst16.count_4_15\
        );

    \I__1476\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__15409\,
            I => \b2v_inst16.count_4_14\
        );

    \I__1474\ : InMux
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__1473\ : InMux
    port map (
            O => \N__15405\,
            I => \N__15400\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__15400\,
            I => \b2v_inst16.count_rst_3\
        );

    \I__1471\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15394\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__15394\,
            I => \b2v_inst16.countZ0Z_14\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__15391\,
            I => \N__15386\
        );

    \I__1468\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15383\
        );

    \I__1467\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15380\
        );

    \I__1466\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15377\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__15383\,
            I => \N__15374\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__15380\,
            I => \N__15371\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__15377\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__15374\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1461\ : Odrv4
    port map (
            O => \N__15371\,
            I => \b2v_inst16.countZ0Z_3\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__15364\,
            I => \b2v_inst16.countZ0Z_14_cascade_\
        );

    \I__1459\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15357\
        );

    \I__1458\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15354\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__15357\,
            I => \b2v_inst16.countZ0Z_13\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__15354\,
            I => \b2v_inst16.countZ0Z_13\
        );

    \I__1455\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15345\
        );

    \I__1454\ : InMux
    port map (
            O => \N__15348\,
            I => \N__15341\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__15345\,
            I => \N__15338\
        );

    \I__1452\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15335\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__15341\,
            I => \N__15332\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__15338\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__15335\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__15332\,
            I => \b2v_inst16.countZ0Z_8\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \b2v_inst16.N_416_cascade_\
        );

    \I__1446\ : InMux
    port map (
            O => \N__15322\,
            I => \N__15318\
        );

    \I__1445\ : InMux
    port map (
            O => \N__15321\,
            I => \N__15315\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__15318\,
            I => \N__15310\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__15315\,
            I => \N__15310\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__15310\,
            I => \b2v_inst16.un4_count_1_cry_7_THRU_CO\
        );

    \I__1441\ : InMux
    port map (
            O => \N__15307\,
            I => \N__15304\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__15304\,
            I => \b2v_inst16.count_rst_13\
        );

    \I__1439\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15298\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__15298\,
            I => \b2v_inst16.count_rst_5\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__15295\,
            I => \N__15291\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__15294\,
            I => \N__15288\
        );

    \I__1435\ : InMux
    port map (
            O => \N__15291\,
            I => \N__15285\
        );

    \I__1434\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15282\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__15285\,
            I => \N__15279\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__15282\,
            I => \b2v_inst16.un4_count_1_cry_4_THRU_CO\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__15279\,
            I => \b2v_inst16.un4_count_1_cry_4_THRU_CO\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__15274\,
            I => \b2v_inst16.count_rst_10_cascade_\
        );

    \I__1429\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15268\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__15268\,
            I => \b2v_inst16.count_4_5\
        );

    \I__1427\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15259\
        );

    \I__1426\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15256\
        );

    \I__1425\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15253\
        );

    \I__1424\ : InMux
    port map (
            O => \N__15262\,
            I => \N__15250\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__15259\,
            I => \N__15247\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__15256\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__15253\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__15250\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__15247\,
            I => \b2v_inst16.countZ0Z_5\
        );

    \I__1418\ : InMux
    port map (
            O => \N__15238\,
            I => \N__15232\
        );

    \I__1417\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15232\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__15232\,
            I => \N__15229\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__15229\,
            I => \b2v_inst16.count_rst\
        );

    \I__1414\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15223\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__15223\,
            I => \b2v_inst16.count_4_10\
        );

    \I__1412\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15214\
        );

    \I__1411\ : InMux
    port map (
            O => \N__15219\,
            I => \N__15214\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__15214\,
            I => \b2v_inst16.count_rst_11\
        );

    \I__1409\ : InMux
    port map (
            O => \N__15211\,
            I => \N__15208\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__15208\,
            I => \b2v_inst16.count_4_6\
        );

    \I__1407\ : InMux
    port map (
            O => \N__15205\,
            I => \bfn_1_16_0_\
        );

    \I__1406\ : InMux
    port map (
            O => \N__15202\,
            I => \b2v_inst20.counter_1_cry_25\
        );

    \I__1405\ : InMux
    port map (
            O => \N__15199\,
            I => \b2v_inst20.counter_1_cry_26\
        );

    \I__1404\ : InMux
    port map (
            O => \N__15196\,
            I => \b2v_inst20.counter_1_cry_27\
        );

    \I__1403\ : InMux
    port map (
            O => \N__15193\,
            I => \b2v_inst20.counter_1_cry_28\
        );

    \I__1402\ : InMux
    port map (
            O => \N__15190\,
            I => \b2v_inst20.counter_1_cry_29\
        );

    \I__1401\ : InMux
    port map (
            O => \N__15187\,
            I => \b2v_inst20.counter_1_cry_30\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__15184\,
            I => \b2v_inst16.countZ0Z_0_cascade_\
        );

    \I__1399\ : InMux
    port map (
            O => \N__15181\,
            I => \b2v_inst20.counter_1_cry_15\
        );

    \I__1398\ : InMux
    port map (
            O => \N__15178\,
            I => \bfn_1_15_0_\
        );

    \I__1397\ : InMux
    port map (
            O => \N__15175\,
            I => \b2v_inst20.counter_1_cry_17\
        );

    \I__1396\ : InMux
    port map (
            O => \N__15172\,
            I => \b2v_inst20.counter_1_cry_18\
        );

    \I__1395\ : InMux
    port map (
            O => \N__15169\,
            I => \b2v_inst20.counter_1_cry_19\
        );

    \I__1394\ : InMux
    port map (
            O => \N__15166\,
            I => \b2v_inst20.counter_1_cry_20\
        );

    \I__1393\ : InMux
    port map (
            O => \N__15163\,
            I => \b2v_inst20.counter_1_cry_21\
        );

    \I__1392\ : InMux
    port map (
            O => \N__15160\,
            I => \b2v_inst20.counter_1_cry_22\
        );

    \I__1391\ : InMux
    port map (
            O => \N__15157\,
            I => \b2v_inst20.counter_1_cry_23\
        );

    \I__1390\ : InMux
    port map (
            O => \N__15154\,
            I => \b2v_inst20.counter_1_cry_6\
        );

    \I__1389\ : InMux
    port map (
            O => \N__15151\,
            I => \b2v_inst20.counter_1_cry_7\
        );

    \I__1388\ : InMux
    port map (
            O => \N__15148\,
            I => \bfn_1_14_0_\
        );

    \I__1387\ : InMux
    port map (
            O => \N__15145\,
            I => \b2v_inst20.counter_1_cry_9\
        );

    \I__1386\ : InMux
    port map (
            O => \N__15142\,
            I => \b2v_inst20.counter_1_cry_10\
        );

    \I__1385\ : InMux
    port map (
            O => \N__15139\,
            I => \b2v_inst20.counter_1_cry_11\
        );

    \I__1384\ : InMux
    port map (
            O => \N__15136\,
            I => \b2v_inst20.counter_1_cry_12\
        );

    \I__1383\ : InMux
    port map (
            O => \N__15133\,
            I => \b2v_inst20.counter_1_cry_13\
        );

    \I__1382\ : InMux
    port map (
            O => \N__15130\,
            I => \b2v_inst20.counter_1_cry_14\
        );

    \I__1381\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15123\
        );

    \I__1380\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15120\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__15123\,
            I => \N__15115\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__15120\,
            I => \N__15115\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__15115\,
            I => \b2v_inst11.un2_count_clk_17_0_o2_4\
        );

    \I__1376\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15109\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__15109\,
            I => \b2v_inst11.count_clk_0_11\
        );

    \I__1374\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15103\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__15100\,
            I => \b2v_inst11.count_clk_0_4\
        );

    \I__1371\ : InMux
    port map (
            O => \N__15097\,
            I => \b2v_inst20.counter_1_cry_1\
        );

    \I__1370\ : InMux
    port map (
            O => \N__15094\,
            I => \b2v_inst20.counter_1_cry_2\
        );

    \I__1369\ : InMux
    port map (
            O => \N__15091\,
            I => \b2v_inst20.counter_1_cry_3\
        );

    \I__1368\ : InMux
    port map (
            O => \N__15088\,
            I => \b2v_inst20.counter_1_cry_4\
        );

    \I__1367\ : InMux
    port map (
            O => \N__15085\,
            I => \b2v_inst20.counter_1_cry_5\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__15082\,
            I => \b2v_inst11.count_clk_en_cascade_\
        );

    \I__1365\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15076\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__15076\,
            I => \b2v_inst11.count_clk_0_13\
        );

    \I__1363\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15070\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__15070\,
            I => \b2v_inst11.count_clk_0_15\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__15067\,
            I => \N__15064\
        );

    \I__1360\ : InMux
    port map (
            O => \N__15064\,
            I => \N__15061\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__15061\,
            I => \b2v_inst11.count_clk_0_12\
        );

    \I__1358\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15055\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__15055\,
            I => \b2v_inst11.count_clk_0_10\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__15052\,
            I => \b2v_inst11.count_clkZ0Z_10_cascade_\
        );

    \I__1355\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15046\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__15046\,
            I => \N__15043\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__15043\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2\
        );

    \I__1352\ : InMux
    port map (
            O => \N__15040\,
            I => \N__15037\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__15037\,
            I => \b2v_inst11.count_clk_RNIVS8U1Z0Z_14\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__15034\,
            I => \N__15031\
        );

    \I__1349\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15028\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__15028\,
            I => \b2v_inst11.N_428\
        );

    \I__1347\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15022\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__15022\,
            I => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__15019\,
            I => \N__15016\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__15016\,
            I => \b2v_inst11.N_175\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__15013\,
            I => \b2v_inst11.N_175_cascade_\
        );

    \I__1342\ : InMux
    port map (
            O => \N__15010\,
            I => \N__15007\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__15007\,
            I => \b2v_inst11.N_190\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__15004\,
            I => \b2v_inst11.N_190_cascade_\
        );

    \I__1339\ : InMux
    port map (
            O => \N__15001\,
            I => \N__14998\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__14998\,
            I => \b2v_inst11.un2_count_clk_17_0_o3_0_4\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__14995\,
            I => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__14992\,
            I => \b2v_inst11.N_379_cascade_\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__14989\,
            I => \N__14986\
        );

    \I__1334\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14983\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__14983\,
            I => \SLP_S3n_ibuf_RNIF6NLZ0\
        );

    \I__1332\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14974\
        );

    \I__1331\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14974\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__14974\,
            I => \N__14971\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__14971\,
            I => \b2v_inst11.N_379\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__14968\,
            I => \N__14965\
        );

    \I__1327\ : InMux
    port map (
            O => \N__14965\,
            I => \N__14962\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__14962\,
            I => \b2v_inst11.count_clk_RNI_0Z0Z_13\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__14959\,
            I => \b2v_inst11.g3_cascade_\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__14956\,
            I => \b2v_inst11.g1_0_1_cascade_\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__14953\,
            I => \b2v_inst11.N_7_3_0_cascade_\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__14950\,
            I => \b2v_inst11.g2_1_0_0_cascade_\
        );

    \I__1321\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14944\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__14944\,
            I => \b2v_inst11.g2_2_0\
        );

    \I__1319\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14938\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__14938\,
            I => \N__14935\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__14935\,
            I => \N__14932\
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__14932\,
            I => \b2v_inst11.g2_1_0\
        );

    \I__1315\ : InMux
    port map (
            O => \N__14929\,
            I => \N__14926\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__14926\,
            I => \b2v_inst11.g0_12_0\
        );

    \I__1313\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14920\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__14920\,
            I => \b2v_inst16.delayed_vddq_pwrgd_en\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__14917\,
            I => \N__14913\
        );

    \I__1310\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14908\
        );

    \I__1309\ : InMux
    port map (
            O => \N__14913\,
            I => \N__14908\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__14908\,
            I => \b2v_inst16.delayed_vddq_pwrgdZ0\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__14905\,
            I => \b2v_inst16.delayed_vddq_pwrgd_en_cascade_\
        );

    \I__1306\ : IoInMux
    port map (
            O => \N__14902\,
            I => \N__14899\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__14899\,
            I => \N__14896\
        );

    \I__1304\ : IoSpan4Mux
    port map (
            O => \N__14896\,
            I => \N__14893\
        );

    \I__1303\ : IoSpan4Mux
    port map (
            O => \N__14893\,
            I => \N__14890\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__14890\,
            I => b2v_inst16_un2_vpp_en_0_i
        );

    \I__1301\ : IoInMux
    port map (
            O => \N__14887\,
            I => \N__14884\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__14884\,
            I => \N__14881\
        );

    \I__1299\ : Span4Mux_s0_h
    port map (
            O => \N__14881\,
            I => \N__14878\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__14878\,
            I => \b2v_inst200.count_enZ0\
        );

    \I__1297\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14871\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14868\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__14871\,
            I => \N__14865\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__14868\,
            I => \N__14862\
        );

    \I__1293\ : Odrv12
    port map (
            O => \N__14865\,
            I => \b2v_inst16.count_rst_7\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__14862\,
            I => \b2v_inst16.count_rst_7\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__14857\,
            I => \b2v_inst16.count_en_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14851\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__14851\,
            I => \b2v_inst16.count_4_2\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__14848\,
            I => \N__14845\
        );

    \I__1287\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14838\
        );

    \I__1286\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14838\
        );

    \I__1285\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14835\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__14838\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__14835\,
            I => \b2v_inst16.countZ0Z_7\
        );

    \I__1282\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14824\
        );

    \I__1281\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14824\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__14824\,
            I => \b2v_inst16.un4_count_1_cry_6_THRU_CO\
        );

    \I__1279\ : InMux
    port map (
            O => \N__14821\,
            I => \b2v_inst16.un4_count_1_cry_6\
        );

    \I__1278\ : InMux
    port map (
            O => \N__14818\,
            I => \b2v_inst16.un4_count_1_cry_7\
        );

    \I__1277\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14810\
        );

    \I__1276\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14805\
        );

    \I__1275\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14805\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__14810\,
            I => \N__14802\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__14805\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__14802\,
            I => \b2v_inst16.countZ0Z_9\
        );

    \I__1271\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14791\
        );

    \I__1270\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14791\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__14791\,
            I => \N__14788\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__14788\,
            I => \b2v_inst16.un4_count_1_cry_8_THRU_CO\
        );

    \I__1267\ : InMux
    port map (
            O => \N__14785\,
            I => \bfn_1_4_0_\
        );

    \I__1266\ : InMux
    port map (
            O => \N__14782\,
            I => \b2v_inst16.un4_count_1_cry_9\
        );

    \I__1265\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14773\
        );

    \I__1264\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14773\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__14773\,
            I => \N__14770\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__14770\,
            I => \b2v_inst16.un4_count_1_cry_10_THRU_CO\
        );

    \I__1261\ : InMux
    port map (
            O => \N__14767\,
            I => \b2v_inst16.un4_count_1_cry_10\
        );

    \I__1260\ : InMux
    port map (
            O => \N__14764\,
            I => \b2v_inst16.un4_count_1_cry_11\
        );

    \I__1259\ : InMux
    port map (
            O => \N__14761\,
            I => \b2v_inst16.un4_count_1_cry_12\
        );

    \I__1258\ : InMux
    port map (
            O => \N__14758\,
            I => \b2v_inst16.un4_count_1_cry_13\
        );

    \I__1257\ : InMux
    port map (
            O => \N__14755\,
            I => \b2v_inst16.un4_count_1_cry_14\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__14752\,
            I => \b2v_inst16.count_rst_12_cascade_\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__14749\,
            I => \b2v_inst16.countZ0Z_7_cascade_\
        );

    \I__1254\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14743\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__14743\,
            I => \b2v_inst16.count_4_7\
        );

    \I__1252\ : InMux
    port map (
            O => \N__14740\,
            I => \b2v_inst16.un4_count_1_cry_1\
        );

    \I__1251\ : InMux
    port map (
            O => \N__14737\,
            I => \N__14731\
        );

    \I__1250\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14731\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__14731\,
            I => \N__14728\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__14728\,
            I => \b2v_inst16.un4_count_1_cry_2_THRU_CO\
        );

    \I__1247\ : InMux
    port map (
            O => \N__14725\,
            I => \b2v_inst16.un4_count_1_cry_2\
        );

    \I__1246\ : InMux
    port map (
            O => \N__14722\,
            I => \b2v_inst16.un4_count_1_cry_3\
        );

    \I__1245\ : InMux
    port map (
            O => \N__14719\,
            I => \b2v_inst16.un4_count_1_cry_4\
        );

    \I__1244\ : InMux
    port map (
            O => \N__14716\,
            I => \b2v_inst16.un4_count_1_cry_5\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__14713\,
            I => \b2v_inst16.countZ0Z_8_cascade_\
        );

    \I__1242\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14707\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__14707\,
            I => \b2v_inst16.count_4_8\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__14704\,
            I => \b2v_inst16.count_rst_8_cascade_\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__14701\,
            I => \b2v_inst16.countZ0Z_3_cascade_\
        );

    \I__1238\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__14695\,
            I => \b2v_inst16.count_4_3\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__14692\,
            I => \b2v_inst16.countZ0Z_9_cascade_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14686\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__14686\,
            I => \b2v_inst16.count_rst_14\
        );

    \I__1233\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14680\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__14680\,
            I => \b2v_inst16.count_4_9\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__14677\,
            I => \b2v_inst16.count_rst_0_cascade_\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__14674\,
            I => \b2v_inst16.countZ0Z_11_cascade_\
        );

    \I__1229\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14668\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__14668\,
            I => \b2v_inst16.count_4_11\
        );

    \IN_MUX_bfv_12_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_1_0_\
        );

    \IN_MUX_bfv_12_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst6.un2_count_1_cry_8\,
            carryinitout => \bfn_12_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst5.un2_count_1_cry_8\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst36.un2_count_1_cry_8\,
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_2_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_15_0_\
        );

    \IN_MUX_bfv_2_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => b2v_inst20_un4_counter_7,
            carryinitout => \bfn_2_16_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_8\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_16\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst20.counter_1_cry_24\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst16.un4_count_1_cry_8\,
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_4_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_4_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un3_count_off_1_cry_8\,
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_cry_8\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_count_clk_2_cry_8\,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_5_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_1_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_7\,
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst200.un2_count_1_cry_15\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_7\,
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \b2v_inst11.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \b2v_inst200.count_en_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14887\,
            GLOBALBUFFEROUTPUT => \b2v_inst200.count_en_g\
        );

    \N_606_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__27603\,
            GLOBALBUFFEROUTPUT => \N_606_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__15882\,
            in1 => \N__14778\,
            in2 => \N__16053\,
            in3 => \N__15452\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIDGU31_11_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20937\,
            in1 => \_gnd_net_\,
            in2 => \N__14677\,
            in3 => \N__14671\,
            lcout => \b2v_inst16.countZ0Z_11\,
            ltout => \b2v_inst16.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_11_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__15883\,
            in1 => \N__16037\,
            in2 => \N__14674\,
            in3 => \N__14779\,
            lcout => \b2v_inst16.count_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36609\,
            ce => \N__20949\,
            sr => \N__20799\
        );

    \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20936\,
            in1 => \N__14710\,
            in2 => \_gnd_net_\,
            in3 => \N__15307\,
            lcout => \b2v_inst16.countZ0Z_8\,
            ltout => \b2v_inst16.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_8_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__15884\,
            in1 => \N__16038\,
            in2 => \N__14713\,
            in3 => \N__15322\,
            lcout => \b2v_inst16.count_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36609\,
            ce => \N__20949\,
            sr => \N__20799\
        );

    \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__14736\,
            in1 => \N__16030\,
            in2 => \N__15391\,
            in3 => \N__15881\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14698\,
            in2 => \N__14704\,
            in3 => \N__20935\,
            lcout => \b2v_inst16.countZ0Z_3\,
            ltout => \b2v_inst16.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_3_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__14737\,
            in1 => \N__16034\,
            in2 => \N__14701\,
            in3 => \N__15885\,
            lcout => \b2v_inst16.count_4_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36609\,
            ce => \N__20949\,
            sr => \N__20799\
        );

    \b2v_inst16.count_RNIRP4K1_9_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20941\,
            in1 => \N__14683\,
            in2 => \_gnd_net_\,
            in3 => \N__14689\,
            lcout => \b2v_inst16.countZ0Z_9\,
            ltout => \b2v_inst16.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_5_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15262\,
            in1 => \N__14844\,
            in2 => \N__14692\,
            in3 => \N__15344\,
            lcout => \b2v_inst16.count_4_i_a3_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000100000"
        )
    port map (
            in0 => \N__14814\,
            in1 => \N__15888\,
            in2 => \N__16054\,
            in3 => \N__14796\,
            lcout => \b2v_inst16.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_9_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__14797\,
            in1 => \N__16044\,
            in2 => \N__15898\,
            in3 => \N__14813\,
            lcout => \b2v_inst16.count_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36601\,
            ce => \N__20928\,
            sr => \N__20785\
        );

    \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__16039\,
            in1 => \N__15887\,
            in2 => \N__14848\,
            in3 => \N__14829\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNINJ2K1_7_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14746\,
            in2 => \N__14752\,
            in3 => \N__20940\,
            lcout => \b2v_inst16.countZ0Z_7\,
            ltout => \b2v_inst16.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_7_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__16043\,
            in1 => \N__15890\,
            in2 => \N__14749\,
            in3 => \N__14830\,
            lcout => \b2v_inst16.count_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36601\,
            ce => \N__20928\,
            sr => \N__20785\
        );

    \b2v_inst16.count_5_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__15889\,
            in1 => \N__15263\,
            in2 => \N__15294\,
            in3 => \N__16045\,
            lcout => \b2v_inst16.count_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36601\,
            ce => \N__20928\,
            sr => \N__20785\
        );

    \b2v_inst16.un4_count_1_cry_1_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15582\,
            in2 => \N__15709\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16036\,
            in1 => \N__15519\,
            in2 => \_gnd_net_\,
            in3 => \N__14740\,
            lcout => \b2v_inst16.count_rst_7\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_1\,
            carryout => \b2v_inst16.un4_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15389\,
            in2 => \_gnd_net_\,
            in3 => \N__14725\,
            lcout => \b2v_inst16.un4_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_2\,
            carryout => \b2v_inst16.un4_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15632\,
            in2 => \_gnd_net_\,
            in3 => \N__14722\,
            lcout => \b2v_inst16.un4_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_3\,
            carryout => \b2v_inst16.un4_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15265\,
            in2 => \_gnd_net_\,
            in3 => \N__14719\,
            lcout => \b2v_inst16.un4_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_4\,
            carryout => \b2v_inst16.un4_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16035\,
            in1 => \N__15564\,
            in2 => \_gnd_net_\,
            in3 => \N__14716\,
            lcout => \b2v_inst16.count_rst_11\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_5\,
            carryout => \b2v_inst16.un4_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14843\,
            in2 => \_gnd_net_\,
            in3 => \N__14821\,
            lcout => \b2v_inst16.un4_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_6\,
            carryout => \b2v_inst16.un4_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15348\,
            in2 => \_gnd_net_\,
            in3 => \N__14818\,
            lcout => \b2v_inst16.un4_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_7\,
            carryout => \b2v_inst16.un4_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14815\,
            in2 => \_gnd_net_\,
            in3 => \N__14785\,
            lcout => \b2v_inst16.un4_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => \b2v_inst16.un4_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16055\,
            in1 => \_gnd_net_\,
            in2 => \N__15540\,
            in3 => \N__14782\,
            lcout => \b2v_inst16.count_rst\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_9\,
            carryout => \b2v_inst16.un4_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15456\,
            in2 => \_gnd_net_\,
            in3 => \N__14767\,
            lcout => \b2v_inst16.un4_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_10\,
            carryout => \b2v_inst16.un4_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_11_c_RNIFJV31_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16056\,
            in1 => \N__15552\,
            in2 => \_gnd_net_\,
            in3 => \N__14764\,
            lcout => \b2v_inst16.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_11\,
            carryout => \b2v_inst16.un4_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16023\,
            in1 => \N__15360\,
            in2 => \_gnd_net_\,
            in3 => \N__14761\,
            lcout => \b2v_inst16.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_12\,
            carryout => \b2v_inst16.un4_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16057\,
            in1 => \N__15397\,
            in2 => \_gnd_net_\,
            in3 => \N__14758\,
            lcout => \b2v_inst16.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst16.un4_count_1_cry_13\,
            carryout => \b2v_inst16.un4_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16024\,
            in1 => \N__15481\,
            in2 => \_gnd_net_\,
            in3 => \N__14755\,
            lcout => \b2v_inst16.count_rst_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIKN901_12_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20962\,
            in1 => \N__20913\,
            in2 => \_gnd_net_\,
            in3 => \N__20973\,
            lcout => \b2v_inst16.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_2_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14874\,
            lcout => \b2v_inst16.count_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36588\,
            ce => \N__20943\,
            sr => \N__20763\
        );

    \b2v_inst16.delayed_vddq_pwrgd_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__15803\,
            in1 => \N__14923\,
            in2 => \N__14917\,
            in3 => \N__15777\,
            lcout => \b2v_inst16.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36585\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI2ABP4_0_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15757\,
            in2 => \_gnd_net_\,
            in3 => \N__36406\,
            lcout => \b2v_inst16.delayed_vddq_pwrgd_en\,
            ltout => \b2v_inst16.delayed_vddq_pwrgd_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.delayed_vddq_pwrgd_RNI8SES8_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100111011"
        )
    port map (
            in0 => \N__14916\,
            in1 => \N__21202\,
            in2 => \N__14905\,
            in3 => \N__15907\,
            lcout => b2v_inst16_un2_vpp_en_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_en_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36404\,
            in2 => \_gnd_net_\,
            in3 => \N__22623\,
            lcout => \b2v_inst200.count_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GPIO_FPGA_SoC_4_ibuf_RNINPGR_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__24390\,
            in1 => \N__24643\,
            in2 => \N__24148\,
            in3 => \N__16102\,
            lcout => \N_15_i_0_a4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIKEBL_1_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__15975\,
            in1 => \N__15802\,
            in2 => \_gnd_net_\,
            in3 => \N__36405\,
            lcout => \b2v_inst16.count_en\,
            ltout => \b2v_inst16.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNID4TJ1_2_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__14875\,
            in1 => \_gnd_net_\,
            in2 => \N__14857\,
            in3 => \N__14854\,
            lcout => \b2v_inst16.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI_0_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.N_2987_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI863D_6_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24162\,
            in2 => \_gnd_net_\,
            in3 => \N__26612\,
            lcout => OPEN,
            ltout => \b2v_inst11.g3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIDGAL3_0_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011111111"
        )
    port map (
            in0 => \N__24389\,
            in1 => \N__16090\,
            in2 => \N__14959\,
            in3 => \N__23904\,
            lcout => OPEN,
            ltout => \b2v_inst11.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI24DD8_7_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101010101"
        )
    port map (
            in0 => \N__14947\,
            in1 => \N__26789\,
            in2 => \N__14956\,
            in3 => \N__25859\,
            lcout => \b2v_inst11.dutycycle_RNI24DD8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIF6NL_7_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__26790\,
            in1 => \N__23722\,
            in2 => \N__24166\,
            in3 => \N__14929\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_7_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI608H1_7_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__14941\,
            in1 => \N__23164\,
            in2 => \N__14953\,
            in3 => \N__26611\,
            lcout => OPEN,
            ltout => \b2v_inst11.g2_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIMMPP2_7_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__23165\,
            in1 => \N__26791\,
            in2 => \N__14950\,
            in3 => \N__23903\,
            lcout => \b2v_inst11.g2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNINPGR_7_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15919\,
            in1 => \N__24642\,
            in2 => \N__26831\,
            in3 => \N__23166\,
            lcout => \b2v_inst11.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI70K8_0_0_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__23182\,
            in1 => \N__24387\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.g0_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S3n_ibuf_RNI9HQH3_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100110011"
        )
    port map (
            in0 => \N__23880\,
            in1 => \N__33782\,
            in2 => \N__14989\,
            in3 => \N__17590\,
            lcout => \SLP_S3n_ibuf_RNI9HQHZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_4_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__16287\,
            in1 => \N__17875\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_2_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18430\,
            in1 => \N__18361\,
            in2 => \N__14995\,
            in3 => \N__17904\,
            lcout => \b2v_inst11.N_379\,
            ltout => \b2v_inst11.N_379_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_1_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16374\,
            in1 => \N__15049\,
            in2 => \N__14992\,
            in3 => \N__15019\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_7_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14980\,
            in1 => \N__15010\,
            in2 => \_gnd_net_\,
            in3 => \N__16572\,
            lcout => \b2v_inst11.N_428\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_2_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__16286\,
            in1 => \N__17903\,
            in2 => \N__18429\,
            in3 => \N__18356\,
            lcout => \b2v_inst11.un2_count_clk_17_0_o3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S3n_ibuf_RNIF6NL_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__30295\,
            in1 => \N__24388\,
            in2 => \_gnd_net_\,
            in3 => \N__24127\,
            lcout => \SLP_S3n_ibuf_RNIF6NLZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVS8U1_13_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15040\,
            in1 => \N__14979\,
            in2 => \N__14968\,
            in3 => \N__15127\,
            lcout => \b2v_inst11.count_clk_RNIVS8U1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINPGR_1_1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__24511\,
            in1 => \N__24212\,
            in2 => \N__26641\,
            in3 => \N__16174\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_13_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16567\,
            in1 => \N__16369\,
            in2 => \N__18322\,
            in3 => \N__16445\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_5_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18259\,
            in1 => \N__18320\,
            in2 => \_gnd_net_\,
            in3 => \N__16568\,
            lcout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI3BJF_4_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__16886\,
            in1 => \N__16273\,
            in2 => \N__18084\,
            in3 => \N__15106\,
            lcout => \b2v_inst11.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVS8U1_14_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__18258\,
            in1 => \N__16407\,
            in2 => \N__16222\,
            in3 => \N__16341\,
            lcout => \b2v_inst11.count_clk_RNIVS8U1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI608H1_1_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__24512\,
            in1 => \N__23698\,
            in2 => \N__15034\,
            in3 => \N__15025\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_13_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16330\,
            in1 => \N__16406\,
            in2 => \N__16449\,
            in3 => \N__15126\,
            lcout => \b2v_inst11.N_175\,
            ltout => \b2v_inst11.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__16368\,
            in1 => \N__18257\,
            in2 => \N__15013\,
            in3 => \N__18316\,
            lcout => \b2v_inst11.N_190\,
            ltout => \b2v_inst11.N_190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_6_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__16566\,
            in1 => \N__17870\,
            in2 => \N__15004\,
            in3 => \N__15001\,
            lcout => \b2v_inst11.N_3038_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_14_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16927\,
            lcout => \b2v_inst11.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__18082\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIMATB8_0_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__17959\,
            in1 => \N__25858\,
            in2 => \N__23179\,
            in3 => \N__16078\,
            lcout => \b2v_inst11.count_clk_en\,
            ltout => \b2v_inst11.count_clk_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI3T3F_13_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16429\,
            in1 => \_gnd_net_\,
            in2 => \N__15082\,
            in3 => \N__15079\,
            lcout => \b2v_inst11.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_13_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16428\,
            lcout => \b2v_inst11.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__18082\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_15_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16794\,
            lcout => \b2v_inst11.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__18082\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI736F_15_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__18083\,
            in1 => \_gnd_net_\,
            in2 => \N__16795\,
            in3 => \N__15073\,
            lcout => \b2v_inst11.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_2_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18384\,
            lcout => \b2v_inst11.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36582\,
            ce => \N__18082\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI1Q2F_12_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__16865\,
            in1 => \N__18054\,
            in2 => \N__15067\,
            in3 => \N__16462\,
            lcout => \b2v_inst11.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_12_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16461\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16870\,
            lcout => \b2v_inst11.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36584\,
            ce => \N__18107\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_10_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16512\,
            lcout => \b2v_inst11.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36584\,
            ce => \N__18107\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIMAMA_10_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__18055\,
            in1 => \N__15058\,
            in2 => \N__16516\,
            in3 => \N__16866\,
            lcout => \b2v_inst11.count_clkZ0Z_10\,
            ltout => \b2v_inst11.count_clkZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_15_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16501\,
            in1 => \N__16474\,
            in2 => \N__15052\,
            in3 => \N__16899\,
            lcout => \b2v_inst11.un2_count_clk_17_0_o2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVM1F_11_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__18056\,
            in1 => \N__15112\,
            in2 => \N__16489\,
            in3 => \N__16867\,
            lcout => \b2v_inst11.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_11_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16485\,
            lcout => \b2v_inst11.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36584\,
            ce => \N__18107\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_4_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16266\,
            in2 => \_gnd_net_\,
            in3 => \N__16871\,
            lcout => \b2v_inst11.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36584\,
            ce => \N__18107\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20326\,
            in2 => \N__18748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \b2v_inst20.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18595\,
            in2 => \_gnd_net_\,
            in3 => \N__15097\,
            lcout => \b2v_inst20.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_1\,
            carryout => \b2v_inst20.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18454\,
            in2 => \_gnd_net_\,
            in3 => \N__15094\,
            lcout => \b2v_inst20.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_2\,
            carryout => \b2v_inst20.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18676\,
            in2 => \_gnd_net_\,
            in3 => \N__15091\,
            lcout => \b2v_inst20.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_3\,
            carryout => \b2v_inst20.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20374\,
            in2 => \_gnd_net_\,
            in3 => \N__15088\,
            lcout => \b2v_inst20.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_4\,
            carryout => \b2v_inst20.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20350\,
            in2 => \_gnd_net_\,
            in3 => \N__15085\,
            lcout => \b2v_inst20.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_5\,
            carryout => \b2v_inst20.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_7_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20388\,
            in2 => \_gnd_net_\,
            in3 => \N__15154\,
            lcout => \b2v_inst20.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_6\,
            carryout => \b2v_inst20.counter_1_cry_7\,
            clk => \N__36587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_8_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16741\,
            in2 => \_gnd_net_\,
            in3 => \N__15151\,
            lcout => \b2v_inst20.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_7\,
            carryout => \b2v_inst20.counter_1_cry_8\,
            clk => \N__36587\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_9_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16768\,
            in2 => \_gnd_net_\,
            in3 => \N__15148\,
            lcout => \b2v_inst20.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \b2v_inst20.counter_1_cry_9\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_10_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16755\,
            in2 => \_gnd_net_\,
            in3 => \N__15145\,
            lcout => \b2v_inst20.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_9\,
            carryout => \b2v_inst20.counter_1_cry_10\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_11_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16780\,
            in2 => \_gnd_net_\,
            in3 => \N__15142\,
            lcout => \b2v_inst20.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_10\,
            carryout => \b2v_inst20.counter_1_cry_11\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_12_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16690\,
            in2 => \_gnd_net_\,
            in3 => \N__15139\,
            lcout => \b2v_inst20.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_11\,
            carryout => \b2v_inst20.counter_1_cry_12\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_13_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16704\,
            in2 => \_gnd_net_\,
            in3 => \N__15136\,
            lcout => \b2v_inst20.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_12\,
            carryout => \b2v_inst20.counter_1_cry_13\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_14_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16717\,
            in2 => \_gnd_net_\,
            in3 => \N__15133\,
            lcout => \b2v_inst20.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_13\,
            carryout => \b2v_inst20.counter_1_cry_14\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_15_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16729\,
            in2 => \_gnd_net_\,
            in3 => \N__15130\,
            lcout => \b2v_inst20.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_14\,
            carryout => \b2v_inst20.counter_1_cry_15\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_16_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16639\,
            in2 => \_gnd_net_\,
            in3 => \N__15181\,
            lcout => \b2v_inst20.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_15\,
            carryout => \b2v_inst20.counter_1_cry_16\,
            clk => \N__36590\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_17_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16666\,
            in2 => \_gnd_net_\,
            in3 => \N__15178\,
            lcout => \b2v_inst20.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \b2v_inst20.counter_1_cry_17\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_18_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16653\,
            in2 => \_gnd_net_\,
            in3 => \N__15175\,
            lcout => \b2v_inst20.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_17\,
            carryout => \b2v_inst20.counter_1_cry_18\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_19_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16678\,
            in2 => \_gnd_net_\,
            in3 => \N__15172\,
            lcout => \b2v_inst20.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_18\,
            carryout => \b2v_inst20.counter_1_cry_19\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_20_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16588\,
            in2 => \_gnd_net_\,
            in3 => \N__15169\,
            lcout => \b2v_inst20.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_19\,
            carryout => \b2v_inst20.counter_1_cry_20\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_21_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16615\,
            in2 => \_gnd_net_\,
            in3 => \N__15166\,
            lcout => \b2v_inst20.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_20\,
            carryout => \b2v_inst20.counter_1_cry_21\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_22_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16602\,
            in2 => \_gnd_net_\,
            in3 => \N__15163\,
            lcout => \b2v_inst20.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_21\,
            carryout => \b2v_inst20.counter_1_cry_22\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_23_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16627\,
            in2 => \_gnd_net_\,
            in3 => \N__15160\,
            lcout => \b2v_inst20.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_22\,
            carryout => \b2v_inst20.counter_1_cry_23\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_24_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17011\,
            in2 => \_gnd_net_\,
            in3 => \N__15157\,
            lcout => \b2v_inst20.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_23\,
            carryout => \b2v_inst20.counter_1_cry_24\,
            clk => \N__36596\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_25_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17038\,
            in2 => \_gnd_net_\,
            in3 => \N__15205\,
            lcout => \b2v_inst20.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \b2v_inst20.counter_1_cry_25\,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_26_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17025\,
            in2 => \_gnd_net_\,
            in3 => \N__15202\,
            lcout => \b2v_inst20.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_25\,
            carryout => \b2v_inst20.counter_1_cry_26\,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_27_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17050\,
            in2 => \_gnd_net_\,
            in3 => \N__15199\,
            lcout => \b2v_inst20.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_26\,
            carryout => \b2v_inst20.counter_1_cry_27\,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_28_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17068\,
            in2 => \_gnd_net_\,
            in3 => \N__15196\,
            lcout => \b2v_inst20.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_27\,
            carryout => \b2v_inst20.counter_1_cry_28\,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_29_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17095\,
            in2 => \_gnd_net_\,
            in3 => \N__15193\,
            lcout => \b2v_inst20.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_28\,
            carryout => \b2v_inst20.counter_1_cry_29\,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_30_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17082\,
            in2 => \_gnd_net_\,
            in3 => \N__15190\,
            lcout => \b2v_inst20.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \b2v_inst20.counter_1_cry_29\,
            carryout => \b2v_inst20.counter_1_cry_30\,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_31_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17107\,
            in2 => \_gnd_net_\,
            in3 => \N__15187\,
            lcout => \b2v_inst20.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI1I651_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15676\,
            in1 => \N__20932\,
            in2 => \_gnd_net_\,
            in3 => \N__15301\,
            lcout => \b2v_inst16.countZ0Z_0\,
            ltout => \b2v_inst16.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_0_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15184\,
            in3 => \N__15727\,
            lcout => \b2v_inst16.N_416\,
            ltout => \b2v_inst16.N_416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001000"
        )
    port map (
            in0 => \N__16029\,
            in1 => \N__15349\,
            in2 => \N__15325\,
            in3 => \N__15321\,
            lcout => \b2v_inst16.count_rst_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_0_0_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__15698\,
            in1 => \N__16027\,
            in2 => \_gnd_net_\,
            in3 => \N__15726\,
            lcout => \b2v_inst16.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__16028\,
            in1 => \N__15264\,
            in2 => \N__15295\,
            in3 => \N__15886\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__20933\,
            in1 => \_gnd_net_\,
            in2 => \N__15274\,
            in3 => \N__15271\,
            lcout => \b2v_inst16.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI4M8F1_10_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15226\,
            in1 => \N__20934\,
            in2 => \_gnd_net_\,
            in3 => \N__15237\,
            lcout => \b2v_inst16.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_10_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15238\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36615\,
            ce => \N__20942\,
            sr => \N__20798\
        );

    \b2v_inst16.count_RNILG1K1_6_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15211\,
            in1 => \N__15219\,
            in2 => \_gnd_net_\,
            in3 => \N__20938\,
            lcout => \b2v_inst16.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_6_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15220\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36610\,
            ce => \N__20945\,
            sr => \N__20797\
        );

    \b2v_inst16.count_RNILS241_15_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15433\,
            in1 => \N__15418\,
            in2 => \_gnd_net_\,
            in3 => \N__20939\,
            lcout => \b2v_inst16.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_15_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15432\,
            lcout => \b2v_inst16.count_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36610\,
            ce => \N__20945\,
            sr => \N__20797\
        );

    \b2v_inst200.count_RNI3TN71_12_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25212\,
            in1 => \N__17143\,
            in2 => \_gnd_net_\,
            in3 => \N__18904\,
            lcout => \b2v_inst200.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73351_5_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17128\,
            in1 => \N__25210\,
            in2 => \_gnd_net_\,
            in3 => \N__18802\,
            lcout => \b2v_inst200.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9551_7_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25211\,
            in1 => \N__17119\,
            in2 => \_gnd_net_\,
            in3 => \N__18778\,
            lcout => \b2v_inst200.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_14_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.count_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__20944\,
            sr => \N__20796\
        );

    \b2v_inst16.count_RNIJP141_14_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15412\,
            in1 => \N__20912\,
            in2 => \_gnd_net_\,
            in3 => \N__15405\,
            lcout => \b2v_inst16.countZ0Z_14\,
            ltout => \b2v_inst16.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_13_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__15633\,
            in1 => \N__15390\,
            in2 => \N__15364\,
            in3 => \N__15361\,
            lcout => \b2v_inst16.count_4_i_a3_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIHM041_13_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15592\,
            in1 => \N__20911\,
            in2 => \_gnd_net_\,
            in3 => \N__15600\,
            lcout => \b2v_inst16.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15618\,
            in1 => \N__16025\,
            in2 => \N__15637\,
            in3 => \N__15895\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIHAVJ1_4_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15607\,
            in2 => \N__15640\,
            in3 => \N__20910\,
            lcout => \b2v_inst16.countZ0Z_4\,
            ltout => \b2v_inst16.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_4_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__15619\,
            in1 => \N__16026\,
            in2 => \N__15610\,
            in3 => \N__15896\,
            lcout => \b2v_inst16.count_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__20944\,
            sr => \N__20796\
        );

    \b2v_inst16.count_13_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15601\,
            lcout => \b2v_inst16.count_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36602\,
            ce => \N__20944\,
            sr => \N__20796\
        );

    \b2v_inst16.count_RNI2J651_0_1_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15502\,
            in1 => \N__20882\,
            in2 => \_gnd_net_\,
            in3 => \N__15490\,
            lcout => \b2v_inst16.un4_count_1_axb_1\,
            ltout => \b2v_inst16.un4_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI_1_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__15712\,
            in1 => \_gnd_net_\,
            in2 => \N__15586\,
            in3 => \N__15982\,
            lcout => \b2v_inst16.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_1_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__15710\,
            in2 => \_gnd_net_\,
            in3 => \N__15583\,
            lcout => \b2v_inst16.count_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36597\,
            ce => \N__20914\,
            sr => \N__20789\
        );

    \b2v_inst16.count_RNIKN901_0_12_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15571\,
            in1 => \N__15553\,
            in2 => \N__15541\,
            in3 => \N__15520\,
            lcout => \b2v_inst16.count_4_i_a3_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI2J651_1_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20915\,
            in1 => \N__15501\,
            in2 => \_gnd_net_\,
            in3 => \N__15489\,
            lcout => OPEN,
            ltout => \b2v_inst16.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNI2J651_2_1_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__15477\,
            in1 => \_gnd_net_\,
            in2 => \N__15463\,
            in3 => \N__15460\,
            lcout => OPEN,
            ltout => \b2v_inst16.count_4_i_a3_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_RNIMAG52_12_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15751\,
            in1 => \N__15742\,
            in2 => \N__15736\,
            in3 => \N__15733\,
            lcout => \b2v_inst16.N_414\,
            ltout => \b2v_inst16.N_414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_0_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__15711\,
            in1 => \_gnd_net_\,
            in2 => \N__15679\,
            in3 => \N__15984\,
            lcout => \b2v_inst16.count_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36597\,
            ce => \N__20914\,
            sr => \N__20789\
        );

    \b2v_inst11.count_off_RNI5BGAF_1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__19318\,
            in1 => \N__15655\,
            in2 => \N__19485\,
            in3 => \N__15664\,
            lcout => \b2v_inst11.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4AGAF_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__17170\,
            in1 => \N__19431\,
            in2 => \N__15649\,
            in3 => \N__19317\,
            lcout => \b2v_inst11.count_offZ0Z_0\,
            ltout => \b2v_inst11.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_1_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15667\,
            in3 => \N__19145\,
            lcout => \b2v_inst11.count_off_RNIZ0Z_1\,
            ltout => \b2v_inst11.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_1_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15658\,
            in3 => \N__19323\,
            lcout => \b2v_inst11.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36592\,
            ce => \N__19484\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_0_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__19320\,
            in1 => \N__17171\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36592\,
            ce => \N__19484\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_10_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17241\,
            in2 => \_gnd_net_\,
            in3 => \N__19321\,
            lcout => \b2v_inst11.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36592\,
            ce => \N__19484\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIRKFDF_10_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__19319\,
            in1 => \N__15913\,
            in2 => \N__19486\,
            in3 => \N__17242\,
            lcout => \b2v_inst11.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_13_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17373\,
            in2 => \_gnd_net_\,
            in3 => \N__19322\,
            lcout => \b2v_inst11.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36592\,
            ce => \N__19484\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI3B692_0_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15773\,
            in2 => \_gnd_net_\,
            in3 => \N__15807\,
            lcout => \b2v_inst16.N_1440\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI3B692_0_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__21140\,
            in1 => \N__35904\,
            in2 => \N__15811\,
            in3 => \N__15817\,
            lcout => \b2v_inst16.curr_state_RNI3B692Z0Z_0\,
            ltout => \b2v_inst16.curr_state_RNI3B692Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_1_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__15809\,
            in1 => \N__21142\,
            in2 => \N__15901\,
            in3 => \N__15897\,
            lcout => \b2v_inst16.curr_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36589\,
            ce => \N__36369\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIERV34_0_0_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001011111"
        )
    port map (
            in0 => \N__21139\,
            in1 => \N__15894\,
            in2 => \N__15778\,
            in3 => \N__15810\,
            lcout => OPEN,
            ltout => \b2v_inst16.curr_state_7_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI7NCI4_1_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__35903\,
            in1 => \_gnd_net_\,
            in2 => \N__15829\,
            in3 => \N__15826\,
            lcout => \b2v_inst16.curr_stateZ0Z_1\,
            ltout => \b2v_inst16.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__21141\,
            in1 => \_gnd_net_\,
            in2 => \N__15820\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst16.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36589\,
            ce => \N__36369\,
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNIERV34_0_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__15808\,
            in1 => \N__15772\,
            in2 => \_gnd_net_\,
            in3 => \N__21138\,
            lcout => \b2v_inst16.N_268\,
            ltout => \b2v_inst16.N_268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_RNI68A74_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16060\,
            in3 => \N__35902\,
            lcout => \b2v_inst16.N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNILCR74_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__16113\,
            in1 => \N__17834\,
            in2 => \N__16141\,
            in3 => \N__16213\,
            lcout => \b2v_inst11.N_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__24397\,
            in1 => \N__24641\,
            in2 => \_gnd_net_\,
            in3 => \N__23381\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__21201\,
            in1 => \N__23704\,
            in2 => \N__15925\,
            in3 => \N__17746\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_329_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIF6NL_9_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__24393\,
            in1 => \N__24149\,
            in2 => \N__17752\,
            in3 => \N__23382\,
            lcout => \b2v_inst11.N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINPGR_2_1_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__24640\,
            in1 => \N__24396\,
            in2 => \N__24161\,
            in3 => \N__27142\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_RNINPGR_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI608H1_0_1_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100011111"
        )
    port map (
            in0 => \N__23705\,
            in1 => \N__26632\,
            in2 => \N__15922\,
            in3 => \N__23426\,
            lcout => \b2v_inst11.func_state_RNI608H1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__24150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24394\,
            lcout => b2v_inst11_dutycycle_1_0_iv_0_o3_out,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_0_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100111111"
        )
    port map (
            in0 => \N__24395\,
            in1 => \N__24151\,
            in2 => \N__23720\,
            in3 => \N__19849\,
            lcout => \b2v_inst11.g0_20_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16114\,
            in1 => \N__23887\,
            in2 => \N__18718\,
            in3 => \N__16189\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__23702\,
            in1 => \N__16084\,
            in2 => \N__16144\,
            in3 => \N__16134\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_func_state25_6_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_en_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__17575\,
            in1 => \N__16123\,
            in2 => \N__16117\,
            in3 => \N__27722\,
            lcout => \b2v_inst11.count_off_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIC9BO3_1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001100"
        )
    port map (
            in0 => \N__24469\,
            in1 => \N__24213\,
            in2 => \N__35938\,
            in3 => \N__16195\,
            lcout => \b2v_inst11.N_430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_0_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23701\,
            in2 => \_gnd_net_\,
            in3 => \N__19841\,
            lcout => \b2v_inst11.func_state_RNI_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_1_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__23703\,
            in1 => \_gnd_net_\,
            in2 => \N__27149\,
            in3 => \N__29398\,
            lcout => \N_236_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIEJ1N1_0_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__24639\,
            in1 => \N__18496\,
            in2 => \N__24519\,
            in3 => \N__19842\,
            lcout => \b2v_inst11.g1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23886\,
            in1 => \N__18717\,
            in2 => \N__27148\,
            in3 => \N__17745\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_331_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIH4KN3_0_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__24606\,
            in1 => \N__33781\,
            in2 => \N__16069\,
            in3 => \N__16162\,
            lcout => \b2v_inst11.count_clk_en_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_0_1_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26941\,
            in1 => \N__23696\,
            in2 => \N__23390\,
            in3 => \N__17741\,
            lcout => \b2v_inst11.N_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIMFI92_1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17798\,
            in1 => \N__22496\,
            in2 => \_gnd_net_\,
            in3 => \N__16187\,
            lcout => \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI5M9V2_9_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__23068\,
            in1 => \N__16204\,
            in2 => \N__27150\,
            in3 => \N__17799\,
            lcout => \b2v_inst11.func_state_1_ss0_i_0_o3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI8JP5_1_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24605\,
            in1 => \N__16188\,
            in2 => \N__17751\,
            in3 => \N__21672\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_9_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17740\,
            lcout => \b2v_inst11.count_off_RNIZ0Z_9\,
            ltout => \b2v_inst11.count_off_RNIZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_1_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__23695\,
            in1 => \_gnd_net_\,
            in2 => \N__16168\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.func_state_RNI_1Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNI_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_3_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000111"
        )
    port map (
            in0 => \N__19843\,
            in1 => \N__23697\,
            in2 => \N__16165\,
            in3 => \N__17797\,
            lcout => \b2v_inst11.un1_func_state25_4_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16878\,
            in1 => \N__16370\,
            in2 => \_gnd_net_\,
            in3 => \N__16334\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI2UQ9_1_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16150\,
            in2 => \N__16156\,
            in3 => \N__18048\,
            lcout => \b2v_inst11.count_clkZ0Z_1\,
            ltout => \b2v_inst11.count_clkZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_1_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__16879\,
            in1 => \_gnd_net_\,
            in2 => \N__16153\,
            in3 => \N__16336\,
            lcout => \b2v_inst11.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36583\,
            ce => \N__18118\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_0_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16880\,
            lcout => \b2v_inst11.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36583\,
            ce => \N__18118\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI1TQ9_0_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18050\,
            in1 => \N__16246\,
            in2 => \_gnd_net_\,
            in3 => \N__16228\,
            lcout => \b2v_inst11.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI9KMF_7_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16543\,
            in1 => \N__16240\,
            in2 => \_gnd_net_\,
            in3 => \N__18049\,
            lcout => \b2v_inst11.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_7_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16542\,
            lcout => \b2v_inst11.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36583\,
            ce => \N__18118\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICQPCF_6_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19072\,
            in1 => \N__19458\,
            in2 => \_gnd_net_\,
            in3 => \N__19567\,
            lcout => \b2v_inst11.un3_count_off_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__23878\,
            in1 => \N__24366\,
            in2 => \_gnd_net_\,
            in3 => \N__24132\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_168_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNICGI84_0_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__24500\,
            in1 => \N__35892\,
            in2 => \N__16234\,
            in3 => \N__16381\,
            lcout => \b2v_inst11.func_state_RNICGI84_0_0\,
            ltout => \b2v_inst11.func_state_RNICGI84_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_0_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16231\,
            in3 => \N__16337\,
            lcout => \b2v_inst11.count_clk_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_0_0_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__26942\,
            in1 => \N__23365\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.func_state_RNIVS8U1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI505F_14_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16926\,
            in2 => \N__18068\,
            in3 => \N__16393\,
            lcout => \b2v_inst11.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIN9J12_1_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__24211\,
            in1 => \N__23877\,
            in2 => \N__24515\,
            in3 => \N__35891\,
            lcout => \b2v_inst11.N_338\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI608H1_0_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__17750\,
            in1 => \N__23699\,
            in2 => \N__19840\,
            in3 => \N__16387\,
            lcout => \b2v_inst11.un1_count_clk_1_sqmuxa_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_0_1_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__23700\,
            in1 => \N__23366\,
            in2 => \N__29400\,
            in3 => \N__23472\,
            lcout => b2v_inst11_un1_dutycycle_172_m3_amcf1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16375\,
            in2 => \N__16342\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16877\,
            in1 => \N__18360\,
            in2 => \_gnd_net_\,
            in3 => \N__16297\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_1\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16872\,
            in1 => \N__17905\,
            in2 => \_gnd_net_\,
            in3 => \N__16294\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_2\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16291\,
            in2 => \_gnd_net_\,
            in3 => \N__16252\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_3\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16873\,
            in1 => \N__18321\,
            in2 => \_gnd_net_\,
            in3 => \N__16249\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_4\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16875\,
            in1 => \N__17874\,
            in2 => \_gnd_net_\,
            in3 => \N__16576\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_5\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16874\,
            in1 => \N__16573\,
            in2 => \_gnd_net_\,
            in3 => \N__16531\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_6\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16876\,
            in1 => \N__18428\,
            in2 => \_gnd_net_\,
            in3 => \N__16528\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_7_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16885\,
            in1 => \N__18256\,
            in2 => \_gnd_net_\,
            in3 => \N__16525\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5\,
            ltout => OPEN,
            carryin => \bfn_2_13_0_\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16522\,
            in2 => \_gnd_net_\,
            in3 => \N__16504\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_9_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16500\,
            in2 => \_gnd_net_\,
            in3 => \N__16477\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_10_cZ0\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16473\,
            in2 => \_gnd_net_\,
            in3 => \N__16453\,
            lcout => \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_11\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16884\,
            in1 => \N__16450\,
            in2 => \_gnd_net_\,
            in3 => \N__16414\,
            lcout => \b2v_inst11.count_clk_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_12\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__16887\,
            in1 => \N__16411\,
            in2 => \_gnd_net_\,
            in3 => \N__16906\,
            lcout => \b2v_inst11.count_clk_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_clk_2_cry_13\,
            carryout => \b2v_inst11.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__16903\,
            in1 => \_gnd_net_\,
            in2 => \N__16888\,
            in3 => \N__16798\,
            lcout => \b2v_inst11.count_clk_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_9_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36591\,
            ce => \N__18091\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_RNO_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16779\,
            in1 => \N__16767\,
            in2 => \N__16756\,
            in3 => \N__16740\,
            lcout => \b2v_inst20.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_RNO_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16728\,
            in1 => \N__16716\,
            in2 => \N__16705\,
            in3 => \N__16689\,
            lcout => \b2v_inst20.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_RNO_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16677\,
            in1 => \N__16665\,
            in2 => \N__16654\,
            in3 => \N__16638\,
            lcout => \b2v_inst20.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_RNO_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16626\,
            in1 => \N__16614\,
            in2 => \N__16603\,
            in3 => \N__16587\,
            lcout => \b2v_inst20.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_4_1_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19947\,
            in1 => \N__23879\,
            in2 => \_gnd_net_\,
            in3 => \N__29388\,
            lcout => \func_state_RNIVS8U1_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.un1_vddq_en_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__21199\,
            in1 => \N__16981\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \VDDQ_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18520\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_15_0_\,
            carryout => \b2v_inst20.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20302\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_0\,
            carryout => \b2v_inst20.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_2_c_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16957\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_1\,
            carryout => \b2v_inst20.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_3_c_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16948\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_2\,
            carryout => \b2v_inst20.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_4_c_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16939\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_3\,
            carryout => \b2v_inst20.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_5_c_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16933\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_4\,
            carryout => \b2v_inst20.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16999\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_5\,
            carryout => \b2v_inst20.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17056\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst20.un4_counter_6\,
            carryout => b2v_inst20_un4_counter_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17110\,
            lcout => \b2v_inst20_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_7_c_RNO_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17106\,
            in1 => \N__17094\,
            in2 => \N__17083\,
            in3 => \N__17067\,
            lcout => \b2v_inst20.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_6_c_RNO_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17049\,
            in1 => \N__17037\,
            in2 => \N__17026\,
            in3 => \N__17010\,
            lcout => \b2v_inst20.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_1_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18829\,
            in1 => \N__18853\,
            in2 => \N__18571\,
            in3 => \N__18544\,
            lcout => \b2v_inst200.un25_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIP16E1_1_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18555\,
            in1 => \N__16993\,
            in2 => \_gnd_net_\,
            in3 => \N__25206\,
            lcout => \b2v_inst200.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_1_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18556\,
            lcout => \b2v_inst200.count_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36627\,
            ce => \N__25154\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QV41_2_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__16987\,
            in1 => \N__18531\,
            in2 => \_gnd_net_\,
            in3 => \N__25207\,
            lcout => \b2v_inst200.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_2_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18532\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36627\,
            ce => \N__25154\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI3T051_3_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17149\,
            in1 => \N__25208\,
            in2 => \_gnd_net_\,
            in3 => \N__18840\,
            lcout => \b2v_inst200.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_3_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36627\,
            ce => \N__25154\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50251_4_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17134\,
            in1 => \N__25209\,
            in2 => \_gnd_net_\,
            in3 => \N__18816\,
            lcout => \b2v_inst200.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_12_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18903\,
            lcout => \b2v_inst200.count_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36623\,
            ce => \N__25153\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_13_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20644\,
            lcout => \b2v_inst200.count_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36623\,
            ce => \N__25153\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_4_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18817\,
            lcout => \b2v_inst200.count_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36623\,
            ce => \N__25153\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_5_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18798\,
            lcout => \b2v_inst200.count_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36623\,
            ce => \N__25153\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_7_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18774\,
            lcout => \b2v_inst200.count_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36623\,
            ce => \N__25153\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_17_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18865\,
            lcout => \b2v_inst200.count_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36623\,
            ce => \N__25153\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICFRGF_15_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19533\,
            in1 => \N__17221\,
            in2 => \N__19351\,
            in3 => \N__17328\,
            lcout => \b2v_inst11.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_15_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17332\,
            in3 => \N__19347\,
            lcout => \b2v_inst11.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36617\,
            ce => \N__19536\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI89PGF_13_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19531\,
            in1 => \N__17215\,
            in2 => \N__17377\,
            in3 => \N__19348\,
            lcout => \b2v_inst11.count_offZ0Z_13\,
            ltout => \b2v_inst11.count_offZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI_15_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18934\,
            in1 => \N__17191\,
            in2 => \N__17203\,
            in3 => \N__17346\,
            lcout => \b2v_inst11.un34_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_8_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17256\,
            in2 => \_gnd_net_\,
            in3 => \N__19350\,
            lcout => \b2v_inst11.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36617\,
            ce => \N__19536\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIG0SCF_8_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19349\,
            in1 => \N__17200\,
            in2 => \N__17260\,
            in3 => \N__19532\,
            lcout => \b2v_inst11.count_offZ0Z_8\,
            ltout => \b2v_inst11.count_offZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIETQCF_0_7_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__19549\,
            in1 => \N__19534\,
            in2 => \N__17194\,
            in3 => \N__19216\,
            lcout => \b2v_inst11.un34_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIETQCF_7_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19535\,
            in1 => \N__19548\,
            in2 => \_gnd_net_\,
            in3 => \N__19215\,
            lcout => \b2v_inst11.un3_count_off_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19149\,
            in2 => \N__17190\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_4_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18913\,
            in2 => \_gnd_net_\,
            in3 => \N__17155\,
            lcout => \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_1\,
            carryout => \b2v_inst11.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19012\,
            in2 => \_gnd_net_\,
            in3 => \N__17152\,
            lcout => \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_2\,
            carryout => \b2v_inst11.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19006\,
            in2 => \_gnd_net_\,
            in3 => \N__17302\,
            lcout => \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_3\,
            carryout => \b2v_inst11.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19164\,
            in2 => \_gnd_net_\,
            in3 => \N__17299\,
            lcout => \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_4\,
            carryout => \b2v_inst11.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17296\,
            in2 => \_gnd_net_\,
            in3 => \N__17281\,
            lcout => \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_5\,
            carryout => \b2v_inst11.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17278\,
            in3 => \N__17269\,
            lcout => \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_6\,
            carryout => \b2v_inst11.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17266\,
            in2 => \_gnd_net_\,
            in3 => \N__17248\,
            lcout => \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_7\,
            carryout => \b2v_inst11.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19021\,
            in2 => \_gnd_net_\,
            in3 => \N__17245\,
            lcout => \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \b2v_inst11.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17454\,
            in2 => \_gnd_net_\,
            in3 => \N__17227\,
            lcout => \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_9\,
            carryout => \b2v_inst11.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17317\,
            in2 => \_gnd_net_\,
            in3 => \N__17224\,
            lcout => \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_10\,
            carryout => \b2v_inst11.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17472\,
            in2 => \_gnd_net_\,
            in3 => \N__17389\,
            lcout => \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_11\,
            carryout => \b2v_inst11.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17386\,
            in2 => \_gnd_net_\,
            in3 => \N__17356\,
            lcout => \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_12\,
            carryout => \b2v_inst11.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18933\,
            in2 => \_gnd_net_\,
            in3 => \N__17353\,
            lcout => \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un3_count_off_1_cry_13\,
            carryout => \b2v_inst11.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17350\,
            in2 => \_gnd_net_\,
            in3 => \N__17335\,
            lcout => \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_1_c_RNIJE0A4_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19186\,
            in2 => \_gnd_net_\,
            in3 => \N__19343\,
            lcout => \b2v_inst11.count_off_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_12_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17493\,
            in2 => \_gnd_net_\,
            in3 => \N__19341\,
            lcout => \b2v_inst11.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36599\,
            ce => \N__19517\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI43NGF_11_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17311\,
            in1 => \N__17409\,
            in2 => \_gnd_net_\,
            in3 => \N__19516\,
            lcout => \b2v_inst11.un3_count_off_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_10_c_RNI3CGD4_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17419\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19342\,
            lcout => \b2v_inst11.count_off_1_11\,
            ltout => \b2v_inst11.count_off_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI43NGF_0_11_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__17473\,
            in1 => \N__17410\,
            in2 => \N__17305\,
            in3 => \N__19518\,
            lcout => \b2v_inst11.un34_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI66OGF_12_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__19515\,
            in1 => \N__17494\,
            in2 => \N__17482\,
            in3 => \N__19339\,
            lcout => \b2v_inst11.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNII3TCF_0_9_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__19036\,
            in1 => \N__19042\,
            in2 => \N__17461\,
            in3 => \N__19519\,
            lcout => OPEN,
            ltout => \b2v_inst11.un34_clk_100khz_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIQTKGS2_9_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17437\,
            in1 => \N__19099\,
            in2 => \N__17431\,
            in3 => \N__17428\,
            lcout => \b2v_inst11.count_off_RNIQTKGS2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_11_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19340\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17418\,
            lcout => \b2v_inst11.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36599\,
            ce => \N__19517\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_7_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001100110011"
        )
    port map (
            in0 => \N__17554\,
            in1 => \N__17395\,
            in2 => \N__23043\,
            in3 => \N__17539\,
            lcout => \b2v_inst11.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36594\,
            ce => 'H',
            sr => \N__25981\
        );

    \b2v_inst11.dutycycle_RNI863D_2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101011111"
        )
    port map (
            in0 => \N__24103\,
            in1 => \N__23694\,
            in2 => \N__27151\,
            in3 => \N__30298\,
            lcout => OPEN,
            ltout => \b2v_inst11.g4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIGT0G4_2_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__22991\,
            in1 => \N__24622\,
            in2 => \N__17401\,
            in3 => \N__33784\,
            lcout => \b2v_inst11.g1_0_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIVTQU_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__24392\,
            in1 => \N__21481\,
            in2 => \N__24128\,
            in3 => \N__23693\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_17_N_3L3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIVGS13_7_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110111011"
        )
    port map (
            in0 => \N__27724\,
            in1 => \N__17553\,
            in2 => \N__17398\,
            in3 => \N__23894\,
            lcout => \b2v_inst11.dutycycle_RNIVGS13Z0Z_7\,
            ltout => \b2v_inst11.dutycycle_RNIVGS13Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIJI0UD_7_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101100001111"
        )
    port map (
            in0 => \N__17552\,
            in1 => \N__17538\,
            in2 => \N__17524\,
            in3 => \N__22987\,
            lcout => \b2v_inst11.dutycycleZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_ss0_i_0_x2_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24391\,
            in2 => \_gnd_net_\,
            in3 => \N__24104\,
            lcout => \b2v_inst11.N_160_i\,
            ltout => \b2v_inst11.N_160_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_5_1_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23895\,
            in1 => \N__23376\,
            in2 => \N__17521\,
            in3 => \N__17842\,
            lcout => \b2v_inst11.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_1_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__23714\,
            in1 => \N__23482\,
            in2 => \N__23907\,
            in3 => \N__21419\,
            lcout => \b2v_inst11.N_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_3_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__28756\,
            in1 => \N__21602\,
            in2 => \N__29539\,
            in3 => \N__26977\,
            lcout => g0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIUPHS3_6_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111100"
        )
    port map (
            in0 => \N__17560\,
            in1 => \N__25840\,
            in2 => \N__19195\,
            in3 => \N__19639\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIERM9C_2_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__22986\,
            in1 => \N__17518\,
            in2 => \N__17509\,
            in3 => \N__33783\,
            lcout => \b2v_inst11.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_8_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__26188\,
            in1 => \N__26329\,
            in2 => \_gnd_net_\,
            in3 => \N__29526\,
            lcout => \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNISM1B4_6_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011110000"
        )
    port map (
            in0 => \N__18508\,
            in1 => \N__17506\,
            in2 => \N__26197\,
            in3 => \N__23899\,
            lcout => \b2v_inst11.N_231_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_3_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28758\,
            in3 => \N__29525\,
            lcout => \b2v_inst11.N_354\,
            ltout => \b2v_inst11.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29399\,
            in1 => \N__21603\,
            in2 => \N__17593\,
            in3 => \N__26976\,
            lcout => b2v_inst11_g0_i_m2_i_a6_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__23356\,
            in1 => \N__19728\,
            in2 => \N__19847\,
            in3 => \N__20038\,
            lcout => \b2v_inst11.N_159\,
            ltout => \b2v_inst11.N_159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_6_0_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__20695\,
            in1 => \_gnd_net_\,
            in2 => \N__17581\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_425\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI7J1P_0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__24361\,
            in1 => \N__24052\,
            in2 => \N__19848\,
            in3 => \N__35897\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m0_0_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIT2K23_1_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__17727\,
            in1 => \N__22498\,
            in2 => \N__17578\,
            in3 => \N__23716\,
            lcout => \b2v_inst11.func_state_1_m0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27064\,
            in1 => \N__20697\,
            in2 => \N__26947\,
            in3 => \N__20040\,
            lcout => \b2v_inst11.un1_func_state25_6_0_o_N_313_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI_0_6_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27063\,
            in2 => \_gnd_net_\,
            in3 => \N__26587\,
            lcout => \b2v_inst11.N_19_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIF6NL_6_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101111"
        )
    port map (
            in0 => \N__23499\,
            in1 => \N__20696\,
            in2 => \N__26633\,
            in3 => \N__20039\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIVS8U1_6_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__22036\,
            in1 => \N__20293\,
            in2 => \N__17563\,
            in3 => \N__22120\,
            lcout => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_5_1_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24190\,
            in2 => \_gnd_net_\,
            in3 => \N__23322\,
            lcout => \b2v_inst11.func_state_RNI_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_2_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23638\,
            lcout => \b2v_inst11.func_state_RNI_2Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_6_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__27102\,
            in1 => \N__20694\,
            in2 => \N__17638\,
            in3 => \N__19726\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m2s2_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICME96_6_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__23060\,
            in1 => \N__17635\,
            in2 => \N__17623\,
            in3 => \N__17620\,
            lcout => \b2v_inst11.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_6_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19727\,
            in2 => \_gnd_net_\,
            in3 => \N__20693\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_5Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIOSKL1_6_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21665\,
            in1 => \N__24102\,
            in2 => \N__17608\,
            in3 => \N__23852\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIH3TI8_6_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111111"
        )
    port map (
            in0 => \N__19738\,
            in1 => \N__17605\,
            in2 => \N__17596\,
            in3 => \N__23059\,
            lcout => \b2v_inst11.dutycycle_e_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_1_1_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23125\,
            in1 => \N__23639\,
            in2 => \N__23519\,
            in3 => \N__26568\,
            lcout => \b2v_inst11.un1_clk_100khz_43_and_i_0_ccf1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI5M9V2_0_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__17763\,
            in1 => \N__22483\,
            in2 => \N__23375\,
            in3 => \N__19760\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m2_am_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIR5S85_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__17841\,
            in1 => \N__23061\,
            in2 => \N__17809\,
            in3 => \N__17806\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_RNIR5S85Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIMLUM9_0_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17661\,
            in1 => \_gnd_net_\,
            in2 => \N__17782\,
            in3 => \N__19879\,
            lcout => \b2v_inst11.func_state_1_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI7762C_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__17948\,
            in1 => \N__21164\,
            in2 => \N__17776\,
            in3 => \N__17646\,
            lcout => \b2v_inst11.func_state\,
            ltout => \b2v_inst11.func_state_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_2_0_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17779\,
            in3 => \_gnd_net_\,
            lcout => \func_state_RNI_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__17775\,
            in1 => \N__21165\,
            in2 => \N__17955\,
            in3 => \N__17647\,
            lcout => \b2v_inst11.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36593\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_0_0_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__17764\,
            in1 => \N__17736\,
            in2 => \N__17662\,
            in3 => \N__19761\,
            lcout => OPEN,
            ltout => \b2v_inst11.func_state_1_m2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIOIMG7_1_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__19896\,
            in1 => \N__17674\,
            in2 => \N__17665\,
            in3 => \N__17657\,
            lcout => \b2v_inst11.func_state_1_m2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_1_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__21177\,
            in1 => \N__17947\,
            in2 => \N__17971\,
            in3 => \N__17923\,
            lcout => \b2v_inst11.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__22035\,
            in1 => \N__20289\,
            in2 => \N__23532\,
            in3 => \N__22114\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_fast_RNITMQQ5_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111100"
        )
    port map (
            in0 => \N__27163\,
            in1 => \N__19988\,
            in2 => \N__17986\,
            in3 => \N__19964\,
            lcout => \N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_1_1_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__26634\,
            in1 => \N__23857\,
            in2 => \N__23533\,
            in3 => \N__23632\,
            lcout => \b2v_inst11.N_326_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_en_0_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__24920\,
            in1 => \N__24845\,
            in2 => \N__24101\,
            in3 => \N__33725\,
            lcout => \b2v_inst11.count_clk_enZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.VCCST_EN_i_0_o3_0_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111111011111"
        )
    port map (
            in0 => \N__21987\,
            in1 => \N__35820\,
            in2 => \N__24100\,
            in3 => \N__22113\,
            lcout => \VCCST_EN_i_0_o3_0\,
            ltout => \VCCST_EN_i_0_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI6BE8E_1_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__17967\,
            in1 => \N__17946\,
            in2 => \N__17926\,
            in3 => \N__17922\,
            lcout => \func_state_RNI6BE8E_0_1\,
            ltout => \func_state_RNI6BE8E_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_1_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17914\,
            in3 => \N__23349\,
            lcout => \b2v_inst11.N_172\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIU6GN_7_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__24691\,
            in1 => \N__35827\,
            in2 => \_gnd_net_\,
            in3 => \N__17911\,
            lcout => \b2v_inst11.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_7_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24690\,
            lcout => \b2v_inst11.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36603\,
            ce => \N__36363\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI18IF_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18232\,
            in2 => \N__18114\,
            in3 => \N__18214\,
            lcout => \b2v_inst11.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI7HLF_6_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18178\,
            in1 => \N__18154\,
            in2 => \_gnd_net_\,
            in3 => \N__18106\,
            lcout => \b2v_inst11.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIBNNF_8_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18148\,
            in2 => \N__18112\,
            in3 => \N__18124\,
            lcout => \b2v_inst11.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIV4HF_2_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18391\,
            in1 => \N__18373\,
            in2 => \_gnd_net_\,
            in3 => \N__18102\,
            lcout => \b2v_inst11.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI5EKF_5_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18184\,
            in2 => \N__18113\,
            in3 => \N__18208\,
            lcout => \b2v_inst11.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIDQOF_9_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18283\,
            in1 => \N__18268\,
            in2 => \_gnd_net_\,
            in3 => \N__18095\,
            lcout => \b2v_inst11.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_3_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18231\,
            lcout => \b2v_inst11.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36611\,
            ce => \N__18111\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_5_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18207\,
            lcout => \b2v_inst11.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36611\,
            ce => \N__18111\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_6_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18177\,
            lcout => \b2v_inst11.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36611\,
            ce => \N__18111\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_8_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18147\,
            lcout => \b2v_inst11.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36611\,
            ce => \N__18111\,
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_0_c_RNO_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18736\,
            in1 => \N__18587\,
            in2 => \N__18450\,
            in3 => \N__18668\,
            lcout => \b2v_inst20.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__24581\,
            in1 => \N__24924\,
            in2 => \N__24520\,
            in3 => \N__23757\,
            lcout => \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINPGR_0_1_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011000100"
        )
    port map (
            in0 => \N__24318\,
            in1 => \N__23655\,
            in2 => \N__24056\,
            in3 => \N__24582\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI608H1_1_1_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110011"
        )
    port map (
            in0 => \N__24021\,
            in1 => \N__24317\,
            in2 => \N__18511\,
            in3 => \N__26642\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1\,
            ltout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNITPOC2_0_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__18699\,
            in1 => \_gnd_net_\,
            in2 => \N__18499\,
            in3 => \N__19839\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNINPGR_1_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000100010"
        )
    port map (
            in0 => \N__23656\,
            in1 => \N__24319\,
            in2 => \N__24604\,
            in3 => \N__24025\,
            lcout => \b2v_inst11.N_381_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_RNIQDE62_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__18484\,
            in1 => \N__21991\,
            in2 => \N__20287\,
            in3 => \N__22119\,
            lcout => \N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_3_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18466\,
            in1 => \N__18446\,
            in2 => \_gnd_net_\,
            in3 => \N__24849\,
            lcout => \b2v_inst20.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36616\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_0_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__24838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18741\,
            lcout => \b2v_inst20.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_1_LC_4_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18740\,
            in1 => \N__20322\,
            in2 => \_gnd_net_\,
            in3 => \N__24841\,
            lcout => \b2v_inst20.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_4_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__24562\,
            in1 => \N__23991\,
            in2 => \_gnd_net_\,
            in3 => \N__24308\,
            lcout => \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_4_LC_4_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__24837\,
            in1 => \N__18688\,
            in2 => \_gnd_net_\,
            in3 => \N__18672\,
            lcout => \b2v_inst20.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_5_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18652\,
            in1 => \N__20370\,
            in2 => \_gnd_net_\,
            in3 => \N__24840\,
            lcout => \b2v_inst20.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_0_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33688\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delayed_vccin_vccinaux_ok_RNI8L1J7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_2_LC_4_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18607\,
            in1 => \N__18591\,
            in2 => \_gnd_net_\,
            in3 => \N__24839\,
            lcout => \b2v_inst20.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36622\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_0_0_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__22317\,
            in1 => \N__20622\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_1_0\,
            ltout => OPEN,
            carryin => \bfn_5_1_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_1_cy\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_5_0_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18567\,
            in2 => \_gnd_net_\,
            in3 => \N__18547\,
            lcout => \b2v_inst200.count_RNIC03N_5Z0Z_0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_1_cy\,
            carryout => \b2v_inst200.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18543\,
            in2 => \_gnd_net_\,
            in3 => \N__18523\,
            lcout => \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_1\,
            carryout => \b2v_inst200.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18852\,
            in2 => \_gnd_net_\,
            in3 => \N__18832\,
            lcout => \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_2\,
            carryout => \b2v_inst200.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18828\,
            in2 => \_gnd_net_\,
            in3 => \N__18805\,
            lcout => \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_3\,
            carryout => \b2v_inst200.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20589\,
            in2 => \_gnd_net_\,
            in3 => \N__18784\,
            lcout => \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_4\,
            carryout => \b2v_inst200.un2_count_1_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20479\,
            in2 => \_gnd_net_\,
            in3 => \N__18781\,
            lcout => \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_5_cZ0\,
            carryout => \b2v_inst200.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20610\,
            in2 => \_gnd_net_\,
            in3 => \N__18760\,
            lcout => \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_6\,
            carryout => \b2v_inst200.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20469\,
            in2 => \_gnd_net_\,
            in3 => \N__18757\,
            lcout => \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0\,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25258\,
            in2 => \_gnd_net_\,
            in3 => \N__18754\,
            lcout => \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_8\,
            carryout => \b2v_inst200.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20995\,
            in3 => \N__18751\,
            lcout => \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_9\,
            carryout => \b2v_inst200.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21079\,
            in2 => \_gnd_net_\,
            in3 => \N__18907\,
            lcout => \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_10\,
            carryout => \b2v_inst200.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20409\,
            in2 => \_gnd_net_\,
            in3 => \N__18889\,
            lcout => \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_11\,
            carryout => \b2v_inst200.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20632\,
            in2 => \_gnd_net_\,
            in3 => \N__18886\,
            lcout => \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_12\,
            carryout => \b2v_inst200.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20520\,
            in2 => \_gnd_net_\,
            in3 => \N__18883\,
            lcout => \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_13\,
            carryout => \b2v_inst200.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20562\,
            in2 => \_gnd_net_\,
            in3 => \N__18880\,
            lcout => \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69\,
            ltout => OPEN,
            carryin => \b2v_inst200.un2_count_1_cry_14\,
            carryout => \b2v_inst200.un2_count_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21057\,
            in2 => \_gnd_net_\,
            in3 => \N__18877\,
            lcout => \b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \b2v_inst200.un2_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__21073\,
            in1 => \N__22313\,
            in2 => \_gnd_net_\,
            in3 => \N__18874\,
            lcout => \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDCT71_17_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18871\,
            in1 => \N__18864\,
            in2 => \_gnd_net_\,
            in3 => \N__25219\,
            lcout => \b2v_inst200.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_2_c_RNIKG1A4_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18990\,
            in2 => \_gnd_net_\,
            in3 => \N__19330\,
            lcout => \b2v_inst11.count_off_1_3\,
            ltout => \b2v_inst11.count_off_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI6HMCF_3_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18981\,
            in2 => \N__19015\,
            in3 => \N__19487\,
            lcout => \b2v_inst11.un3_count_off_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI8KNCF_4_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__19488\,
            in1 => \N__18969\,
            in2 => \N__18961\,
            in3 => \N__19331\,
            lcout => \b2v_inst11.count_offZ0Z_4\,
            ltout => \b2v_inst11.count_offZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI6HMCF_0_3_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__19000\,
            in1 => \N__18982\,
            in2 => \N__18994\,
            in3 => \N__19490\,
            lcout => \b2v_inst11.un34_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_3_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18991\,
            in2 => \_gnd_net_\,
            in3 => \N__19335\,
            lcout => \b2v_inst11.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36619\,
            ce => \N__19525\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_4_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19333\,
            in1 => \_gnd_net_\,
            in2 => \N__18973\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36619\,
            ce => \N__19525\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_14_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18942\,
            in2 => \_gnd_net_\,
            in3 => \N__19334\,
            lcout => \b2v_inst11.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36619\,
            ce => \N__19525\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIACQGF_14_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19332\,
            in1 => \N__18952\,
            in2 => \N__18946\,
            in3 => \N__19489\,
            lcout => \b2v_inst11.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4ELCF_0_2_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__19174\,
            in1 => \N__18921\,
            in2 => \N__19537\,
            in3 => \N__19165\,
            lcout => \b2v_inst11.un34_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4ELCF_2_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__18922\,
            in1 => \N__19173\,
            in2 => \_gnd_net_\,
            in3 => \N__19494\,
            lcout => \b2v_inst11.un3_count_off_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19185\,
            in2 => \_gnd_net_\,
            in3 => \N__19338\,
            lcout => \b2v_inst11.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36612\,
            ce => \N__19526\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNIANOCF_5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__19495\,
            in1 => \N__19092\,
            in2 => \N__19081\,
            in3 => \N__19336\,
            lcout => \b2v_inst11.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNICQPCF_0_6_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__19065\,
            in1 => \N__19563\,
            in2 => \N__19153\,
            in3 => \N__19530\,
            lcout => OPEN,
            ltout => \b2v_inst11.un34_clk_100khz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNI4N0JT1_2_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19123\,
            in1 => \N__19117\,
            in2 => \N__19111\,
            in3 => \N__19108\,
            lcout => \b2v_inst11.un34_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19337\,
            in1 => \_gnd_net_\,
            in2 => \N__19093\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36612\,
            ce => \N__19526\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_6_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19579\,
            in2 => \_gnd_net_\,
            in3 => \N__19328\,
            lcout => \b2v_inst11.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36605\,
            ce => \N__19521\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_9_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19327\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19050\,
            lcout => \b2v_inst11.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36605\,
            ce => \N__19521\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_8_c_RNIQS7A4_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19329\,
            lcout => \b2v_inst11.count_off_1_9\,
            ltout => \b2v_inst11.count_off_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_RNII3TCF_9_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19035\,
            in2 => \N__19024\,
            in3 => \N__19520\,
            lcout => \b2v_inst11.un3_count_off_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_5_c_RNINM4A4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19578\,
            in2 => \_gnd_net_\,
            in3 => \N__19325\,
            lcout => \b2v_inst11.count_off_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_off_7_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19362\,
            lcout => \b2v_inst11.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36605\,
            ce => \N__19521\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un3_count_off_1_cry_6_c_RNIOO5A4_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19324\,
            lcout => \b2v_inst11.count_off_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_15_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__29614\,
            in1 => \N__29731\,
            in2 => \_gnd_net_\,
            in3 => \N__22687\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIDGA72_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__23452\,
            in1 => \N__21508\,
            in2 => \N__23906\,
            in3 => \N__23721\,
            lcout => \b2v_inst11.N_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_12_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__29047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21402\,
            lcout => \b2v_inst11.N_360\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101010"
        )
    port map (
            in0 => \N__26328\,
            in1 => \N__29533\,
            in2 => \N__26196\,
            in3 => \N__26712\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_14_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__29730\,
            in1 => \N__26452\,
            in2 => \N__26750\,
            in3 => \N__21108\,
            lcout => \b2v_inst11.un2_count_clk_17_0_a2_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_6_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101011111"
        )
    port map (
            in0 => \N__23380\,
            in1 => \N__19732\,
            in2 => \N__21869\,
            in3 => \N__20698\,
            lcout => \b2v_inst11.g0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_1_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__21857\,
            in1 => \N__21271\,
            in2 => \N__21823\,
            in3 => \N__26650\,
            lcout => \b2v_inst11.dutycycle_RNI_9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_4_1_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21819\,
            in2 => \_gnd_net_\,
            in3 => \N__21853\,
            lcout => \b2v_inst11.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI2T5T7_3_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__23044\,
            in1 => \N__23229\,
            in2 => \N__19588\,
            in3 => \N__19603\,
            lcout => \b2v_inst11.dutycycle_eena_8\,
            ltout => \b2v_inst11.dutycycle_eena_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_3_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__19624\,
            in1 => \N__19630\,
            in2 => \N__19633\,
            in3 => \N__27721\,
            lcout => \b2v_inst11.dutycycle_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36595\,
            ce => 'H',
            sr => \N__25976\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_c_RNIBC872_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__23835\,
            in1 => \N__23709\,
            in2 => \N__23521\,
            in3 => \N__21343\,
            lcout => \b2v_inst11.dutycycle_rst_7\,
            ltout => \b2v_inst11.dutycycle_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIP1UUA_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__19623\,
            in1 => \N__27720\,
            in2 => \N__19615\,
            in3 => \N__19612\,
            lcout => \b2v_inst11.dutycycleZ0Z_3\,
            ltout => \b2v_inst11.dutycycleZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_3_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19606\,
            in3 => \N__23157\,
            lcout => \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_2_1_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23836\,
            in2 => \_gnd_net_\,
            in3 => \N__19597\,
            lcout => \b2v_inst11.un1_clk_100khz_43_and_i_0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIVS8U1_12_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001101"
        )
    port map (
            in0 => \N__23837\,
            in1 => \N__23483\,
            in2 => \N__29048\,
            in3 => \N__23710\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_307_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI9R6T4_12_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010101010"
        )
    port map (
            in0 => \N__27723\,
            in1 => \N__19699\,
            in2 => \N__19702\,
            in3 => \N__23045\,
            lcout => \b2v_inst11.dutycycle_RNI9R6T4Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_2_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__23231\,
            in1 => \N__25816\,
            in2 => \N__21301\,
            in3 => \N__19651\,
            lcout => \b2v_inst11.N_234_N\,
            ltout => \b2v_inst11.N_234_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI9R6T4_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__23047\,
            in1 => \N__19693\,
            in2 => \N__19684\,
            in3 => \N__27719\,
            lcout => \b2v_inst11.func_state_RNI9R6T4Z0Z_1\,
            ltout => \b2v_inst11.func_state_RNI9R6T4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIA3KA7_11_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__21457\,
            in1 => \N__19668\,
            in2 => \N__19681\,
            in3 => \N__25817\,
            lcout => \b2v_inst11.dutycycleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_11_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__25818\,
            in1 => \N__21456\,
            in2 => \N__19672\,
            in3 => \N__19678\,
            lcout => \b2v_inst11.dutycycleZ1Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36586\,
            ce => 'H',
            sr => \N__25948\
        );

    \b2v_inst11.dutycycle_RNI_2_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__26637\,
            in1 => \N__19660\,
            in2 => \N__21323\,
            in3 => \N__30279\,
            lcout => \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_14_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010101"
        )
    port map (
            in0 => \N__25815\,
            in1 => \N__23230\,
            in2 => \N__29737\,
            in3 => \N__26636\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_155_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIMBHI8_14_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__27718\,
            in1 => \N__23132\,
            in2 => \N__19645\,
            in3 => \N__23046\,
            lcout => \b2v_inst11.dutycycle_en_11\,
            ltout => \b2v_inst11.dutycycle_en_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_14_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__25819\,
            in1 => \N__22710\,
            in2 => \N__19642\,
            in3 => \N__22741\,
            lcout => \b2v_inst11.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36586\,
            ce => 'H',
            sr => \N__25948\
        );

    \b2v_inst11.func_state_RNIVS8U1_3_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111101"
        )
    port map (
            in0 => \N__22031\,
            in1 => \N__20288\,
            in2 => \N__19858\,
            in3 => \N__22115\,
            lcout => \func_state_RNIVS8U1_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI70K8_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24331\,
            in2 => \_gnd_net_\,
            in3 => \N__19762\,
            lcout => \b2v_inst11.N_305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIEIB72_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__23715\,
            in1 => \N__21496\,
            in2 => \N__23520\,
            in3 => \N__23874\,
            lcout => \b2v_inst11.N_301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_3_1_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21813\,
            lcout => \b2v_inst11.N_3060_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21379\,
            in1 => \N__29344\,
            in2 => \_gnd_net_\,
            in3 => \N__26102\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_6\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_6_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19708\,
            in3 => \N__20699\,
            lcout => \b2v_inst11.N_426_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_3_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111001110000"
        )
    port map (
            in0 => \N__28772\,
            in1 => \N__26337\,
            in2 => \N__26844\,
            in3 => \N__29482\,
            lcout => OPEN,
            ltout => \b2v_inst11.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_9_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101101000010"
        )
    port map (
            in0 => \N__26103\,
            in1 => \N__26448\,
            in2 => \N__19705\,
            in3 => \N__26830\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111011111"
        )
    port map (
            in0 => \N__24328\,
            in1 => \N__20277\,
            in2 => \N__21986\,
            in3 => \N__22093\,
            lcout => \N_15_i_0_a4_1_N_3L3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__24587\,
            in1 => \N__24934\,
            in2 => \N__24513\,
            in3 => \N__23853\,
            lcout => \b2v_inst11.N_382\,
            ltout => \b2v_inst11.N_382_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQ6_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__23057\,
            in1 => \N__19912\,
            in2 => \N__19906\,
            in3 => \N__27078\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNIF6NL_0_6_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__23509\,
            in1 => \N__26649\,
            in2 => \N__20041\,
            in3 => \N__20706\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_clk_RNI5FOR1_6_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__21978\,
            in1 => \N__35896\,
            in2 => \N__19903\,
            in3 => \N__22095\,
            lcout => \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIRF2E4_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111100001111"
        )
    port map (
            in0 => \N__24113\,
            in1 => \N__24330\,
            in2 => \N__19900\,
            in3 => \N__19756\,
            lcout => \b2v_inst11.func_state_RNIRF2E4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__21977\,
            in1 => \N__24111\,
            in2 => \N__35929\,
            in3 => \N__22094\,
            lcout => \VCCST_EN_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIF6NL_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__24112\,
            in1 => \N__24329\,
            in2 => \_gnd_net_\,
            in3 => \N__23587\,
            lcout => \b2v_inst11.un1_clk_100khz_2_i_o3_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIVS8U1_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__19813\,
            in1 => \N__26915\,
            in2 => \N__33617\,
            in3 => \N__23617\,
            lcout => \b2v_inst11.dutycycle_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI98672_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110001"
        )
    port map (
            in0 => \N__23618\,
            in1 => \N__21361\,
            in2 => \N__26931\,
            in3 => \N__19814\,
            lcout => \b2v_inst11.dutycycle_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI_0_0_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19815\,
            in1 => \N__20707\,
            in2 => \_gnd_net_\,
            in3 => \N__20021\,
            lcout => \b2v_inst11.func_state_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__21944\,
            in1 => \N__25548\,
            in2 => \_gnd_net_\,
            in3 => \N__22096\,
            lcout => \b2v_inst5.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36604\,
            ce => \N__36364\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21924\,
            lcout => \b2v_inst5.N_2897_i\,
            ltout => \b2v_inst5.N_2897_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22098\,
            in2 => \N__19930\,
            in3 => \N__25547\,
            lcout => OPEN,
            ltout => \b2v_inst5.m4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI1CVE1_0_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19927\,
            in2 => \N__19921\,
            in3 => \N__35819\,
            lcout => \b2v_inst5.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.g0_8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111111011"
        )
    port map (
            in0 => \N__23510\,
            in1 => \N__21979\,
            in2 => \N__24932\,
            in3 => \N__22097\,
            lcout => \b2v_inst11.N_165_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_1_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__21420\,
            in1 => \N__21324\,
            in2 => \_gnd_net_\,
            in3 => \N__33321\,
            lcout => OPEN,
            ltout => \b2v_inst11.g2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_12_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__29049\,
            in1 => \N__33595\,
            in2 => \N__19918\,
            in3 => \N__26190\,
            lcout => \b2v_inst11.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNISSAOS1_5_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__20146\,
            in1 => \N__20158\,
            in2 => \N__20167\,
            in3 => \N__27534\,
            lcout => \dutycycle_RNISSAOS1_0_5\,
            ltout => \dutycycle_RNISSAOS1_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19915\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_5\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_1_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26192\,
            in1 => \N__33597\,
            in2 => \N__20044\,
            in3 => \N__33322\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.N_224_i_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__24484\,
            in1 => \N__35826\,
            in2 => \N__23905\,
            in3 => \N__24586\,
            lcout => \b2v_inst11.N_224_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__29050\,
            in2 => \N__33353\,
            in3 => \N__21325\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_73_mux_i_i_o7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__33596\,
            in1 => \N__26635\,
            in2 => \N__20008\,
            in3 => \N__26191\,
            lcout => \N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI52GVC_5_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__20124\,
            in1 => \N__27688\,
            in2 => \N__27285\,
            in3 => \N__20005\,
            lcout => \b2v_inst11.N_73_mux_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIUNGA5_5_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100011011"
        )
    port map (
            in0 => \N__27687\,
            in1 => \N__20123\,
            in2 => \N__23058\,
            in3 => \N__20083\,
            lcout => \b2v_inst11.dutycycle_RNIUNGA5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI4NJR6_5_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__20125\,
            in1 => \N__19990\,
            in2 => \N__20101\,
            in3 => \N__19965\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_73_mux_i_i_a7_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI7JLNN_5_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19999\,
            in2 => \N__19993\,
            in3 => \N__26053\,
            lcout => \b2v_inst11.N_73_mux_i_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_0_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19989\,
            in2 => \_gnd_net_\,
            in3 => \N__19966\,
            lcout => OPEN,
            ltout => \N_73_mux_i_i_a7_4_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_fast_RNIVS8U1_0_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__19951\,
            in1 => \N__23792\,
            in2 => \N__19933\,
            in3 => \N__29329\,
            lcout => OPEN,
            ltout => \N_73_mux_i_i_a7_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI74U7G_5_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__20122\,
            in1 => \N__27552\,
            in2 => \N__20170\,
            in3 => \N__20094\,
            lcout => \b2v_inst11.N_73_mux_i_i_1\,
            ltout => \b2v_inst11.N_73_mux_i_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_5_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__20157\,
            in1 => \N__20145\,
            in2 => \N__20128\,
            in3 => \N__27535\,
            lcout => \b2v_inst11.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36618\,
            ce => 'H',
            sr => \N__25937\
        );

    \b2v_inst11.func_state_RNIDGAL3_0_0_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000111"
        )
    port map (
            in0 => \N__22066\,
            in1 => \N__20259\,
            in2 => \N__22021\,
            in3 => \N__20110\,
            lcout => \b2v_inst11.N_140_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_fast_RNIGMH81_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22009\,
            in2 => \N__20276\,
            in3 => \N__22065\,
            lcout => \RSMRSTn_fast_RNIGMH81\,
            ltout => \RSMRSTn_fast_RNIGMH81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_rep1_RNIABFM6_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__20065\,
            in1 => \_gnd_net_\,
            in2 => \N__20104\,
            in3 => \N__20082\,
            lcout => \N_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35887\,
            lcout => \SYNTHESIZED_WIRE_1keep_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_rep1_RNI07F73_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__24510\,
            in1 => \N__24580\,
            in2 => \N__24933\,
            in3 => \N__20081\,
            lcout => \b2v_inst20.tmp_1_rep1_RNI07FZ0Z73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.counter_6_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000110"
        )
    port map (
            in0 => \N__20059\,
            in1 => \N__20342\,
            in2 => \N__24864\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst20.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.un4_counter_1_c_RNO_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20392\,
            in1 => \N__20366\,
            in2 => \N__20346\,
            in3 => \N__20318\,
            lcout => \b2v_inst20.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_fast_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__20260\,
            in1 => \_gnd_net_\,
            in2 => \N__24865\,
            in3 => \_gnd_net_\,
            lcout => \SYNTHESIZED_WIRE_1keep_3_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36624\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_ATP_RNIQFGQ_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__35815\,
            in1 => \N__20215\,
            in2 => \N__20191\,
            in3 => \N__20203\,
            lcout => \HDA_SDO_ATP_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI_0_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__22186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22229\,
            lcout => \b2v_inst200.N_205\,
            ltout => \b2v_inst200.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010111011"
        )
    port map (
            in0 => \N__22595\,
            in1 => \N__20202\,
            in2 => \N__20209\,
            in3 => \N__33686\,
            lcout => \G_2734\,
            ltout => \G_2734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNI52VB_2_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20176\,
            in2 => \N__20206\,
            in3 => \N__35814\,
            lcout => \b2v_inst200.curr_stateZ0Z_2\,
            ltout => \b2v_inst200.curr_stateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.HDA_SDO_ATP_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__22230\,
            in1 => \_gnd_net_\,
            in2 => \N__20194\,
            in3 => \N__22190\,
            lcout => \b2v_inst200.HDA_SDO_ATP_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36628\,
            ce => \N__36357\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_2_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20182\,
            lcout => \b2v_inst200.curr_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36628\,
            ce => \N__36357\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_0_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011001101"
        )
    port map (
            in0 => \N__33687\,
            in1 => \N__22249\,
            in2 => \N__22195\,
            in3 => \N__22231\,
            lcout => \b2v_inst200.curr_state_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36628\,
            ce => \N__36357\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIDC651_8_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__25205\,
            in1 => \N__20431\,
            in2 => \N__22329\,
            in3 => \N__20439\,
            lcout => \b2v_inst200.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI96451_6_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20457\,
            in1 => \N__22318\,
            in2 => \N__20449\,
            in3 => \N__25204\,
            lcout => \b2v_inst200.countZ0Z_6\,
            ltout => \b2v_inst200.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_6_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20473\,
            in3 => \N__20470\,
            lcout => \b2v_inst200.un25_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_6_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22324\,
            lcout => \b2v_inst200.count_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36642\,
            ce => \N__25158\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_8_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20440\,
            lcout => \b2v_inst200.count_3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36642\,
            ce => \N__25158\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_0_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20416\,
            in1 => \N__20425\,
            in2 => \_gnd_net_\,
            in3 => \N__25203\,
            lcout => \b2v_inst200.countZ0Z_0\,
            ltout => \b2v_inst200.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_0_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__22322\,
            in1 => \_gnd_net_\,
            in2 => \N__20419\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36642\,
            ce => \N__25158\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_16_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22323\,
            in2 => \_gnd_net_\,
            in3 => \N__20497\,
            lcout => \b2v_inst200.count_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36642\,
            ce => \N__25158\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_9_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25257\,
            in2 => \_gnd_net_\,
            in3 => \N__20410\,
            lcout => \b2v_inst200.un25_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI50P71_13_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20653\,
            in1 => \N__25216\,
            in2 => \_gnd_net_\,
            in3 => \N__20643\,
            lcout => \b2v_inst200.countZ0Z_13\,
            ltout => \b2v_inst200.countZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_1_0_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20521\,
            in1 => \N__20563\,
            in2 => \N__20626\,
            in3 => \N__20623\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_3_0_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__20611\,
            in1 => \N__20590\,
            in2 => \N__20572\,
            in3 => \N__20569\,
            lcout => \b2v_inst200.un25_clk_100khz_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_14_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20536\,
            lcout => \b2v_inst200.count_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36636\,
            ce => \N__25156\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI96R71_15_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20550\,
            in1 => \N__20542\,
            in2 => \_gnd_net_\,
            in3 => \N__25218\,
            lcout => \b2v_inst200.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_15_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20551\,
            lcout => \b2v_inst200.count_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36636\,
            ce => \N__25156\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI73Q71_14_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20535\,
            in1 => \N__20527\,
            in2 => \_gnd_net_\,
            in3 => \N__25217\,
            lcout => \b2v_inst200.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIB9S71_16_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__25215\,
            in1 => \N__20509\,
            in2 => \N__20496\,
            in3 => \N__22310\,
            lcout => \b2v_inst200.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_11_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22312\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21097\,
            lcout => \b2v_inst200.count_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36630\,
            ce => \N__25155\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_10_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21012\,
            in2 => \_gnd_net_\,
            in3 => \N__22311\,
            lcout => \b2v_inst200.count_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36630\,
            ce => \N__25155\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI1QM71_11_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__22309\,
            in1 => \N__21096\,
            in2 => \N__21088\,
            in3 => \N__25214\,
            lcout => \b2v_inst200.countZ0Z_11\,
            ltout => \b2v_inst200.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_17_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20994\,
            in1 => \N__21072\,
            in2 => \N__21061\,
            in3 => \N__21058\,
            lcout => OPEN,
            ltout => \b2v_inst200.un25_clk_100khz_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIC03N_6_0_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21046\,
            in1 => \N__21037\,
            in2 => \N__21025\,
            in3 => \N__21022\,
            lcout => \b2v_inst200.count_RNIC03N_6Z0Z_0\,
            ltout => \b2v_inst200.count_RNIC03N_6Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNI_0_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21016\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst200.count_RNI_0_0\,
            ltout => \b2v_inst200.count_RNI_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIOMPC1_10_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__21013\,
            in1 => \N__21004\,
            in2 => \N__20998\,
            in3 => \N__25213\,
            lcout => \b2v_inst200.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.count_12_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20980\,
            lcout => \b2v_inst16.count_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36626\,
            ce => \N__20950\,
            sr => \N__20800\
        );

    \b2v_inst11.dutycycle_RNI_1_2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30287\,
            in2 => \_gnd_net_\,
            in3 => \N__21280\,
            lcout => \b2v_inst11.N_366\,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25444\,
            in2 => \N__21242\,
            in3 => \N__21262\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_2_c\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28249\,
            in2 => \N__21244\,
            in3 => \N__21259\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_3_c\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28231\,
            in2 => \N__32519\,
            in3 => \N__21256\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_4_c\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28210\,
            in2 => \N__32520\,
            in3 => \N__21253\,
            lcout => \b2v_inst11.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_5_c\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31706\,
            in1 => \N__28192\,
            in2 => \N__21243\,
            in3 => \N__21250\,
            lcout => \b2v_inst11.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un152_sum_cry_6_c\,
            carryout => \b2v_inst11.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28408\,
            in2 => \_gnd_net_\,
            in3 => \N__21247\,
            lcout => \b2v_inst11.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21220\,
            in2 => \_gnd_net_\,
            in3 => \N__21200\,
            lcout => \b2v_inst16.N_208_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__26777\,
            in1 => \N__21378\,
            in2 => \N__21118\,
            in3 => \N__26647\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_10_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26326\,
            in2 => \_gnd_net_\,
            in3 => \N__29216\,
            lcout => OPEN,
            ltout => \b2v_inst11.un2_count_clk_17_0_a2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_15_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__28895\,
            in1 => \N__21334\,
            in2 => \N__21328\,
            in3 => \N__29612\,
            lcout => \b2v_inst11.N_363\,
            ltout => \b2v_inst11.N_363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_15_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21297\,
            in2 => \N__21283\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_365\,
            ltout => \b2v_inst11.N_365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__33613\,
            in1 => \N__26179\,
            in2 => \N__21274\,
            in3 => \N__33352\,
            lcout => \b2v_inst11.N_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__24365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24155\,
            lcout => \N_161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_6_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101110111"
        )
    port map (
            in0 => \N__26776\,
            in1 => \N__29534\,
            in2 => \_gnd_net_\,
            in3 => \N__26178\,
            lcout => \b2v_inst11.g0_13_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_11_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__29102\,
            in1 => \N__26301\,
            in2 => \N__21439\,
            in3 => \N__26800\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_8_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101011111"
        )
    port map (
            in0 => \N__26299\,
            in1 => \N__29498\,
            in2 => \N__26832\,
            in3 => \N__26183\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_3_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100000"
        )
    port map (
            in0 => \N__28755\,
            in1 => \N__26798\,
            in2 => \N__29532\,
            in3 => \N__26300\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_8_3_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110111"
        )
    port map (
            in0 => \N__26445\,
            in1 => \N__29499\,
            in2 => \N__26327\,
            in3 => \N__28754\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_30_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_9_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010001010"
        )
    port map (
            in0 => \N__26184\,
            in1 => \N__26799\,
            in2 => \N__21442\,
            in3 => \N__26446\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_13_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111111111"
        )
    port map (
            in0 => \N__28896\,
            in1 => \N__29198\,
            in2 => \N__21413\,
            in3 => \N__29037\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_9_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__21430\,
            in1 => \N__26447\,
            in2 => \N__21424\,
            in3 => \N__21406\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_11_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29101\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_7_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__33360\,
            in1 => \N__33621\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.dutycycle_RNI_7Z0Z_1\,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33359\,
            in2 => \N__27132\,
            in3 => \N__21349\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27108\,
            in2 => \N__30278\,
            in3 => \N__21346\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27059\,
            in2 => \N__28757\,
            in3 => \N__21337\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_2\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29509\,
            in2 => \N__27104\,
            in3 => \N__21511\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_3\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27054\,
            in2 => \N__29389\,
            in3 => \N__21499\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_4_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26157\,
            in2 => \N__27103\,
            in3 => \N__21484\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27058\,
            in2 => \N__26842\,
            in3 => \N__21469\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27088\,
            in2 => \N__26336\,
            in3 => \N__21466\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49\,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26438\,
            in2 => \N__27129\,
            in3 => \N__21463\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_8_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27092\,
            in2 => \N__29215\,
            in3 => \N__21460\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_9\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_10_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29115\,
            in2 => \N__27130\,
            in3 => \N__21448\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_10_cZ0\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27096\,
            in2 => \N__29046\,
            in3 => \N__21445\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_11\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28899\,
            in2 => \N__27131\,
            in3 => \N__21574\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_12\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27100\,
            in2 => \N__29725\,
            in3 => \N__21571\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_94_cry_13\,
            carryout => \b2v_inst11.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__27101\,
            in1 => \N__29608\,
            in2 => \_gnd_net_\,
            in3 => \N__21568\,
            lcout => \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_4_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__21556\,
            in1 => \N__23053\,
            in2 => \N__21550\,
            in3 => \N__21523\,
            lcout => \b2v_inst11.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36606\,
            ce => 'H',
            sr => \N__25972\
        );

    \b2v_inst11.dutycycle_RNIP7P13_4_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__27710\,
            in1 => \N__25811\,
            in2 => \N__21549\,
            in3 => \N__21565\,
            lcout => \b2v_inst11.dutycycle_RNIP7P13Z0Z_4\,
            ltout => \b2v_inst11.dutycycle_RNIP7P13Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIKF34B_4_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__21545\,
            in1 => \N__23051\,
            in2 => \N__21529\,
            in3 => \N__21522\,
            lcout => \b2v_inst11.dutycycleZ0Z_7\,
            ltout => \b2v_inst11.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_4_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__23167\,
            in1 => \N__23259\,
            in2 => \N__21526\,
            in3 => \N__23232\,
            lcout => \b2v_inst11.dutycycle_e_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_15_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000011"
        )
    port map (
            in0 => \N__23233\,
            in1 => \N__26648\,
            in2 => \N__25853\,
            in3 => \N__29613\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_158_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIMBHI8_15_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__23052\,
            in1 => \N__23175\,
            in2 => \N__21514\,
            in3 => \N__27664\,
            lcout => \b2v_inst11.dutycycle_en_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__21691\,
            in1 => \N__21699\,
            in2 => \N__27700\,
            in3 => \N__21712\,
            lcout => \b2v_inst11.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36606\,
            ce => 'H',
            sr => \N__25972\
        );

    \b2v_inst11.dutycycle_RNIQGT7G_6_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__21711\,
            in1 => \N__27663\,
            in2 => \N__21703\,
            in3 => \N__21690\,
            lcout => \b2v_inst11.dutycycleZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNIMJCJ5_1_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24637\,
            in2 => \N__33754\,
            in3 => \N__21790\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8E1K7_1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110111111"
        )
    port map (
            in0 => \N__21676\,
            in1 => \N__24125\,
            in2 => \N__21646\,
            in3 => \N__33729\,
            lcout => \b2v_inst11.N_117_f0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIVS8U1_6_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111111"
        )
    port map (
            in0 => \N__21643\,
            in1 => \N__25824\,
            in2 => \N__21877\,
            in3 => \N__23391\,
            lcout => \b2v_inst11.N_5572_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_12_1_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__21613\,
            in1 => \_gnd_net_\,
            in2 => \N__23395\,
            in3 => \N__21875\,
            lcout => OPEN,
            ltout => \b2v_inst11_g0_i_m2_i_a6_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S3n_ibuf_RNI4G1E7_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__21580\,
            in1 => \N__25823\,
            in2 => \N__21631\,
            in3 => \N__21628\,
            lcout => \N_15_i_0_a4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_5_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001100110"
        )
    port map (
            in0 => \N__21612\,
            in1 => \N__21874\,
            in2 => \_gnd_net_\,
            in3 => \N__29330\,
            lcout => OPEN,
            ltout => \b2v_inst11.g0_i_m2_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIS1UT1_5_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101001000000"
        )
    port map (
            in0 => \N__21870\,
            in1 => \N__21589\,
            in2 => \N__21583\,
            in3 => \N__26876\,
            lcout => \N_15_i_0_a4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI4C1Q3_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010001"
        )
    port map (
            in0 => \N__21883\,
            in1 => \N__21876\,
            in2 => \N__21832\,
            in3 => \N__21812\,
            lcout => \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_0_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__21778\,
            in1 => \N__27659\,
            in2 => \N__21769\,
            in3 => \N__21784\,
            lcout => \b2v_inst11.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36620\,
            ce => 'H',
            sr => \N__25897\
        );

    \b2v_inst11.dutycycle_RNI8I5HB_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111011"
        )
    port map (
            in0 => \N__33587\,
            in1 => \N__23026\,
            in2 => \N__33780\,
            in3 => \N__21751\,
            lcout => \b2v_inst11.dutycycle_eena\,
            ltout => \b2v_inst11.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIG4U9E_0_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__21777\,
            in1 => \N__21765\,
            in2 => \N__21754\,
            in3 => \N__27658\,
            lcout => \b2v_inst11.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI8I5HB_1_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111011"
        )
    port map (
            in0 => \N__33755\,
            in1 => \N__23025\,
            in2 => \N__33354\,
            in3 => \N__21750\,
            lcout => \b2v_inst11.dutycycle_eena_0\,
            ltout => \b2v_inst11.dutycycle_eena_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIRGRIE_1_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__21735\,
            in1 => \N__21720\,
            in2 => \N__21742\,
            in3 => \N__27657\,
            lcout => \b2v_inst11.dutycycle\,
            ltout => \b2v_inst11.dutycycle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_1_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__33588\,
            in1 => \_gnd_net_\,
            in2 => \N__21739\,
            in3 => \N__29537\,
            lcout => \b2v_inst11.dutycycle_RNI_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_1_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__21736\,
            in1 => \N__21727\,
            in2 => \N__27714\,
            in3 => \N__21721\,
            lcout => \b2v_inst11.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36620\,
            ce => 'H',
            sr => \N__25897\
        );

    \b2v_inst11.dutycycle_RNI_1_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33586\,
            in1 => \N__29538\,
            in2 => \_gnd_net_\,
            in3 => \N__33320\,
            lcout => \b2v_inst11.g3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI_1_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25569\,
            lcout => \b2v_inst5.curr_state_RNIZ0Z_1\,
            ltout => \b2v_inst5.curr_state_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIR6ES_0_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__34721\,
            in1 => \_gnd_net_\,
            in2 => \N__22123\,
            in3 => \N__21925\,
            lcout => \b2v_inst5_RSMRSTn_latmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_fast_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21928\,
            in1 => \N__34716\,
            in2 => \_gnd_net_\,
            in3 => \N__21904\,
            lcout => \b2v_inst5_RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36625\,
            ce => \N__36361\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21903\,
            in1 => \N__34712\,
            in2 => \_gnd_net_\,
            in3 => \N__21927\,
            lcout => \RSMRSTn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36625\,
            ce => \N__36361\,
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIFLPH1_1_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__21946\,
            in1 => \N__21901\,
            in2 => \N__34722\,
            in3 => \N__36403\,
            lcout => \b2v_inst5.curr_state_RNIFLPH1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNIJJOV_1_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21900\,
            in1 => \N__21945\,
            in2 => \N__34723\,
            in3 => \N__35745\,
            lcout => \b2v_inst5.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m6_i_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__21926\,
            in1 => \N__21902\,
            in2 => \N__25555\,
            in3 => \N__34717\,
            lcout => \b2v_inst5.N_51\,
            ltout => \b2v_inst5.N_51_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_RNI2DVE1_1_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35744\,
            in2 => \N__21886\,
            in3 => \N__30454\,
            lcout => \b2v_inst5.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI2DIN_9_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35813\,
            in1 => \N__22150\,
            in2 => \_gnd_net_\,
            in3 => \N__24669\,
            lcout => \b2v_inst11.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_9_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24673\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36629\,
            ce => \N__36358\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIB49T_10_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22144\,
            in2 => \N__24658\,
            in3 => \N__35811\,
            lcout => \b2v_inst11.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_10_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24657\,
            lcout => \b2v_inst11.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36629\,
            ce => \N__36358\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIK61M_11_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35812\,
            in1 => \N__22138\,
            in2 => \_gnd_net_\,
            in3 => \N__24783\,
            lcout => \b2v_inst11.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_11_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24787\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36629\,
            ce => \N__36358\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIKNAN_2_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22132\,
            in2 => \N__24721\,
            in3 => \N__35810\,
            lcout => \b2v_inst11.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_2_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24720\,
            lcout => \b2v_inst11.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36629\,
            ce => \N__36358\,
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m8_i_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__22206\,
            in1 => \N__22192\,
            in2 => \N__22600\,
            in3 => \N__33684\,
            lcout => OPEN,
            ltout => \b2v_inst200.N_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNICM0V7_1_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22162\,
            in2 => \N__22126\,
            in3 => \N__35775\,
            lcout => \b2v_inst200.curr_stateZ0Z_1\,
            ltout => \b2v_inst200.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22333\,
            in3 => \N__22227\,
            lcout => \N_411\,
            ltout => \N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__22330\,
            in1 => \N__22264\,
            in2 => \N__22252\,
            in3 => \N__22207\,
            lcout => \b2v_inst200.m6_i_0\,
            ltout => \b2v_inst200.m6_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m6_i_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111001"
        )
    port map (
            in0 => \N__22194\,
            in1 => \N__22228\,
            in2 => \N__22243\,
            in3 => \N__33683\,
            lcout => OPEN,
            ltout => \b2v_inst200.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_RNIGPR58_0_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22240\,
            in2 => \N__22234\,
            in3 => \N__35774\,
            lcout => \b2v_inst200.curr_stateZ0Z_0\,
            ltout => \b2v_inst200.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m8_i_a3_0_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22191\,
            in2 => \N__22210\,
            in3 => \_gnd_net_\,
            lcout => \N_412\,
            ltout => \N_412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_1_LC_6_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__33685\,
            in1 => \N__22596\,
            in2 => \N__22198\,
            in3 => \N__22193\,
            lcout => \b2v_inst200.curr_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36635\,
            ce => \N__36356\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_4_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27834\,
            in1 => \N__27802\,
            in2 => \N__27996\,
            in3 => \N__27762\,
            lcout => \b2v_inst36.un12_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNINEG01_6_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22156\,
            in1 => \N__30696\,
            in2 => \_gnd_net_\,
            in3 => \N__27786\,
            lcout => \b2v_inst36.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_6_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27787\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36650\,
            ce => \N__30699\,
            sr => \N__30591\
        );

    \b2v_inst36.count_RNIHJCV_12_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22360\,
            in1 => \N__30698\,
            in2 => \_gnd_net_\,
            in3 => \N__27975\,
            lcout => \b2v_inst36.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIJ8E01_4_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27819\,
            in1 => \N__22372\,
            in2 => \_gnd_net_\,
            in3 => \N__30695\,
            lcout => \b2v_inst36.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_4_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27820\,
            lcout => \b2v_inst36.count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36650\,
            ce => \N__30699\,
            sr => \N__30591\
        );

    \b2v_inst36.count_RNITNJ01_9_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22366\,
            in1 => \N__30697\,
            in2 => \_gnd_net_\,
            in3 => \N__27747\,
            lcout => \b2v_inst36.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_14_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27934\,
            lcout => \b2v_inst36.count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36644\,
            ce => \N__30732\,
            sr => \N__30587\
        );

    \b2v_inst36.count_9_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27748\,
            lcout => \b2v_inst36.count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36644\,
            ce => \N__30732\,
            sr => \N__30587\
        );

    \b2v_inst36.count_12_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36644\,
            ce => \N__30732\,
            sr => \N__30587\
        );

    \b2v_inst36.curr_state_RNI8TT2_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__22398\,
            in1 => \_gnd_net_\,
            in2 => \N__25354\,
            in3 => \N__25289\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_RNI8TT2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_RNIUDI9_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22414\,
            in1 => \_gnd_net_\,
            in2 => \N__22354\,
            in3 => \N__35933\,
            lcout => \DSW_PWROK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_0_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__30845\,
            in1 => \N__22393\,
            in2 => \N__25352\,
            in3 => \N__25287\,
            lcout => \b2v_inst36.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36638\,
            ce => \N__36367\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.DSW_PWROK_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__25286\,
            in1 => \_gnd_net_\,
            in2 => \N__22399\,
            in3 => \N__25340\,
            lcout => \b2v_inst36.DSW_PWROK_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36638\,
            ce => \N__36367\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m4_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011000000"
        )
    port map (
            in0 => \N__30844\,
            in1 => \N__22397\,
            in2 => \N__25353\,
            in3 => \N__25285\,
            lcout => OPEN,
            ltout => \b2v_inst36.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI2MTL_0_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22408\,
            in2 => \N__22402\,
            in3 => \N__35932\,
            lcout => \b2v_inst36.curr_stateZ0Z_0\,
            ltout => \b2v_inst36.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI_0_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22378\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.N_2939_i\,
            ltout => \b2v_inst36.N_2939_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_7_1_0__m6_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011100000"
        )
    port map (
            in0 => \N__25288\,
            in1 => \N__25347\,
            in2 => \N__22375\,
            in3 => \N__30843\,
            lcout => \b2v_inst36.curr_state_7_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_11_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31444\,
            lcout => \b2v_inst5.count_1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36631\,
            ce => \N__31928\,
            sr => \N__32173\
        );

    \b2v_inst5.count_12_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31411\,
            lcout => \b2v_inst5.count_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36631\,
            ce => \N__31928\,
            sr => \N__32173\
        );

    \b2v_inst5.count_14_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31324\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36631\,
            ce => \N__31928\,
            sr => \N__32173\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28657\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25450\,
            in2 => \N__22507\,
            in3 => \N__22444\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22671\,
            in2 => \N__22660\,
            in3 => \N__22441\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32548\,
            in2 => \N__22558\,
            in3 => \N__22438\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22546\,
            in2 => \N__32556\,
            in3 => \N__22435\,
            lcout => \b2v_inst11.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25474\,
            in1 => \N__22536\,
            in2 => \N__22426\,
            in3 => \N__22432\,
            lcout => \b2v_inst11.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un131_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22525\,
            in3 => \N__22429\,
            lcout => \b2v_inst11.mult1_un131_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22537\,
            in2 => \_gnd_net_\,
            in3 => \N__32547\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28626\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25495\,
            in2 => \N__25593\,
            in3 => \N__22417\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25589\,
            in2 => \N__25435\,
            in3 => \N__22549\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25642\,
            in2 => \N__32586\,
            in3 => \N__22540\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32582\,
            in2 => \N__25633\,
            in3 => \N__22528\,
            lcout => \b2v_inst11.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32552\,
            in1 => \N__25621\,
            in2 => \N__25594\,
            in3 => \N__22516\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un124_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25612\,
            in3 => \N__22513\,
            lcout => \b2v_inst11.mult1_un124_sum_s_8\,
            ltout => \b2v_inst11.mult1_un124_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22510\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIPFFQ6_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110011"
        )
    port map (
            in0 => \N__22497\,
            in1 => \N__23067\,
            in2 => \N__22456\,
            in3 => \N__27147\,
            lcout => b2v_inst11_dutycycle_set_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28677\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_14_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22686\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__22672\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32546\,
            lcout => \b2v_inst11.mult1_un131_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_9_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100011101010"
        )
    port map (
            in0 => \N__26335\,
            in1 => \N__26449\,
            in2 => \N__26823\,
            in3 => \N__22648\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_13_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26450\,
            in1 => \N__28900\,
            in2 => \N__22642\,
            in3 => \N__29223\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22639\,
            in2 => \_gnd_net_\,
            in3 => \N__22627\,
            lcout => \b2v_inst200.m11_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_3_c_RNIB6L91_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__31491\,
            in1 => \N__31131\,
            in2 => \N__31152\,
            in3 => \N__32094\,
            lcout => \b2v_inst5.count_rst_10\,
            ltout => \b2v_inst5.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIP7CS2_4_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__31835\,
            in1 => \_gnd_net_\,
            in2 => \N__22570\,
            in3 => \N__22770\,
            lcout => \b2v_inst5.un2_count_1_axb_4\,
            ltout => \b2v_inst5.un2_count_1_axb_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_4_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__31492\,
            in1 => \N__31132\,
            in2 => \N__22567\,
            in3 => \N__32096\,
            lcout => \b2v_inst5.count_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36608\,
            ce => \N__31941\,
            sr => \N__32135\
        );

    \b2v_inst5.count_8_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__32095\,
            in1 => \N__31493\,
            in2 => \N__31066\,
            in3 => \N__31085\,
            lcout => \b2v_inst5.count_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36608\,
            ce => \N__31941\,
            sr => \N__32135\
        );

    \b2v_inst5.count_RNI1KGS2_8_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__22564\,
            in1 => \N__31836\,
            in2 => \_gnd_net_\,
            in3 => \N__28282\,
            lcout => \b2v_inst5.countZ0Z_8\,
            ltout => \b2v_inst5.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIP7CS2_0_4_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__31942\,
            in1 => \N__22780\,
            in2 => \N__22774\,
            in3 => \N__22771\,
            lcout => OPEN,
            ltout => \b2v_inst5.un12_clk_100khz_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIAEONB_2_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28294\,
            in1 => \N__28048\,
            in2 => \N__22762\,
            in3 => \N__31615\,
            lcout => \b2v_inst5.un12_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_9_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__29491\,
            in1 => \N__26425\,
            in2 => \N__26836\,
            in3 => \N__26155\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_10_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__26308\,
            in1 => \N__26435\,
            in2 => \N__22759\,
            in3 => \N__29199\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_10_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010101001010"
        )
    port map (
            in0 => \N__29200\,
            in1 => \N__22756\,
            in2 => \N__22744\,
            in3 => \N__22693\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNITS10B_14_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__22737\,
            in1 => \N__22726\,
            in2 => \N__22717\,
            in3 => \N__25864\,
            lcout => \b2v_inst11.dutycycleZ0Z_12\,
            ltout => \b2v_inst11.dutycycleZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_11_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22696\,
            in3 => \N__29116\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_6_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__26153\,
            in1 => \N__29490\,
            in2 => \_gnd_net_\,
            in3 => \N__26808\,
            lcout => \b2v_inst11.N_15_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_9_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26426\,
            in2 => \N__29530\,
            in3 => \N__26154\,
            lcout => \b2v_inst11.dutycycle_RNI_3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_9_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26156\,
            in1 => \N__26436\,
            in2 => \N__29397\,
            in3 => \N__22849\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI5K4VA_9_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__25836\,
            in1 => \N__22809\,
            in2 => \N__22828\,
            in3 => \N__22834\,
            lcout => \b2v_inst11.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIRP00B_13_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__23271\,
            in1 => \N__22788\,
            in2 => \N__22801\,
            in3 => \N__25837\,
            lcout => \b2v_inst11.dutycycleZ0Z_8\,
            ltout => \b2v_inst11.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_13_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010101"
        )
    port map (
            in0 => \N__25835\,
            in1 => \N__23242\,
            in2 => \N__22843\,
            in3 => \N__26570\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_153_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIMBHI8_13_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__27671\,
            in1 => \N__23181\,
            in2 => \N__22840\,
            in3 => \N__23066\,
            lcout => \b2v_inst11.dutycycle_en_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_9_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010101"
        )
    port map (
            in0 => \N__25834\,
            in1 => \N__23241\,
            in2 => \N__26451\,
            in3 => \N__26569\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_156_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIMBHI8_9_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__27670\,
            in1 => \N__23180\,
            in2 => \N__22837\,
            in3 => \N__23065\,
            lcout => \b2v_inst11.dutycycle_e_1_9\,
            ltout => \b2v_inst11.dutycycle_e_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__25838\,
            in1 => \N__22824\,
            in2 => \N__22813\,
            in3 => \N__22810\,
            lcout => \b2v_inst11.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36607\,
            ce => 'H',
            sr => \N__25946\
        );

    \b2v_inst11.dutycycle_13_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__22797\,
            in1 => \N__22789\,
            in2 => \N__23275\,
            in3 => \N__25839\,
            lcout => \b2v_inst11.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36607\,
            ce => 'H',
            sr => \N__25946\
        );

    \b2v_inst11.dutycycle_RNI0084B_8_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__23055\,
            in1 => \N__22880\,
            in2 => \N__22861\,
            in3 => \N__23076\,
            lcout => \b2v_inst11.dutycycleZ0Z_5\,
            ltout => \b2v_inst11.dutycycleZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_8_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__23234\,
            in1 => \N__23173\,
            in2 => \N__23263\,
            in3 => \N__23260\,
            lcout => \b2v_inst11.dutycycle_e_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNICDJJ5_10_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010101"
        )
    port map (
            in0 => \N__25860\,
            in1 => \N__23235\,
            in2 => \N__29217\,
            in3 => \N__26643\,
            lcout => OPEN,
            ltout => \b2v_inst11.N_154_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIMBHI8_10_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101010"
        )
    port map (
            in0 => \N__27672\,
            in1 => \N__23174\,
            in2 => \N__23083\,
            in3 => \N__23054\,
            lcout => \b2v_inst11.dutycycle_en_4\,
            ltout => \b2v_inst11.dutycycle_en_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIEOB3B_10_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__25861\,
            in1 => \N__22896\,
            in2 => \N__23080\,
            in3 => \N__22909\,
            lcout => \b2v_inst11.dutycycleZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_8_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__23077\,
            in1 => \N__22857\,
            in2 => \N__22885\,
            in3 => \N__23056\,
            lcout => \b2v_inst11.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36613\,
            ce => 'H',
            sr => \N__25980\
        );

    \b2v_inst11.dutycycle_10_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__25863\,
            in1 => \N__22915\,
            in2 => \N__22900\,
            in3 => \N__22908\,
            lcout => \b2v_inst11.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36613\,
            ce => 'H',
            sr => \N__25980\
        );

    \b2v_inst11.dutycycle_RNI1KT13_8_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__22881\,
            in1 => \N__22870\,
            in2 => \N__27701\,
            in3 => \N__25862\,
            lcout => \b2v_inst11.dutycycle_RNI1KT13Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI8JP5_0_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__23389\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24638\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI6P011_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__24514\,
            in1 => \N__24931\,
            in2 => \N__24400\,
            in3 => \N__23672\,
            lcout => \b2v_inst11.N_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIU8G3G_2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__23919\,
            in1 => \N__27668\,
            in2 => \N__23947\,
            in3 => \N__23934\,
            lcout => \dutycycle_RNIU8G3G_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIF6NL_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111110101010"
        )
    port map (
            in0 => \N__24370\,
            in1 => \N__24226\,
            in2 => \N__24217\,
            in3 => \N__24126\,
            lcout => OPEN,
            ltout => \b2v_inst11.g1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.func_state_RNI5M9V2_1_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__23876\,
            in1 => \_gnd_net_\,
            in2 => \N__23956\,
            in3 => \N__23953\,
            lcout => \b2v_inst11.g1\,
            ltout => \b2v_inst11.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_2_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__23920\,
            in1 => \N__27669\,
            in2 => \N__23938\,
            in3 => \N__23935\,
            lcout => \b2v_inst11.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36621\,
            ce => 'H',
            sr => \N__25945\
        );

    \b2v_inst5.RSMRSTn_fast_RNIVS8U1_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__23875\,
            in1 => \N__23671\,
            in2 => \N__23531\,
            in3 => \N__23388\,
            lcout => \b2v_inst5.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32439\,
            in2 => \N__32400\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \b2v_inst11.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27448\,
            in1 => \N__32357\,
            in2 => \_gnd_net_\,
            in3 => \N__24706\,
            lcout => \b2v_inst11.count_1_2\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_1\,
            carryout => \b2v_inst11.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27452\,
            in1 => \N__32306\,
            in2 => \_gnd_net_\,
            in3 => \N__24703\,
            lcout => \b2v_inst11.count_1_3\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_2\,
            carryout => \b2v_inst11.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27449\,
            in1 => \N__32940\,
            in2 => \_gnd_net_\,
            in3 => \N__24700\,
            lcout => \b2v_inst11.count_1_4\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_3\,
            carryout => \b2v_inst11.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27453\,
            in1 => \N__32901\,
            in2 => \_gnd_net_\,
            in3 => \N__24697\,
            lcout => \b2v_inst11.count_1_5\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_4\,
            carryout => \b2v_inst11.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27450\,
            in1 => \N__32847\,
            in2 => \_gnd_net_\,
            in3 => \N__24694\,
            lcout => \b2v_inst11.count_1_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_5\,
            carryout => \b2v_inst11.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27454\,
            in1 => \N__32804\,
            in2 => \_gnd_net_\,
            in3 => \N__24679\,
            lcout => \b2v_inst11.count_1_7\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_6\,
            carryout => \b2v_inst11.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27451\,
            in1 => \N__32766\,
            in2 => \_gnd_net_\,
            in3 => \N__24676\,
            lcout => \b2v_inst11.count_1_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_7\,
            carryout => \b2v_inst11.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27438\,
            in1 => \N__32711\,
            in2 => \_gnd_net_\,
            in3 => \N__24661\,
            lcout => \b2v_inst11.count_1_9\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \b2v_inst11.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27455\,
            in1 => \N__32657\,
            in2 => \_gnd_net_\,
            in3 => \N__24646\,
            lcout => \b2v_inst11.count_1_10\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_9\,
            carryout => \b2v_inst11.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27437\,
            in1 => \N__32615\,
            in2 => \_gnd_net_\,
            in3 => \N__24775\,
            lcout => \b2v_inst11.count_1_11\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_10\,
            carryout => \b2v_inst11.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27456\,
            in1 => \N__33120\,
            in2 => \_gnd_net_\,
            in3 => \N__24772\,
            lcout => \b2v_inst11.count_1_12\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_11\,
            carryout => \b2v_inst11.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27439\,
            in1 => \N__33087\,
            in2 => \_gnd_net_\,
            in3 => \N__24769\,
            lcout => \b2v_inst11.count_1_13\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_12\,
            carryout => \b2v_inst11.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27457\,
            in1 => \N__33051\,
            in2 => \_gnd_net_\,
            in3 => \N__24766\,
            lcout => \b2v_inst11.count_1_14\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_count_cry_13\,
            carryout => \b2v_inst11.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__27440\,
            in1 => \N__33018\,
            in2 => \_gnd_net_\,
            in3 => \N__24763\,
            lcout => \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQF4M_14_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35901\,
            in1 => \N__24727\,
            in2 => \_gnd_net_\,
            in3 => \N__24738\,
            lcout => \b2v_inst11.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIQ0EN_5_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35886\,
            in1 => \N__24745\,
            in2 => \_gnd_net_\,
            in3 => \N__24756\,
            lcout => \b2v_inst11.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_5_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24760\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36637\,
            ce => \N__36355\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_14_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24739\,
            lcout => \b2v_inst11.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36637\,
            ce => \N__36355\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIS3FN_6_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35885\,
            in1 => \N__24973\,
            in2 => \_gnd_net_\,
            in3 => \N__24984\,
            lcout => \b2v_inst11.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_6_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24988\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36637\,
            ce => \N__36355\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNISI5M_15_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24955\,
            in1 => \N__35870\,
            in2 => \_gnd_net_\,
            in3 => \N__24963\,
            lcout => \b2v_inst11.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_15_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24967\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36637\,
            ce => \N__36355\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__36409\,
            in1 => \N__24940\,
            in2 => \N__32989\,
            in3 => \N__29877\,
            lcout => OPEN,
            ltout => \b2v_inst11.pwm_out_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNIEV5S_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__29876\,
            in1 => \_gnd_net_\,
            in2 => \N__24949\,
            in3 => \N__27484\,
            lcout => \PWRBTN_LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst20.tmp_1_rep1_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24901\,
            in2 => \_gnd_net_\,
            in3 => \N__24836\,
            lcout => \SYNTHESIZED_WIRE_1keep_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35917\,
            in1 => \N__29875\,
            in2 => \_gnd_net_\,
            in3 => \N__29838\,
            lcout => \b2v_inst11.pwm_out_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.G_146_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24900\,
            in2 => \_gnd_net_\,
            in3 => \N__24835\,
            lcout => \G_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_0_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__27349\,
            in1 => \N__30959\,
            in2 => \_gnd_net_\,
            in3 => \N__30842\,
            lcout => \b2v_inst36.count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36657\,
            ce => \N__30700\,
            sr => \N__30590\
        );

    \b2v_inst36.count_RNI471O_1_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25009\,
            in1 => \N__25021\,
            in2 => \_gnd_net_\,
            in3 => \N__30701\,
            lcout => OPEN,
            ltout => \b2v_inst36.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI471O_2_1_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__28027\,
            in1 => \N__27904\,
            in2 => \N__25045\,
            in3 => \N__28150\,
            lcout => OPEN,
            ltout => \b2v_inst36.un12_clk_100khz_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNISMPL1_1_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25000\,
            in1 => \N__25042\,
            in2 => \N__25033\,
            in3 => \N__30382\,
            lcout => \b2v_inst36.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI361O_0_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25030\,
            in1 => \N__24994\,
            in2 => \_gnd_net_\,
            in3 => \N__30693\,
            lcout => \b2v_inst36.countZ0Z_0\,
            ltout => \b2v_inst36.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_1_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__30957\,
            in1 => \_gnd_net_\,
            in2 => \N__25024\,
            in3 => \N__27364\,
            lcout => \b2v_inst36.count_rst_13\,
            ltout => \b2v_inst36.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI471O_0_1_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25008\,
            in2 => \N__25015\,
            in3 => \N__30694\,
            lcout => \b2v_inst36.un2_count_1_axb_1\,
            ltout => \b2v_inst36.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_1_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__30958\,
            in1 => \_gnd_net_\,
            in2 => \N__25012\,
            in3 => \N__27348\,
            lcout => \b2v_inst36.count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36657\,
            ce => \N__30700\,
            sr => \N__30590\
        );

    \b2v_inst36.count_RNIOFOT_0_14_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28060\,
            in1 => \N__27350\,
            in2 => \N__27952\,
            in3 => \N__28108\,
            lcout => \b2v_inst36.un12_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_0_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__27351\,
            in1 => \N__30912\,
            in2 => \_gnd_net_\,
            in3 => \N__30811\,
            lcout => \b2v_inst36.count_rst_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__30813\,
            in1 => \N__28026\,
            in2 => \N__30956\,
            in3 => \N__28008\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIFGBV_11_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25078\,
            in2 => \N__25084\,
            in3 => \N__30661\,
            lcout => \b2v_inst36.countZ0Z_11\,
            ltout => \b2v_inst36.countZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_11_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010001000000"
        )
    port map (
            in0 => \N__30814\,
            in1 => \N__30927\,
            in2 => \N__25081\,
            in3 => \N__28009\,
            lcout => \b2v_inst36.count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36652\,
            ce => \N__30730\,
            sr => \N__30592\
        );

    \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__27849\,
            in1 => \N__30399\,
            in2 => \N__30960\,
            in3 => \N__30812\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIF2C01_2_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30660\,
            in1 => \_gnd_net_\,
            in2 => \N__25072\,
            in3 => \N__25066\,
            lcout => \b2v_inst36.countZ0Z_2\,
            ltout => \b2v_inst36.countZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_2_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__27850\,
            in1 => \N__30916\,
            in2 => \N__25069\,
            in3 => \N__30815\,
            lcout => \b2v_inst36.count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36652\,
            ce => \N__30730\,
            sr => \N__30592\
        );

    \b2v_inst36.curr_state_RNI3NTL_1_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25051\,
            in1 => \N__25060\,
            in2 => \_gnd_net_\,
            in3 => \N__35930\,
            lcout => \b2v_inst36.curr_stateZ0Z_1\,
            ltout => \b2v_inst36.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNIKEBL_1_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000000000"
        )
    port map (
            in0 => \N__30536\,
            in1 => \N__25365\,
            in2 => \N__25054\,
            in3 => \N__36407\,
            lcout => \b2v_inst36.count_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011100000"
        )
    port map (
            in0 => \N__25291\,
            in1 => \N__25336\,
            in2 => \N__25369\,
            in3 => \N__30856\,
            lcout => \b2v_inst36.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36646\,
            ce => \N__36368\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI0A86_1_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__35931\,
            in1 => \N__25364\,
            in2 => \N__25351\,
            in3 => \N__25290\,
            lcout => \b2v_inst36.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100000"
        )
    port map (
            in0 => \N__31004\,
            in1 => \N__30765\,
            in2 => \N__30980\,
            in3 => \N__30857\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIPHH01_7_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30724\,
            in2 => \N__25264\,
            in3 => \N__30745\,
            lcout => \b2v_inst36.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.curr_state_RNI_1_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30535\,
            lcout => \b2v_inst36.N_2942_i\,
            ltout => \b2v_inst36.N_2942_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__30855\,
            in1 => \N__27903\,
            in2 => \N__25261\,
            in3 => \N__27876\,
            lcout => \b2v_inst36.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_RNIFF751_9_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25240\,
            in1 => \N__25225\,
            in2 => \_gnd_net_\,
            in3 => \N__25202\,
            lcout => \b2v_inst200.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst200.count_9_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25239\,
            lcout => \b2v_inst200.count_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36639\,
            ce => \N__25157\,
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIOFOT_14_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25099\,
            in1 => \N__30680\,
            in2 => \_gnd_net_\,
            in3 => \N__27933\,
            lcout => \b2v_inst36.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIL7E23_11_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31443\,
            in1 => \N__25090\,
            in2 => \_gnd_net_\,
            in3 => \N__31911\,
            lcout => \b2v_inst5.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNINAF23_12_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31912\,
            in1 => \N__25423\,
            in2 => \_gnd_net_\,
            in3 => \N__31410\,
            lcout => \b2v_inst5.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIRGH23_14_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__25414\,
            in1 => \N__31913\,
            in2 => \_gnd_net_\,
            in3 => \N__31323\,
            lcout => \b2v_inst5.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNITJI23_15_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__31914\,
            in1 => \N__31285\,
            in2 => \_gnd_net_\,
            in3 => \N__31267\,
            lcout => \b2v_inst5.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28681\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25489\,
            in2 => \N__25517\,
            in3 => \N__25408\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25405\,
            in2 => \N__25519\,
            in3 => \N__25399\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25396\,
            in2 => \N__25483\,
            in3 => \N__25390\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25387\,
            in2 => \N__25482\,
            in3 => \N__25381\,
            lcout => \b2v_inst11.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32466\,
            in1 => \N__25378\,
            in2 => \N__25518\,
            in3 => \N__25372\,
            lcout => \b2v_inst11.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un138_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25522\,
            lcout => \b2v_inst11.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25475\,
            lcout => \b2v_inst11.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28576\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28656\,
            lcout => \b2v_inst11.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25473\,
            lcout => \b2v_inst11.mult1_un131_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28575\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25675\,
            in2 => \N__28506\,
            in3 => \N__25426\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28502\,
            in2 => \N__28360\,
            in3 => \N__25636\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28348\,
            in2 => \N__31689\,
            in3 => \N__25624\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31685\,
            in2 => \N__28339\,
            in3 => \N__25615\,
            lcout => \b2v_inst11.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32578\,
            in1 => \N__28327\,
            in2 => \N__28507\,
            in3 => \N__25603\,
            lcout => \b2v_inst11.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un117_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28525\,
            in3 => \N__25600\,
            lcout => \b2v_inst11.mult1_un117_sum_s_8\,
            ltout => \b2v_inst11.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25597\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31494\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25576\,
            lcout => \N_413\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29251\,
            lcout => \b2v_inst11.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28830\,
            lcout => \b2v_inst11.mult1_un103_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35213\,
            lcout => \b2v_inst11.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28542\,
            lcout => \b2v_inst11.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI4ALGH_5_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28270\,
            in1 => \N__32203\,
            in2 => \N__31762\,
            in3 => \N__25669\,
            lcout => \b2v_inst5.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_14_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29705\,
            in2 => \_gnd_net_\,
            in3 => \N__25663\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_10_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__26433\,
            in1 => \N__26206\,
            in2 => \N__29027\,
            in3 => \N__29219\,
            lcout => OPEN,
            ltout => \b2v_inst11.i7_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_11_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001110010"
        )
    port map (
            in0 => \N__29128\,
            in1 => \N__26035\,
            in2 => \N__25657\,
            in3 => \N__29000\,
            lcout => \b2v_inst11.dutycycle_RNIZ0Z_11\,
            ltout => \b2v_inst11.dutycycle_RNIZ0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_13_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__29001\,
            in1 => \_gnd_net_\,
            in2 => \N__25654\,
            in3 => \N__28882\,
            lcout => \b2v_inst11.dutycycle_RNI_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_8_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001010110000"
        )
    port map (
            in0 => \N__26333\,
            in1 => \N__25651\,
            in2 => \N__26843\,
            in3 => \N__26189\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26434\,
            in1 => \N__29033\,
            in2 => \N__25645\,
            in3 => \N__26334\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_5_10_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100010001"
        )
    port map (
            in0 => \N__29218\,
            in1 => \N__26432\,
            in2 => \N__26338\,
            in3 => \N__26041\,
            lcout => \b2v_inst11.i6_mux_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_13_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \N__29706\,
            in1 => \N__28881\,
            in2 => \N__29028\,
            in3 => \N__26029\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIC6LA7_12_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__25826\,
            in1 => \N__25989\,
            in2 => \N__26008\,
            in3 => \N__26022\,
            lcout => \b2v_inst11.dutycycleZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_12_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__26023\,
            in1 => \N__26004\,
            in2 => \N__25993\,
            in3 => \N__25830\,
            lcout => \b2v_inst11.dutycycleZ1Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36614\,
            ce => 'H',
            sr => \N__25947\
        );

    \b2v_inst11.dutycycle_15_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__25705\,
            in1 => \N__25719\,
            in2 => \N__25857\,
            in3 => \N__25873\,
            lcout => \b2v_inst11.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36614\,
            ce => 'H',
            sr => \N__25947\
        );

    \b2v_inst11.dutycycle_RNIVV20B_15_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__25872\,
            in1 => \N__25825\,
            in2 => \N__25723\,
            in3 => \N__25704\,
            lcout => \b2v_inst11.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_10_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000001"
        )
    port map (
            in0 => \N__26280\,
            in1 => \N__29190\,
            in2 => \N__26845\,
            in3 => \N__25693\,
            lcout => OPEN,
            ltout => \b2v_inst11.un1_dutycycle_53_50_1_i_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_11_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000010"
        )
    port map (
            in0 => \N__29191\,
            in1 => \N__26356\,
            in2 => \N__25681\,
            in3 => \N__29129\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_11_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29130\,
            in1 => \N__29594\,
            in2 => \N__25678\,
            in3 => \N__29005\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_10_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__29189\,
            in1 => \N__26437\,
            in2 => \N__26309\,
            in3 => \N__26059\,
            lcout => \b2v_inst11.un1_dutycycle_53_50_1_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_3_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__28775\,
            in1 => \N__26350\,
            in2 => \N__28606\,
            in3 => \N__26167\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29390\,
            in2 => \N__29535\,
            in3 => \N__33361\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_1\,
            ltout => \b2v_inst11.dutycycle_RNI_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_0_2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__28774\,
            in1 => \N__30242\,
            in2 => \N__26344\,
            in3 => \N__26166\,
            lcout => \b2v_inst11.dutycycle_RNI_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_3_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010001000"
        )
    port map (
            in0 => \N__29517\,
            in1 => \N__26835\,
            in2 => \_gnd_net_\,
            in3 => \N__28773\,
            lcout => OPEN,
            ltout => \b2v_inst11.dutycycle_RNI_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_8_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__26276\,
            in1 => \N__29392\,
            in2 => \N__26341\,
            in3 => \N__29518\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_8_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__26164\,
            in1 => \N__26275\,
            in2 => \N__29536\,
            in3 => \N__26834\,
            lcout => \b2v_inst11.m6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_2_6_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__26833\,
            in1 => \N__29516\,
            in2 => \_gnd_net_\,
            in3 => \N__26165\,
            lcout => \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_fast_RNIUPHS3_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100011"
        )
    port map (
            in0 => \N__26482\,
            in1 => \N__27187\,
            in2 => \N__27181\,
            in3 => \N__26854\,
            lcout => \N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_12_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__26886\,
            in1 => \N__27199\,
            in2 => \_gnd_net_\,
            in3 => \N__26645\,
            lcout => b2v_inst11_un1_dutycycle_164_0,
            ltout => \b2v_inst11_un1_dutycycle_164_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.RSMRSTn_fast_RNIUPHS3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101101"
        )
    port map (
            in0 => \N__27177\,
            in1 => \N__26481\,
            in2 => \N__27166\,
            in3 => \N__26853\,
            lcout => \b2v_inst5.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28784\,
            in1 => \N__26837\,
            in2 => \_gnd_net_\,
            in3 => \N__29531\,
            lcout => \b2v_inst11.dutycycle_RNI_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_4_1_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__26646\,
            in1 => \N__33629\,
            in2 => \N__27146\,
            in3 => \N__33355\,
            lcout => \b2v_inst11.un1_dutycycle_96_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNIVS8U1_2_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010101110"
        )
    port map (
            in0 => \N__26962\,
            in1 => \N__26943\,
            in2 => \N__26887\,
            in3 => \N__30241\,
            lcout => \N_73_mux_i_i_o3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_3_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28785\,
            in1 => \N__26838\,
            in2 => \N__26665\,
            in3 => \N__26644\,
            lcout => g3_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIM92M_12_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35922\,
            in1 => \N__26458\,
            in2 => \_gnd_net_\,
            in3 => \N__26466\,
            lcout => \b2v_inst11.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_12_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26470\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36632\,
            ce => \N__36362\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIMQBN_3_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27244\,
            in1 => \_gnd_net_\,
            in2 => \N__35934\,
            in3 => \N__27252\,
            lcout => \b2v_inst11.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27256\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36632\,
            ce => \N__36362\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOC3M_13_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35923\,
            in1 => \N__27226\,
            in2 => \_gnd_net_\,
            in3 => \N__27234\,
            lcout => \b2v_inst11.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_13_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27238\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36632\,
            ce => \N__36362\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNIOTCN_4_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__35918\,
            in1 => \N__27208\,
            in2 => \_gnd_net_\,
            in3 => \N__27216\,
            lcout => \b2v_inst11.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_4_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27220\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36632\,
            ce => \N__36362\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNO_0_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__35924\,
            in1 => \N__29878\,
            in2 => \_gnd_net_\,
            in3 => \N__29832\,
            lcout => \b2v_inst11.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__33119\,
            in1 => \N__32625\,
            in2 => \N__32673\,
            in3 => \N__32718\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_5_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__32840\,
            in1 => \N__32894\,
            in2 => \N__27202\,
            in3 => \N__27325\,
            lcout => \b2v_inst11.un79_clk_100khzlto15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_2_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32939\,
            in2 => \N__32310\,
            in3 => \N__32361\,
            lcout => \b2v_inst11.un79_clk_100khzlt6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_15_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32811\,
            in1 => \N__32759\,
            in2 => \_gnd_net_\,
            in3 => \N__33017\,
            lcout => OPEN,
            ltout => \b2v_inst11.un79_clk_100khzlto15_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33050\,
            in1 => \N__33086\,
            in2 => \N__27319\,
            in3 => \N__27316\,
            lcout => \b2v_inst11.count_RNIZ0Z_13\,
            ltout => \b2v_inst11.count_RNIZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_RNO_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__35925\,
            in1 => \N__36408\,
            in2 => \N__27310\,
            in3 => \N__29879\,
            lcout => \b2v_inst11.g0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI03G9_0_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27292\,
            in1 => \N__35859\,
            in2 => \_gnd_net_\,
            in3 => \N__27370\,
            lcout => \b2v_inst11.countZ0Z_0\,
            ltout => \b2v_inst11.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_1_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27420\,
            in2 => \N__27307\,
            in3 => \N__32393\,
            lcout => OPEN,
            ltout => \b2v_inst11.count_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI14G9_1_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27298\,
            in2 => \N__27304\,
            in3 => \N__35860\,
            lcout => \b2v_inst11.countZ0Z_1\,
            ltout => \b2v_inst11.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_1_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__32437\,
            in1 => \_gnd_net_\,
            in2 => \N__27301\,
            in3 => \N__27419\,
            lcout => \b2v_inst11.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36645\,
            ce => \N__36359\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_0_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32436\,
            in2 => \_gnd_net_\,
            in3 => \N__27418\,
            lcout => \b2v_inst11.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36645\,
            ce => \N__36359\,
            sr => \_gnd_net_\
        );

    \SLP_S3n_ibuf_RNIHESTE_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__27286\,
            in1 => \N__27595\,
            in2 => \_gnd_net_\,
            in3 => \N__27553\,
            lcout => \N_73_mux_i_i_a7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI0AHN_8_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27511\,
            in1 => \N__27499\,
            in2 => \_gnd_net_\,
            in3 => \N__35861\,
            lcout => \b2v_inst11.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_8_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27510\,
            lcout => \b2v_inst11.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36645\,
            ce => \N__36359\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.pwm_out_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011100000"
        )
    port map (
            in0 => \N__27483\,
            in1 => \N__32988\,
            in2 => \N__29883\,
            in3 => \N__27493\,
            lcout => \b2v_inst11.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36651\,
            ce => 'H',
            sr => \N__27472\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__29874\,
            in1 => \N__29837\,
            in2 => \_gnd_net_\,
            in3 => \N__32987\,
            lcout => OPEN,
            ltout => \b2v_inst11.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIJK34_0_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29806\,
            in2 => \N__27463\,
            in3 => \N__35915\,
            lcout => \b2v_inst11.curr_stateZ0Z_0\,
            ltout => \b2v_inst11.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_RNIOCA3_0_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__35916\,
            in1 => \_gnd_net_\,
            in2 => \N__27460\,
            in3 => \N__29836\,
            lcout => \b2v_inst11.count_0_sqmuxa_i\,
            ltout => \b2v_inst11.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.count_RNI_0_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__32438\,
            in1 => \_gnd_net_\,
            in2 => \N__27373\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27363\,
            in2 => \N__27352\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30398\,
            in2 => \_gnd_net_\,
            in3 => \N__27841\,
            lcout => \b2v_inst36.un2_count_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_1\,
            carryout => \b2v_inst36.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30365\,
            in2 => \_gnd_net_\,
            in3 => \N__27838\,
            lcout => \b2v_inst36.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_2\,
            carryout => \b2v_inst36.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30978\,
            in1 => \N__27835\,
            in2 => \_gnd_net_\,
            in3 => \N__27808\,
            lcout => \b2v_inst36.count_rst_10\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_3\,
            carryout => \b2v_inst36.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30321\,
            in2 => \_gnd_net_\,
            in3 => \N__27805\,
            lcout => \b2v_inst36.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_4\,
            carryout => \b2v_inst36.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30979\,
            in1 => \N__27801\,
            in2 => \_gnd_net_\,
            in3 => \N__27775\,
            lcout => \b2v_inst36.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_5\,
            carryout => \b2v_inst36.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31015\,
            in2 => \_gnd_net_\,
            in3 => \N__27772\,
            lcout => \b2v_inst36.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_6\,
            carryout => \b2v_inst36.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27902\,
            in2 => \_gnd_net_\,
            in3 => \N__27769\,
            lcout => \b2v_inst36.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_7\,
            carryout => \b2v_inst36.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30973\,
            in1 => \N__27766\,
            in2 => \_gnd_net_\,
            in3 => \N__27730\,
            lcout => \b2v_inst36.count_rst_5\,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \b2v_inst36.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28142\,
            in2 => \_gnd_net_\,
            in3 => \N__27727\,
            lcout => \b2v_inst36.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_9\,
            carryout => \b2v_inst36.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28025\,
            in2 => \_gnd_net_\,
            in3 => \N__28000\,
            lcout => \b2v_inst36.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_10\,
            carryout => \b2v_inst36.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30950\,
            in1 => \N__27997\,
            in2 => \_gnd_net_\,
            in3 => \N__27958\,
            lcout => \b2v_inst36.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_11\,
            carryout => \b2v_inst36.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30974\,
            in1 => \N__28107\,
            in2 => \_gnd_net_\,
            in3 => \N__27955\,
            lcout => \b2v_inst36.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_12\,
            carryout => \b2v_inst36.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_13_c_RNILPEV_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__30951\,
            in1 => \N__27948\,
            in2 => \_gnd_net_\,
            in3 => \N__27916\,
            lcout => \b2v_inst36.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst36.un2_count_1_cry_13\,
            carryout => \b2v_inst36.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__28059\,
            in1 => \N__30952\,
            in2 => \_gnd_net_\,
            in3 => \N__27913\,
            lcout => \b2v_inst36.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_15_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28071\,
            lcout => \b2v_inst36.count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36659\,
            ce => \N__30733\,
            sr => \N__30588\
        );

    \b2v_inst36.count_RNIRKI01_8_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27910\,
            in1 => \N__27856\,
            in2 => \_gnd_net_\,
            in3 => \N__30707\,
            lcout => \b2v_inst36.countZ0Z_8\,
            ltout => \b2v_inst36.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_8_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__30859\,
            in1 => \N__27877\,
            in2 => \N__27859\,
            in3 => \N__30977\,
            lcout => \b2v_inst36.count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36653\,
            ce => \N__30710\,
            sr => \N__30580\
        );

    \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__30975\,
            in1 => \N__28125\,
            in2 => \N__28149\,
            in3 => \N__30858\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI6MB61_10_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30708\,
            in1 => \_gnd_net_\,
            in2 => \N__28153\,
            in3 => \N__28114\,
            lcout => \b2v_inst36.countZ0Z_10\,
            ltout => \b2v_inst36.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_10_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__30976\,
            in1 => \N__28126\,
            in2 => \N__28117\,
            in3 => \N__30860\,
            lcout => \b2v_inst36.count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36653\,
            ce => \N__30710\,
            sr => \N__30580\
        );

    \b2v_inst36.count_RNIJMDV_13_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__30709\,
            in1 => \N__28087\,
            in2 => \_gnd_net_\,
            in3 => \N__28095\,
            lcout => \b2v_inst36.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_13_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst36.count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36653\,
            ce => \N__30710\,
            sr => \N__30580\
        );

    \b2v_inst36.count_RNINSFV_15_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28081\,
            in1 => \N__30711\,
            in2 => \_gnd_net_\,
            in3 => \N__28072\,
            lcout => \b2v_inst36.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIL1AS2_0_2_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__31940\,
            in1 => \N__28036\,
            in2 => \N__31219\,
            in3 => \N__31191\,
            lcout => \b2v_inst5.un12_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIL1AS2_2_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__28035\,
            in1 => \N__31873\,
            in2 => \_gnd_net_\,
            in3 => \N__31214\,
            lcout => \b2v_inst5.un2_count_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_2_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31215\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36647\,
            ce => \N__31939\,
            sr => \N__32092\
        );

    \b2v_inst5.count_RNIN4BS2_3_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__28177\,
            in1 => \N__32090\,
            in2 => \N__31177\,
            in3 => \N__31874\,
            lcout => \b2v_inst5.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI_1_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31548\,
            in2 => \_gnd_net_\,
            in3 => \N__31250\,
            lcout => \b2v_inst5.count_RNIZ0Z_1\,
            ltout => \b2v_inst5.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIUHFI2_1_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__28165\,
            in1 => \N__31872\,
            in2 => \N__28180\,
            in3 => \N__32089\,
            lcout => \b2v_inst5.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_3_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__32091\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31176\,
            lcout => \b2v_inst5.count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36647\,
            ce => \N__31939\,
            sr => \N__32092\
        );

    \b2v_inst5.count_1_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28171\,
            in2 => \_gnd_net_\,
            in3 => \N__32093\,
            lcout => \b2v_inst5.count_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36647\,
            ce => \N__31939\,
            sr => \N__32092\
        );

    \b2v_inst5.count_RNIJJOV_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__31555\,
            in1 => \N__31517\,
            in2 => \_gnd_net_\,
            in3 => \N__32085\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_rst_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNITGFI2_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31459\,
            in2 => \N__28159\,
            in3 => \N__31870\,
            lcout => \b2v_inst5.un2_count_1_cry_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_12_c_RNIRRH21_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31386\,
            in1 => \N__31519\,
            in2 => \N__31372\,
            in3 => \N__32087\,
            lcout => \b2v_inst5.count_rst_1\,
            ltout => \b2v_inst5.count_rst_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIPDG23_13_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28305\,
            in2 => \N__28156\,
            in3 => \N__31871\,
            lcout => \b2v_inst5.un2_count_1_axb_13\,
            ltout => \b2v_inst5.un2_count_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_13_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__31525\,
            in1 => \N__32088\,
            in2 => \N__28318\,
            in3 => \N__31371\,
            lcout => \b2v_inst5.count_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36640\,
            ce => \N__31909\,
            sr => \N__32172\
        );

    \b2v_inst5.count_RNIPDG23_0_13_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__31251\,
            in1 => \N__28315\,
            in2 => \N__28309\,
            in3 => \N__31910\,
            lcout => \b2v_inst5.un12_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_c_RNIFEP91_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31059\,
            in1 => \N__31518\,
            in2 => \N__31102\,
            in3 => \N__32086\,
            lcout => \b2v_inst5.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI_15_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31425\,
            in1 => \N__31299\,
            in2 => \N__31345\,
            in3 => \N__31556\,
            lcout => \b2v_inst5.un12_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28707\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28261\,
            in2 => \N__28386\,
            in3 => \N__28240\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28237\,
            in2 => \N__28387\,
            in3 => \N__28222\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32468\,
            in2 => \N__28219\,
            in3 => \N__28201\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28198\,
            in2 => \N__32475\,
            in3 => \N__28183\,
            lcout => \b2v_inst11.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__32497\,
            in1 => \N__28385\,
            in2 => \N__28417\,
            in3 => \N__28399\,
            lcout => \b2v_inst11.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un145_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__28396\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28390\,
            lcout => \b2v_inst11.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32467\,
            lcout => \b2v_inst11.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28543\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28366\,
            in2 => \N__28803\,
            in3 => \N__28351\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28799\,
            in2 => \N__28489\,
            in3 => \N__28342\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28477\,
            in2 => \N__28831\,
            in3 => \N__28330\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28829\,
            in2 => \N__28468\,
            in3 => \N__28321\,
            lcout => \b2v_inst11.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__31681\,
            in1 => \N__28456\,
            in2 => \N__28804\,
            in3 => \N__28516\,
            lcout => \b2v_inst11.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un110_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28429\,
            in3 => \N__28513\,
            lcout => \b2v_inst11.mult1_un110_sum_s_8\,
            ltout => \b2v_inst11.mult1_un110_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28510\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29250\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35077\,
            in2 => \N__28446\,
            in3 => \N__28480\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28442\,
            in2 => \N__34837\,
            in3 => \N__28471\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34810\,
            in2 => \N__35218\,
            in3 => \N__28459\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35217\,
            in2 => \N__34786\,
            in3 => \N__28450\,
            lcout => \b2v_inst11.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__28825\,
            in1 => \N__35269\,
            in2 => \N__28447\,
            in3 => \N__28420\,
            lcout => \b2v_inst11.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un103_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35248\,
            in3 => \N__28834\,
            lcout => \b2v_inst11.mult1_un103_sum_s_8\,
            ltout => \b2v_inst11.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__28807\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_6_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28786\,
            in2 => \N__33634\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_dutycycle_53_axb_0\,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28693\,
            in2 => \N__33633\,
            in3 => \N__28660\,
            lcout => \b2v_inst11.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_0\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30283\,
            in2 => \N__29272\,
            in3 => \N__28639\,
            lcout => \b2v_inst11.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_1\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28636\,
            in2 => \N__30296\,
            in3 => \N__28609\,
            lcout => \b2v_inst11.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_2\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28605\,
            in2 => \N__28588\,
            in3 => \N__28561\,
            lcout => \b2v_inst11.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_3\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29393\,
            in2 => \N__28558\,
            in3 => \N__28528\,
            lcout => \b2v_inst11.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_4\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29260\,
            in2 => \N__29401\,
            in3 => \N__29239\,
            lcout => \b2v_inst11.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_5\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29236\,
            in2 => \N__29224\,
            in3 => \N__29134\,
            lcout => \b2v_inst11.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_6\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29131\,
            in2 => \N__29074\,
            in3 => \N__29059\,
            lcout => \b2v_inst11.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29056\,
            in2 => \N__29029\,
            in3 => \N__28945\,
            lcout => \b2v_inst11.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_8\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28897\,
            in2 => \N__28942\,
            in3 => \N__28927\,
            lcout => \b2v_inst11.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_9\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29736\,
            in2 => \N__28924\,
            in3 => \N__28915\,
            lcout => \b2v_inst11.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_10\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29589\,
            in2 => \N__28912\,
            in3 => \N__28903\,
            lcout => \b2v_inst11.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_11\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28898\,
            in2 => \N__28846\,
            in3 => \N__28837\,
            lcout => \b2v_inst11.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_12\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29732\,
            in2 => \N__29659\,
            in3 => \N__29650\,
            lcout => \b2v_inst11.mult1_un47_sum\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_13\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29590\,
            in2 => \N__29647\,
            in3 => \N__29629\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0\,
            ltout => OPEN,
            carryin => \b2v_inst11.un1_dutycycle_53_cry_14\,
            carryout => \b2v_inst11.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29626\,
            in2 => \N__29607\,
            in3 => \N__29545\,
            lcout => \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0\,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => \b2v_inst11.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.CO2_THRU_LUT4_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29542\,
            lcout => \b2v_inst11.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29923\,
            in3 => \N__29774\,
            lcout => \b2v_inst11.mult1_un47_sum_s_4_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30024\,
            lcout => \b2v_inst11.mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.dutycycle_RNI_1_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__29524\,
            in1 => \N__29391\,
            in2 => \N__30297\,
            in3 => \N__33362\,
            lcout => \b2v_inst11.dutycycle_RNI_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29920\,
            in2 => \N__29779\,
            in3 => \N__29793\,
            lcout => \b2v_inst11.mult1_un40_sum_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.curr_state_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32983\,
            in2 => \N__29887\,
            in3 => \N__29839\,
            lcout => \b2v_inst11.curr_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36633\,
            ce => \N__36365\,
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29922\,
            in2 => \N__29794\,
            in3 => \N__29778\,
            lcout => \b2v_inst11.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30054\,
            in3 => \N__29938\,
            lcout => \b2v_inst11.mult1_un47_sum_s_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__30086\,
            in1 => \N__30087\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33261\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29761\,
            in3 => \N__29749\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30034\,
            in2 => \N__30010\,
            in3 => \N__29746\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30437\,
            in2 => \N__29977\,
            in3 => \N__29743\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30438\,
            in2 => \N__29953\,
            in3 => \N__29740\,
            lcout => \b2v_inst11.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36187\,
            in1 => \N__30088\,
            in2 => \N__30070\,
            in3 => \N__30061\,
            lcout => \b2v_inst11.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un54_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29937\,
            in2 => \N__30058\,
            in3 => \N__30037\,
            lcout => \b2v_inst11.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__30005\,
            in1 => \N__30006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30028\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29896\,
            in3 => \N__29992\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29989\,
            in3 => \N__29968\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30436\,
            in2 => \N__29965\,
            in3 => \N__29944\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un47_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29941\,
            lcout => \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29921\,
            lcout => \b2v_inst11.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30291\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33363\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30190\,
            in2 => \N__30488\,
            in3 => \N__30184\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30181\,
            in2 => \N__30490\,
            in3 => \N__30169\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30166\,
            in2 => \N__31747\,
            in3 => \N__30148\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30145\,
            in2 => \N__31746\,
            in3 => \N__30127\,
            lcout => \b2v_inst11.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__33954\,
            in1 => \N__30124\,
            in2 => \N__30489\,
            in3 => \N__30106\,
            lcout => \b2v_inst11.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un159_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30103\,
            in2 => \_gnd_net_\,
            in3 => \N__30091\,
            lcout => \b2v_inst11.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31739\,
            lcout => \b2v_inst11.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.curr_state_1_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30466\,
            lcout => \b2v_inst5.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36658\,
            ce => \N__36360\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNI_2_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30366\,
            in1 => \N__31013\,
            in2 => \N__30325\,
            in3 => \N__30406\,
            lcout => \b2v_inst36.un12_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__30348\,
            in1 => \N__30981\,
            in2 => \N__30861\,
            in3 => \N__30367\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNIH5D01_3_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30334\,
            in2 => \N__30370\,
            in3 => \N__30725\,
            lcout => \b2v_inst36.countZ0Z_3\,
            ltout => \b2v_inst36.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_3_LC_11_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__30349\,
            in1 => \N__30985\,
            in2 => \N__30337\,
            in3 => \N__30854\,
            lcout => \b2v_inst36.count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36664\,
            ce => \N__30731\,
            sr => \N__30589\
        );

    \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__30852\,
            in1 => \N__31038\,
            in2 => \N__30988\,
            in3 => \N__30320\,
            lcout => OPEN,
            ltout => \b2v_inst36.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_RNILBF01_5_LC_11_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__30726\,
            in1 => \_gnd_net_\,
            in2 => \N__30328\,
            in3 => \N__31021\,
            lcout => \b2v_inst36.countZ0Z_5\,
            ltout => \b2v_inst36.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst36.count_5_LC_11_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000000000"
        )
    port map (
            in0 => \N__30853\,
            in1 => \N__31039\,
            in2 => \N__31024\,
            in3 => \N__30987\,
            lcout => \b2v_inst36.count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36664\,
            ce => \N__30731\,
            sr => \N__30589\
        );

    \b2v_inst36.count_7_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__31014\,
            in1 => \N__30986\,
            in2 => \N__30862\,
            in3 => \N__30766\,
            lcout => \b2v_inst36.count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36664\,
            ce => \N__30731\,
            sr => \N__30589\
        );

    \b2v_inst6.count_14_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__33991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36662\,
            ce => \N__35058\,
            sr => \N__36129\
        );

    \b2v_inst6.count_RNIPG489_14_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30505\,
            in1 => \N__33990\,
            in2 => \_gnd_net_\,
            in3 => \N__35040\,
            lcout => \b2v_inst6.countZ0Z_14\,
            ltout => \b2v_inst6.countZ0Z_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_2_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__34147\,
            in1 => \N__34044\,
            in2 => \N__30499\,
            in3 => \N__33871\,
            lcout => \b2v_inst6.count_1_i_a3_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_13_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34159\,
            lcout => \b2v_inst6.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36662\,
            ce => \N__35058\,
            sr => \N__36129\
        );

    \b2v_inst6.count_RNIRB4V8_6_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34029\,
            in1 => \N__30496\,
            in2 => \_gnd_net_\,
            in3 => \N__35039\,
            lcout => \b2v_inst6.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_6_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34030\,
            lcout => \b2v_inst6.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36662\,
            ce => \N__35058\,
            sr => \N__36129\
        );

    \b2v_inst6.count_RNIJVVU8_2_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34351\,
            in1 => \N__34362\,
            in2 => \_gnd_net_\,
            in3 => \N__35038\,
            lcout => \b2v_inst6.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_1_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31255\,
            in2 => \N__31564\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_1_c_RNI92J91_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32175\,
            in1 => \N__31231\,
            in2 => \_gnd_net_\,
            in3 => \N__31198\,
            lcout => \b2v_inst5.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_1\,
            carryout => \b2v_inst5.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31195\,
            in2 => \_gnd_net_\,
            in3 => \N__31159\,
            lcout => \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_2\,
            carryout => \b2v_inst5.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31156\,
            in2 => \_gnd_net_\,
            in3 => \N__31114\,
            lcout => \b2v_inst5.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_3\,
            carryout => \b2v_inst5.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_4_c_RNIC8M91_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32177\,
            in1 => \N__32269\,
            in2 => \_gnd_net_\,
            in3 => \N__31111\,
            lcout => \b2v_inst5.count_rst_9\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_4\,
            carryout => \b2v_inst5.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_5_c_RNIDAN91_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32176\,
            in1 => \N__32242\,
            in2 => \_gnd_net_\,
            in3 => \N__31108\,
            lcout => \b2v_inst5.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_5\,
            carryout => \b2v_inst5.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_6_c_RNIECO91_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32178\,
            in1 => \N__32191\,
            in2 => \_gnd_net_\,
            in3 => \N__31105\,
            lcout => \b2v_inst5.count_rst_7\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_6\,
            carryout => \b2v_inst5.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31101\,
            in2 => \_gnd_net_\,
            in3 => \N__31042\,
            lcout => \b2v_inst5.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_7\,
            carryout => \b2v_inst5.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31659\,
            in2 => \_gnd_net_\,
            in3 => \N__31450\,
            lcout => \b2v_inst5.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \b2v_inst5.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31599\,
            in2 => \_gnd_net_\,
            in3 => \N__31447\,
            lcout => \b2v_inst5.un2_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_9\,
            carryout => \b2v_inst5.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_10_c_RNIPNF21_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32179\,
            in1 => \N__31956\,
            in2 => \_gnd_net_\,
            in3 => \N__31429\,
            lcout => \b2v_inst5.count_rst_3\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_10\,
            carryout => \b2v_inst5.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_11_c_RNIQPG21_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32180\,
            in1 => \N__31426\,
            in2 => \_gnd_net_\,
            in3 => \N__31393\,
            lcout => \b2v_inst5.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_11\,
            carryout => \b2v_inst5.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31390\,
            in2 => \_gnd_net_\,
            in3 => \N__31348\,
            lcout => \b2v_inst5.un2_count_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_12\,
            carryout => \b2v_inst5.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_13_c_RNISTI21_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__32181\,
            in1 => \N__31341\,
            in2 => \_gnd_net_\,
            in3 => \N__31306\,
            lcout => \b2v_inst5.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst5.un2_count_1_cry_13\,
            carryout => \b2v_inst5.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_14_c_RNITVJ21_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31303\,
            in1 => \N__32182\,
            in2 => \_gnd_net_\,
            in3 => \N__31288\,
            lcout => \b2v_inst5.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_15_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31278\,
            lcout => \b2v_inst5.count_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36655\,
            ce => \N__31927\,
            sr => \N__32174\
        );

    \b2v_inst5.un2_count_1_cry_8_c_RNIGGQ91_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31660\,
            in1 => \N__31520\,
            in2 => \N__31648\,
            in3 => \N__32140\,
            lcout => \b2v_inst5.count_rst_5\,
            ltout => \b2v_inst5.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNI3NHS2_9_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__31633\,
            in1 => \_gnd_net_\,
            in2 => \N__31663\,
            in3 => \N__31882\,
            lcout => \b2v_inst5.un2_count_1_axb_9\,
            ltout => \b2v_inst5.un2_count_1_axb_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_9_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31647\,
            in1 => \N__31522\,
            in2 => \N__31636\,
            in3 => \N__32143\,
            lcout => \b2v_inst5.count_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36648\,
            ce => \N__31883\,
            sr => \N__32170\
        );

    \b2v_inst5.count_RNI3NHS2_0_9_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__31632\,
            in1 => \N__31881\,
            in2 => \N__31624\,
            in3 => \N__31595\,
            lcout => \b2v_inst5.un12_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un2_count_1_cry_9_c_RNIHIR91_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31582\,
            in1 => \N__31523\,
            in2 => \N__31600\,
            in3 => \N__32139\,
            lcout => OPEN,
            ltout => \b2v_inst5.count_rst_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIC1Q93_10_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31570\,
            in2 => \N__31603\,
            in3 => \N__31880\,
            lcout => \b2v_inst5.countZ0Z_10\,
            ltout => \b2v_inst5.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_10_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__31581\,
            in1 => \N__31521\,
            in2 => \N__31573\,
            in3 => \N__32142\,
            lcout => \b2v_inst5.count_1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36648\,
            ce => \N__31883\,
            sr => \N__32170\
        );

    \b2v_inst5.count_0_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32141\,
            in1 => \N__31560\,
            in2 => \_gnd_net_\,
            in3 => \N__31524\,
            lcout => \b2v_inst5.count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36648\,
            ce => \N__31883\,
            sr => \N__32170\
        );

    \b2v_inst5.count_6_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36641\,
            ce => \N__31907\,
            sr => \N__32171\
        );

    \b2v_inst5.count_RNIRADS2_5_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32211\,
            in1 => \N__31884\,
            in2 => \_gnd_net_\,
            in3 => \N__32231\,
            lcout => \b2v_inst5.un2_count_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_5_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36641\,
            ce => \N__31907\,
            sr => \N__32171\
        );

    \b2v_inst5.count_RNITDES2_6_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__32260\,
            in1 => \N__31885\,
            in2 => \_gnd_net_\,
            in3 => \N__32253\,
            lcout => \b2v_inst5.countZ0Z_6\,
            ltout => \b2v_inst5.countZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIRADS2_0_5_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000111"
        )
    port map (
            in0 => \N__31887\,
            in1 => \N__32233\,
            in2 => \N__32215\,
            in3 => \N__32212\,
            lcout => \b2v_inst5.un12_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_RNIVGFS2_7_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__31986\,
            in1 => \N__31886\,
            in2 => \_gnd_net_\,
            in3 => \N__31976\,
            lcout => \b2v_inst5.un2_count_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.count_7_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst5.count_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36641\,
            ce => \N__31907\,
            sr => \N__32171\
        );

    \b2v_inst5.count_RNIVGFS2_0_7_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__31987\,
            in1 => \N__31978\,
            in2 => \N__31963\,
            in3 => \N__31908\,
            lcout => \b2v_inst5.un12_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31730\,
            lcout => \b2v_inst11.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31690\,
            lcout => \b2v_inst11.mult1_un110_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32587\,
            lcout => \b2v_inst11.mult1_un117_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32560\,
            lcout => \b2v_inst11.mult1_un124_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32521\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un145_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32479\,
            lcout => \b2v_inst11.mult1_un138_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32446\,
            in1 => \N__32410\,
            in2 => \N__33889\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32374\,
            in2 => \N__33190\,
            in3 => \N__32404\,
            lcout => \b2v_inst11.N_5530_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_0\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32368\,
            in1 => \N__32323\,
            in2 => \N__32332\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5531_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_1\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32317\,
            in1 => \N__32275\,
            in2 => \N__32287\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5532_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_2\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32950\,
            in1 => \N__32914\,
            in2 => \N__32923\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5533_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_3\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32908\,
            in1 => \N__32866\,
            in2 => \N__32881\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5534_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_4\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32824\,
            in2 => \N__32860\,
            in3 => \N__32851\,
            lcout => \b2v_inst11.N_5535_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_5\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32818\,
            in1 => \N__32776\,
            in2 => \N__32785\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5536_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_6\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32770\,
            in1 => \N__32743\,
            in2 => \N__32734\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5537_i\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32725\,
            in1 => \N__32680\,
            in2 => \N__32695\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5538_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_8\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32674\,
            in1 => \N__34546\,
            in2 => \N__32638\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5539_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_9\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33196\,
            in2 => \N__32596\,
            in3 => \N__32629\,
            lcout => \b2v_inst11.N_5540_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_10\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33175\,
            in2 => \N__33103\,
            in3 => \N__33127\,
            lcout => \b2v_inst11.N_5541_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_11\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33094\,
            in1 => \N__34552\,
            in2 => \N__33070\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5542_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_12\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33061\,
            in1 => \N__35065\,
            in2 => \N__33034\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5543_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_13\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__33025\,
            in1 => \N__33238\,
            in2 => \N__33001\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.N_5544_i\,
            ltout => OPEN,
            carryin => \b2v_inst11.un85_clk_100khz_cry_14\,
            carryout => \b2v_inst11.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32992\,
            lcout => \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33168\,
            lcout => \b2v_inst11.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35337\,
            lcout => \b2v_inst11.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35136\,
            lcout => \b2v_inst11.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35181\,
            lcout => \b2v_inst11.mult1_un89_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33970\,
            lcout => \b2v_inst11.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35382\,
            lcout => \b2v_inst11.mult1_un82_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33169\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33148\,
            in2 => \N__35355\,
            in3 => \N__33142\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35351\,
            in2 => \N__35110\,
            in3 => \N__33139\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35098\,
            in2 => \N__35383\,
            in3 => \N__33136\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35381\,
            in2 => \N__35089\,
            in3 => \N__33133\,
            lcout => \b2v_inst11.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35180\,
            in1 => \N__35410\,
            in2 => \N__35356\,
            in3 => \N__33130\,
            lcout => \b2v_inst11.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un89_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35398\,
            in3 => \N__33367\,
            lcout => \b2v_inst11.mult1_un89_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36230\,
            lcout => \b2v_inst11.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33364\,
            lcout => \b2v_inst11.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33262\,
            lcout => \b2v_inst11.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33229\,
            lcout => \b2v_inst11.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35527\,
            lcout => \b2v_inst11.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35448\,
            lcout => \b2v_inst11.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33228\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33205\,
            in2 => \N__36165\,
            in3 => \N__33199\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36161\,
            in2 => \N__33499\,
            in3 => \N__33484\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33481\,
            in2 => \N__36196\,
            in3 => \N__33472\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36194\,
            in2 => \N__33469\,
            in3 => \N__33457\,
            lcout => \b2v_inst11.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35443\,
            in1 => \N__33454\,
            in2 => \N__36166\,
            in3 => \N__33445\,
            lcout => \b2v_inst11.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un61_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33442\,
            in3 => \N__33430\,
            lcout => \b2v_inst11.mult1_un61_sum_s_8\,
            ltout => \b2v_inst11.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33427\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__35654\,
            in1 => \N__36148\,
            in2 => \_gnd_net_\,
            in3 => \N__36819\,
            lcout => \b2v_inst6.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst31.un6_output_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__34711\,
            in1 => \N__33424\,
            in2 => \N__33802\,
            in3 => \N__33412\,
            lcout => \VCCIN_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIUL1J2_0_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__35652\,
            in1 => \N__36147\,
            in2 => \_gnd_net_\,
            in3 => \N__36817\,
            lcout => \b2v_inst6.N_276_0\,
            ltout => \b2v_inst6.N_276_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__36402\,
            in1 => \N__33820\,
            in2 => \N__33847\,
            in3 => \N__35632\,
            lcout => \b2v_inst6.delayed_vccin_vccinaux_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__33844\,
            in1 => \N__33832\,
            in2 => \_gnd_net_\,
            in3 => \N__33796\,
            lcout => \b2v_inst6.N_192\,
            ltout => \b2v_inst6.N_192_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIUL1J2_0_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__36818\,
            in1 => \_gnd_net_\,
            in2 => \N__33823\,
            in3 => \N__35653\,
            lcout => \b2v_inst6.curr_state_RNIUL1J2Z0Z_0\,
            ltout => \b2v_inst6.curr_state_RNIUL1J2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU0GV5_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__33819\,
            in1 => \N__36401\,
            in2 => \N__33811\,
            in3 => \N__33808\,
            lcout => OPEN,
            ltout => \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__33797\,
            in1 => \_gnd_net_\,
            in2 => \N__33691\,
            in3 => \_gnd_net_\,
            lcout => \N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33628\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33529\,
            in2 => \N__33918\,
            in3 => \N__33955\,
            lcout => \G_2836\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_0\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33914\,
            in2 => \N__33520\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_1\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33508\,
            in2 => \N__33966\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33979\,
            in2 => \N__33965\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33928\,
            in2 => \N__33919\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un166_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__33901\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33892\,
            lcout => \b2v_inst11.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34900\,
            in2 => \N__34459\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_1_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_1_c_RNID55Q2_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36112\,
            in1 => \N__33870\,
            in2 => \_gnd_net_\,
            in3 => \N__33859\,
            lcout => \b2v_inst6.count_rst_12\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_1\,
            carryout => \b2v_inst6.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34535\,
            in2 => \_gnd_net_\,
            in3 => \N__33856\,
            lcout => \b2v_inst6.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_2\,
            carryout => \b2v_inst6.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34227\,
            in2 => \_gnd_net_\,
            in3 => \N__33853\,
            lcout => \b2v_inst6.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_3\,
            carryout => \b2v_inst6.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34096\,
            in2 => \_gnd_net_\,
            in3 => \N__33850\,
            lcout => \b2v_inst6.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_4\,
            carryout => \b2v_inst6.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_5_c_RNIHD9Q2_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__36113\,
            in1 => \_gnd_net_\,
            in2 => \N__34045\,
            in3 => \N__34021\,
            lcout => \b2v_inst6.count_rst_8\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_5\,
            carryout => \b2v_inst6.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34409\,
            in2 => \_gnd_net_\,
            in3 => \N__34018\,
            lcout => \b2v_inst6.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_6\,
            carryout => \b2v_inst6.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34333\,
            in2 => \_gnd_net_\,
            in3 => \N__34015\,
            lcout => \b2v_inst6.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_7\,
            carryout => \b2v_inst6.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34073\,
            in2 => \_gnd_net_\,
            in3 => \N__34012\,
            lcout => \b2v_inst6.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_12_2_0_\,
            carryout => \b2v_inst6.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_9_c_RNILLDQ2_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36085\,
            in1 => \N__34279\,
            in2 => \_gnd_net_\,
            in3 => \N__34009\,
            lcout => \b2v_inst6.count_rst_4\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_9\,
            carryout => \b2v_inst6.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34626\,
            in2 => \_gnd_net_\,
            in3 => \N__34006\,
            lcout => \b2v_inst6.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_10\,
            carryout => \b2v_inst6.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_11_c_RNIUTM13_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__36086\,
            in1 => \_gnd_net_\,
            in2 => \N__34249\,
            in3 => \N__34003\,
            lcout => \b2v_inst6.count_rst_2\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_11\,
            carryout => \b2v_inst6.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_12_c_RNIVVN13_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36088\,
            in1 => \N__34143\,
            in2 => \_gnd_net_\,
            in3 => \N__34000\,
            lcout => \b2v_inst6.count_rst_1\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_12\,
            carryout => \b2v_inst6.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_13_c_RNI02P13_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36087\,
            in1 => \N__33997\,
            in2 => \_gnd_net_\,
            in3 => \N__33982\,
            lcout => \b2v_inst6.count_rst_0\,
            ltout => OPEN,
            carryin => \b2v_inst6.un2_count_1_cry_13\,
            carryout => \b2v_inst6.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_14_c_RNI14Q13_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__36089\,
            in1 => \N__34651\,
            in2 => \_gnd_net_\,
            in3 => \N__34171\,
            lcout => \b2v_inst6.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIND389_13_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34168\,
            in1 => \N__34158\,
            in2 => \_gnd_net_\,
            in3 => \N__35043\,
            lcout => \b2v_inst6.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_5_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__34095\,
            in1 => \N__36124\,
            in2 => \N__36788\,
            in3 => \N__34126\,
            lcout => \b2v_inst6.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36663\,
            ce => \N__35059\,
            sr => \N__36114\
        );

    \b2v_inst6.un2_count_1_cry_8_c_RNIKJCQ2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34059\,
            in1 => \N__36773\,
            in2 => \N__34078\,
            in3 => \N__36083\,
            lcout => \b2v_inst6.count_rst_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIP83V8_5_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34132\,
            in1 => \N__35041\,
            in2 => \_gnd_net_\,
            in3 => \N__34111\,
            lcout => \b2v_inst6.countZ0Z_5\,
            ltout => \b2v_inst6.countZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_4_c_RNIGB8Q2_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34125\,
            in1 => \N__36772\,
            in2 => \N__34114\,
            in3 => \N__36082\,
            lcout => \b2v_inst6.count_rst_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI1L7V8_9_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34051\,
            in1 => \N__35042\,
            in2 => \_gnd_net_\,
            in3 => \N__34105\,
            lcout => \b2v_inst6.countZ0Z_9\,
            ltout => \b2v_inst6.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_5_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34410\,
            in1 => \N__34331\,
            in2 => \N__34099\,
            in3 => \N__34094\,
            lcout => \b2v_inst6.count_1_i_a3_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_9_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__36084\,
            in1 => \N__34074\,
            in2 => \N__36789\,
            in3 => \N__34060\,
            lcout => \b2v_inst6.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36663\,
            ce => \N__35059\,
            sr => \N__36114\
        );

    \b2v_inst6.count_7_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__34411\,
            in1 => \N__36774\,
            in2 => \N__36130\,
            in3 => \N__34438\,
            lcout => \b2v_inst6.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36663\,
            ce => \N__35059\,
            sr => \N__36114\
        );

    \b2v_inst6.count_12_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__34261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36661\,
            ce => \N__35053\,
            sr => \N__36118\
        );

    \b2v_inst6.count_RNIA0P09_10_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__34444\,
            in1 => \N__35020\,
            in2 => \_gnd_net_\,
            in3 => \N__34182\,
            lcout => \b2v_inst6.countZ0Z_10\,
            ltout => \b2v_inst6.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_3_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__34245\,
            in1 => \N__34223\,
            in2 => \N__34270\,
            in3 => \N__34536\,
            lcout => \b2v_inst6.count_1_i_a3_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNILA289_12_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34267\,
            in1 => \N__34260\,
            in2 => \_gnd_net_\,
            in3 => \N__35021\,
            lcout => \b2v_inst6.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_3_c_RNIF97Q2_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34203\,
            in1 => \N__36770\,
            in2 => \N__34228\,
            in3 => \N__36031\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIN52V8_4_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34189\,
            in2 => \N__34231\,
            in3 => \N__35019\,
            lcout => \b2v_inst6.countZ0Z_4\,
            ltout => \b2v_inst6.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_4_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34204\,
            in1 => \N__36771\,
            in2 => \N__34192\,
            in3 => \N__36032\,
            lcout => \b2v_inst6.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36661\,
            ce => \N__35053\,
            sr => \N__36118\
        );

    \b2v_inst6.count_10_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34183\,
            lcout => \b2v_inst6.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36661\,
            ce => \N__35053\,
            sr => \N__36118\
        );

    \b2v_inst6.un2_count_1_cry_6_c_RNIIFAQ2_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__34408\,
            in1 => \N__36781\,
            in2 => \N__36076\,
            in3 => \N__34437\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNITE5V8_7_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34423\,
            in2 => \N__34414\,
            in3 => \N__35022\,
            lcout => \b2v_inst6.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_7_c_RNIJHBQ2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34302\,
            in1 => \N__36782\,
            in2 => \N__34332\,
            in3 => \N__36037\,
            lcout => \b2v_inst6.count_rst_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_15_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34386\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36656\,
            ce => \N__35044\,
            sr => \N__36036\
        );

    \b2v_inst6.count_RNIRJ589_15_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34387\,
            in1 => \N__34375\,
            in2 => \_gnd_net_\,
            in3 => \N__35045\,
            lcout => \b2v_inst6.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_2_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34369\,
            lcout => \b2v_inst6.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36656\,
            ce => \N__35044\,
            sr => \N__36036\
        );

    \b2v_inst6.count_RNIVH6V8_8_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34285\,
            in1 => \N__34339\,
            in2 => \_gnd_net_\,
            in3 => \N__35017\,
            lcout => \b2v_inst6.countZ0Z_8\,
            ltout => \b2v_inst6.countZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_8_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__36030\,
            in1 => \N__36761\,
            in2 => \N__34306\,
            in3 => \N__34303\,
            lcout => \b2v_inst6.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36649\,
            ce => \N__35018\,
            sr => \N__36119\
        );

    \b2v_inst6.count_11_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__36029\,
            in1 => \N__36760\,
            in2 => \N__34492\,
            in3 => \N__34624\,
            lcout => \b2v_inst6.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36649\,
            ce => \N__35018\,
            sr => \N__36119\
        );

    \b2v_inst6.un2_count_1_cry_2_c_RNIE76Q2_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34512\,
            in1 => \N__36758\,
            in2 => \N__34537\,
            in3 => \N__36028\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIL21V8_3_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__35016\,
            in1 => \_gnd_net_\,
            in2 => \N__34540\,
            in3 => \N__34498\,
            lcout => \b2v_inst6.countZ0Z_3\,
            ltout => \b2v_inst6.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__34513\,
            in1 => \N__36759\,
            in2 => \N__34501\,
            in3 => \N__36120\,
            lcout => \b2v_inst6.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36649\,
            ce => \N__35018\,
            sr => \N__36119\
        );

    \b2v_inst6.count_RNIM2CM2_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__34564\,
            in1 => \_gnd_net_\,
            in2 => \N__34899\,
            in3 => \N__36039\,
            lcout => \b2v_inst6.count_RNIM2CM2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34563\,
            in2 => \_gnd_net_\,
            in3 => \N__34892\,
            lcout => \b2v_inst6.N_394\,
            ltout => \b2v_inst6.N_394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.un2_count_1_cry_10_c_RNITRL13_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__34488\,
            in1 => \N__34625\,
            in2 => \N__34471\,
            in3 => \N__36038\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_rst_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIJ7189_11_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34468\,
            in2 => \N__34462\,
            in3 => \N__35023\,
            lcout => \b2v_inst6.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRR6R8_0_1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__34675\,
            in1 => \N__34662\,
            in2 => \N__34995\,
            in3 => \N__36025\,
            lcout => \b2v_inst6.un2_count_1_axb_1\,
            ltout => \b2v_inst6.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNI_1_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34768\,
            in3 => \N__34882\,
            lcout => \b2v_inst6.count_RNI_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34765\,
            in1 => \N__34753\,
            in2 => \N__34738\,
            in3 => \N__34729\,
            lcout => \N_1661\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__36027\,
            in1 => \_gnd_net_\,
            in2 => \N__34666\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36634\,
            ce => \N__35046\,
            sr => \N__36128\
        );

    \b2v_inst6.count_RNIRR6R8_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__34674\,
            in1 => \N__34661\,
            in2 => \N__35057\,
            in3 => \N__36024\,
            lcout => OPEN,
            ltout => \b2v_inst6.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRR6R8_2_1_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__34644\,
            in1 => \_gnd_net_\,
            in2 => \N__34630\,
            in3 => \N__34627\,
            lcout => OPEN,
            ltout => \b2v_inst6.count_1_i_a3_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIRR6R8_3_1_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__34600\,
            in1 => \N__34588\,
            in2 => \N__34579\,
            in3 => \N__34576\,
            lcout => \b2v_inst6.N_389\,
            ltout => \b2v_inst6.N_389_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_0_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__36026\,
            in1 => \_gnd_net_\,
            in2 => \N__34555\,
            in3 => \N__34883\,
            lcout => \b2v_inst6.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36634\,
            ce => \N__35046\,
            sr => \N__36128\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35575\,
            lcout => \b2v_inst11.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35204\,
            lcout => \b2v_inst11.mult1_un96_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34863\,
            lcout => \b2v_inst11.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36232\,
            lcout => \b2v_inst11.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI87PU5_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__36699\,
            in1 => \N__36400\,
            in2 => \_gnd_net_\,
            in3 => \N__36023\,
            lcout => \b2v_inst6.count_en\,
            ltout => \b2v_inst6.count_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.count_RNIQQ6R8_0_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__34921\,
            in1 => \_gnd_net_\,
            in2 => \N__34909\,
            in3 => \N__34906\,
            lcout => \b2v_inst6.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34864\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34843\,
            in2 => \N__35154\,
            in3 => \N__34822\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35150\,
            in2 => \N__34819\,
            in3 => \N__34798\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35176\,
            in2 => \N__34795\,
            in3 => \N__34771\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35275\,
            in2 => \N__35182\,
            in3 => \N__35257\,
            lcout => \b2v_inst11.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35203\,
            in1 => \N__35254\,
            in2 => \N__35155\,
            in3 => \N__35233\,
            lcout => \b2v_inst11.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un96_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35230\,
            in3 => \N__35221\,
            lcout => \b2v_inst11.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35175\,
            lcout => \b2v_inst11.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35137\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35116\,
            in2 => \N__35544\,
            in3 => \N__35101\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35540\,
            in2 => \N__35314\,
            in3 => \N__35092\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35302\,
            in2 => \N__35574\,
            in3 => \N__35080\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35570\,
            in2 => \N__35293\,
            in3 => \N__35401\,
            lcout => \b2v_inst11.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35377\,
            in1 => \N__35281\,
            in2 => \N__35545\,
            in3 => \N__35389\,
            lcout => \b2v_inst11.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un82_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35590\,
            in3 => \N__35386\,
            lcout => \b2v_inst11.mult1_un82_sum_s_8\,
            ltout => \b2v_inst11.mult1_un82_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35359\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35338\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35320\,
            in2 => \N__35607\,
            in3 => \N__35305\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35603\,
            in2 => \N__35497\,
            in3 => \N__35296\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35476\,
            in2 => \N__36231\,
            in3 => \N__35284\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36226\,
            in2 => \N__35461\,
            in3 => \N__35611\,
            lcout => \b2v_inst11.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__35566\,
            in1 => \N__35416\,
            in2 => \N__35608\,
            in3 => \N__35581\,
            lcout => \b2v_inst11.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un75_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36256\,
            in3 => \N__35578\,
            lcout => \b2v_inst11.mult1_un75_sum_s_8\,
            ltout => \b2v_inst11.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__35548\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst11.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35526\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35503\,
            in2 => \N__36273\,
            in3 => \N__35488\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_2\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36269\,
            in2 => \N__35485\,
            in3 => \N__35470\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_3\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35467\,
            in2 => \N__35449\,
            in3 => \N__35452\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_4\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35447\,
            in2 => \N__35425\,
            in3 => \N__36286\,
            lcout => \b2v_inst11.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_5\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__36222\,
            in1 => \N__36283\,
            in2 => \N__36274\,
            in3 => \N__36247\,
            lcout => \b2v_inst11.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \b2v_inst11.mult1_un68_sum_cry_6\,
            carryout => \b2v_inst11.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__36244\,
            in3 => \N__36235\,
            lcout => \b2v_inst11.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36195\,
            lcout => \b2v_inst11.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI59E43_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__35944\,
            in1 => \N__35617\,
            in2 => \_gnd_net_\,
            in3 => \N__35898\,
            lcout => \b2v_inst6.curr_stateZ0Z_0\,
            ltout => \b2v_inst6.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNIM2CM2_0_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__35899\,
            in1 => \N__36146\,
            in2 => \N__36133\,
            in3 => \N__36820\,
            lcout => \b2v_inst6.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_0_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__36802\,
            in1 => \N__35631\,
            in2 => \N__36790\,
            in3 => \N__35655\,
            lcout => \b2v_inst6.curr_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36660\,
            ce => \N__36366\,
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI6AE43_1_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__35900\,
            in1 => \N__36670\,
            in2 => \N__36700\,
            in3 => \N__36706\,
            lcout => \b2v_inst6.curr_stateZ0Z_1\,
            ltout => \b2v_inst6.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m4_0_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__36787\,
            in1 => \N__35656\,
            in2 => \N__35635\,
            in3 => \N__35630\,
            lcout => \b2v_inst6.curr_state_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_RNI_1_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36800\,
            lcout => \b2v_inst6.N_2937_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36801\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36783\,
            lcout => \b2v_inst6.m6_i_a3\,
            ltout => \b2v_inst6.m6_i_a3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b2v_inst6.curr_state_1_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36692\,
            in2 => \N__36673\,
            in3 => \_gnd_net_\,
            lcout => \b2v_inst6.curr_state_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__36660\,
            ce => \N__36366\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
