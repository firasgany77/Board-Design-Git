// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 13 2022 16:56:57

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    input SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    input VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    input VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__37129;
    wire N__37128;
    wire N__37127;
    wire N__37118;
    wire N__37117;
    wire N__37116;
    wire N__37109;
    wire N__37108;
    wire N__37107;
    wire N__37100;
    wire N__37099;
    wire N__37098;
    wire N__37091;
    wire N__37090;
    wire N__37089;
    wire N__37082;
    wire N__37081;
    wire N__37080;
    wire N__37073;
    wire N__37072;
    wire N__37071;
    wire N__37064;
    wire N__37063;
    wire N__37062;
    wire N__37055;
    wire N__37054;
    wire N__37053;
    wire N__37046;
    wire N__37045;
    wire N__37044;
    wire N__37037;
    wire N__37036;
    wire N__37035;
    wire N__37028;
    wire N__37027;
    wire N__37026;
    wire N__37019;
    wire N__37018;
    wire N__37017;
    wire N__37010;
    wire N__37009;
    wire N__37008;
    wire N__37001;
    wire N__37000;
    wire N__36999;
    wire N__36992;
    wire N__36991;
    wire N__36990;
    wire N__36983;
    wire N__36982;
    wire N__36981;
    wire N__36974;
    wire N__36973;
    wire N__36972;
    wire N__36965;
    wire N__36964;
    wire N__36963;
    wire N__36956;
    wire N__36955;
    wire N__36954;
    wire N__36947;
    wire N__36946;
    wire N__36945;
    wire N__36938;
    wire N__36937;
    wire N__36936;
    wire N__36929;
    wire N__36928;
    wire N__36927;
    wire N__36920;
    wire N__36919;
    wire N__36918;
    wire N__36911;
    wire N__36910;
    wire N__36909;
    wire N__36902;
    wire N__36901;
    wire N__36900;
    wire N__36893;
    wire N__36892;
    wire N__36891;
    wire N__36884;
    wire N__36883;
    wire N__36882;
    wire N__36875;
    wire N__36874;
    wire N__36873;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36857;
    wire N__36856;
    wire N__36855;
    wire N__36848;
    wire N__36847;
    wire N__36846;
    wire N__36839;
    wire N__36838;
    wire N__36837;
    wire N__36820;
    wire N__36819;
    wire N__36818;
    wire N__36817;
    wire N__36814;
    wire N__36807;
    wire N__36802;
    wire N__36801;
    wire N__36800;
    wire N__36793;
    wire N__36790;
    wire N__36789;
    wire N__36788;
    wire N__36787;
    wire N__36784;
    wire N__36783;
    wire N__36782;
    wire N__36781;
    wire N__36778;
    wire N__36775;
    wire N__36774;
    wire N__36773;
    wire N__36772;
    wire N__36771;
    wire N__36770;
    wire N__36765;
    wire N__36762;
    wire N__36761;
    wire N__36760;
    wire N__36759;
    wire N__36758;
    wire N__36753;
    wire N__36742;
    wire N__36737;
    wire N__36732;
    wire N__36727;
    wire N__36722;
    wire N__36713;
    wire N__36706;
    wire N__36703;
    wire N__36700;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36678;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36663;
    wire N__36662;
    wire N__36661;
    wire N__36660;
    wire N__36659;
    wire N__36658;
    wire N__36657;
    wire N__36656;
    wire N__36655;
    wire N__36654;
    wire N__36653;
    wire N__36652;
    wire N__36651;
    wire N__36650;
    wire N__36649;
    wire N__36648;
    wire N__36647;
    wire N__36646;
    wire N__36645;
    wire N__36644;
    wire N__36643;
    wire N__36642;
    wire N__36641;
    wire N__36640;
    wire N__36639;
    wire N__36638;
    wire N__36637;
    wire N__36636;
    wire N__36635;
    wire N__36634;
    wire N__36633;
    wire N__36632;
    wire N__36631;
    wire N__36630;
    wire N__36629;
    wire N__36628;
    wire N__36627;
    wire N__36626;
    wire N__36625;
    wire N__36624;
    wire N__36623;
    wire N__36622;
    wire N__36621;
    wire N__36620;
    wire N__36619;
    wire N__36618;
    wire N__36617;
    wire N__36616;
    wire N__36615;
    wire N__36614;
    wire N__36613;
    wire N__36612;
    wire N__36611;
    wire N__36610;
    wire N__36609;
    wire N__36608;
    wire N__36607;
    wire N__36606;
    wire N__36605;
    wire N__36604;
    wire N__36603;
    wire N__36602;
    wire N__36601;
    wire N__36600;
    wire N__36599;
    wire N__36598;
    wire N__36597;
    wire N__36596;
    wire N__36595;
    wire N__36594;
    wire N__36593;
    wire N__36592;
    wire N__36591;
    wire N__36590;
    wire N__36589;
    wire N__36588;
    wire N__36587;
    wire N__36586;
    wire N__36585;
    wire N__36584;
    wire N__36583;
    wire N__36582;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36408;
    wire N__36407;
    wire N__36406;
    wire N__36405;
    wire N__36404;
    wire N__36403;
    wire N__36402;
    wire N__36401;
    wire N__36400;
    wire N__36397;
    wire N__36394;
    wire N__36391;
    wire N__36384;
    wire N__36381;
    wire N__36376;
    wire N__36373;
    wire N__36370;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36366;
    wire N__36365;
    wire N__36364;
    wire N__36363;
    wire N__36362;
    wire N__36361;
    wire N__36360;
    wire N__36359;
    wire N__36358;
    wire N__36357;
    wire N__36356;
    wire N__36355;
    wire N__36352;
    wire N__36349;
    wire N__36346;
    wire N__36343;
    wire N__36340;
    wire N__36337;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36273;
    wire N__36270;
    wire N__36269;
    wire N__36266;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36231;
    wire N__36230;
    wire N__36227;
    wire N__36226;
    wire N__36223;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36191;
    wire N__36188;
    wire N__36187;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36171;
    wire N__36166;
    wire N__36165;
    wire N__36162;
    wire N__36161;
    wire N__36158;
    wire N__36151;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36141;
    wire N__36138;
    wire N__36133;
    wire N__36130;
    wire N__36129;
    wire N__36128;
    wire N__36125;
    wire N__36124;
    wire N__36121;
    wire N__36120;
    wire N__36119;
    wire N__36118;
    wire N__36115;
    wire N__36114;
    wire N__36113;
    wire N__36112;
    wire N__36107;
    wire N__36104;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36089;
    wire N__36088;
    wire N__36087;
    wire N__36086;
    wire N__36085;
    wire N__36084;
    wire N__36083;
    wire N__36082;
    wire N__36077;
    wire N__36076;
    wire N__36067;
    wire N__36062;
    wire N__36057;
    wire N__36050;
    wire N__36043;
    wire N__36040;
    wire N__36039;
    wire N__36038;
    wire N__36037;
    wire N__36036;
    wire N__36033;
    wire N__36032;
    wire N__36031;
    wire N__36030;
    wire N__36029;
    wire N__36028;
    wire N__36027;
    wire N__36026;
    wire N__36025;
    wire N__36024;
    wire N__36023;
    wire N__36018;
    wire N__36009;
    wire N__36004;
    wire N__36001;
    wire N__35996;
    wire N__35991;
    wire N__35984;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35951;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35934;
    wire N__35933;
    wire N__35932;
    wire N__35931;
    wire N__35930;
    wire N__35929;
    wire N__35926;
    wire N__35925;
    wire N__35924;
    wire N__35923;
    wire N__35922;
    wire N__35919;
    wire N__35918;
    wire N__35917;
    wire N__35916;
    wire N__35915;
    wire N__35910;
    wire N__35905;
    wire N__35904;
    wire N__35903;
    wire N__35902;
    wire N__35901;
    wire N__35900;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35896;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35885;
    wire N__35880;
    wire N__35871;
    wire N__35870;
    wire N__35867;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35854;
    wire N__35847;
    wire N__35844;
    wire N__35837;
    wire N__35834;
    wire N__35831;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35821;
    wire N__35820;
    wire N__35819;
    wire N__35816;
    wire N__35815;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35802;
    wire N__35797;
    wire N__35794;
    wire N__35789;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35775;
    wire N__35774;
    wire N__35769;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35746;
    wire N__35745;
    wire N__35744;
    wire N__35741;
    wire N__35736;
    wire N__35731;
    wire N__35726;
    wire N__35715;
    wire N__35710;
    wire N__35707;
    wire N__35702;
    wire N__35699;
    wire N__35684;
    wire N__35679;
    wire N__35656;
    wire N__35655;
    wire N__35654;
    wire N__35653;
    wire N__35652;
    wire N__35647;
    wire N__35640;
    wire N__35635;
    wire N__35632;
    wire N__35631;
    wire N__35630;
    wire N__35627;
    wire N__35622;
    wire N__35617;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35607;
    wire N__35604;
    wire N__35603;
    wire N__35600;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35574;
    wire N__35571;
    wire N__35570;
    wire N__35567;
    wire N__35566;
    wire N__35563;
    wire N__35558;
    wire N__35555;
    wire N__35548;
    wire N__35545;
    wire N__35544;
    wire N__35541;
    wire N__35540;
    wire N__35537;
    wire N__35530;
    wire N__35527;
    wire N__35526;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35448;
    wire N__35447;
    wire N__35444;
    wire N__35443;
    wire N__35440;
    wire N__35435;
    wire N__35432;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35383;
    wire N__35382;
    wire N__35381;
    wire N__35378;
    wire N__35377;
    wire N__35374;
    wire N__35369;
    wire N__35366;
    wire N__35359;
    wire N__35356;
    wire N__35355;
    wire N__35352;
    wire N__35351;
    wire N__35348;
    wire N__35341;
    wire N__35338;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35328;
    wire N__35323;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35263;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35217;
    wire N__35214;
    wire N__35213;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35203;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35182;
    wire N__35181;
    wire N__35180;
    wire N__35177;
    wire N__35176;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35162;
    wire N__35155;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35147;
    wire N__35140;
    wire N__35137;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35058;
    wire N__35057;
    wire N__35054;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35046;
    wire N__35045;
    wire N__35044;
    wire N__35043;
    wire N__35042;
    wire N__35041;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35024;
    wire N__35023;
    wire N__35022;
    wire N__35021;
    wire N__35020;
    wire N__35019;
    wire N__35018;
    wire N__35017;
    wire N__35016;
    wire N__35011;
    wire N__35008;
    wire N__35003;
    wire N__34996;
    wire N__34995;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34971;
    wire N__34964;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34944;
    wire N__34933;
    wire N__34930;
    wire N__34921;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34884;
    wire N__34883;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34871;
    wire N__34864;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34807;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34738;
    wire N__34735;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34723;
    wire N__34722;
    wire N__34721;
    wire N__34718;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34712;
    wire N__34711;
    wire N__34702;
    wire N__34697;
    wire N__34694;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34675;
    wire N__34674;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34662;
    wire N__34661;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34645;
    wire N__34644;
    wire N__34641;
    wire N__34638;
    wire N__34633;
    wire N__34630;
    wire N__34627;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34607;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34573;
    wire N__34570;
    wire N__34567;
    wire N__34564;
    wire N__34563;
    wire N__34558;
    wire N__34555;
    wire N__34552;
    wire N__34549;
    wire N__34546;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34536;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34518;
    wire N__34513;
    wire N__34512;
    wire N__34507;
    wire N__34504;
    wire N__34501;
    wire N__34498;
    wire N__34495;
    wire N__34492;
    wire N__34489;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34438;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34410;
    wire N__34409;
    wire N__34408;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34392;
    wire N__34387;
    wire N__34386;
    wire N__34381;
    wire N__34378;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34332;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34316;
    wire N__34311;
    wire N__34306;
    wire N__34303;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34260;
    wire N__34255;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34245;
    wire N__34242;
    wire N__34239;
    wire N__34236;
    wire N__34231;
    wire N__34228;
    wire N__34227;
    wire N__34224;
    wire N__34223;
    wire N__34220;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34204;
    wire N__34203;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34182;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34147;
    wire N__34144;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34125;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34095;
    wire N__34094;
    wire N__34091;
    wire N__34086;
    wire N__34083;
    wire N__34078;
    wire N__34075;
    wire N__34074;
    wire N__34073;
    wire N__34068;
    wire N__34065;
    wire N__34060;
    wire N__34059;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34044;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34030;
    wire N__34029;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33990;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33966;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33955;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33943;
    wire N__33940;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33918;
    wire N__33915;
    wire N__33914;
    wire N__33911;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33880;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33819;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33805;
    wire N__33802;
    wire N__33801;
    wire N__33798;
    wire N__33797;
    wire N__33796;
    wire N__33793;
    wire N__33792;
    wire N__33785;
    wire N__33784;
    wire N__33783;
    wire N__33782;
    wire N__33781;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33762;
    wire N__33759;
    wire N__33756;
    wire N__33755;
    wire N__33754;
    wire N__33749;
    wire N__33746;
    wire N__33743;
    wire N__33738;
    wire N__33735;
    wire N__33730;
    wire N__33729;
    wire N__33726;
    wire N__33725;
    wire N__33720;
    wire N__33715;
    wire N__33710;
    wire N__33705;
    wire N__33702;
    wire N__33691;
    wire N__33688;
    wire N__33687;
    wire N__33686;
    wire N__33685;
    wire N__33684;
    wire N__33683;
    wire N__33680;
    wire N__33675;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33650;
    wire N__33647;
    wire N__33644;
    wire N__33641;
    wire N__33634;
    wire N__33633;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33625;
    wire N__33622;
    wire N__33621;
    wire N__33618;
    wire N__33617;
    wire N__33614;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33601;
    wire N__33598;
    wire N__33597;
    wire N__33596;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33588;
    wire N__33587;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33566;
    wire N__33563;
    wire N__33558;
    wire N__33551;
    wire N__33544;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33439;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33367;
    wire N__33364;
    wire N__33363;
    wire N__33362;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33356;
    wire N__33355;
    wire N__33354;
    wire N__33353;
    wire N__33352;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33338;
    wire N__33335;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33317;
    wire N__33312;
    wire N__33309;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33290;
    wire N__33287;
    wire N__33282;
    wire N__33277;
    wire N__33262;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33120;
    wire N__33119;
    wire N__33116;
    wire N__33113;
    wire N__33110;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33087;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33051;
    wire N__33050;
    wire N__33047;
    wire N__33044;
    wire N__33041;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33018;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32984;
    wire N__32983;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32966;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32940;
    wire N__32939;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32923;
    wire N__32920;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32894;
    wire N__32889;
    wire N__32886;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32840;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32811;
    wire N__32808;
    wire N__32805;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32759;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32731;
    wire N__32728;
    wire N__32725;
    wire N__32722;
    wire N__32719;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32711;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32587;
    wire N__32586;
    wire N__32583;
    wire N__32582;
    wire N__32579;
    wire N__32578;
    wire N__32575;
    wire N__32570;
    wire N__32567;
    wire N__32560;
    wire N__32557;
    wire N__32556;
    wire N__32553;
    wire N__32552;
    wire N__32549;
    wire N__32548;
    wire N__32547;
    wire N__32546;
    wire N__32543;
    wire N__32540;
    wire N__32533;
    wire N__32530;
    wire N__32521;
    wire N__32520;
    wire N__32519;
    wire N__32516;
    wire N__32513;
    wire N__32510;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32498;
    wire N__32497;
    wire N__32494;
    wire N__32489;
    wire N__32486;
    wire N__32479;
    wire N__32476;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32463;
    wire N__32456;
    wire N__32453;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32439;
    wire N__32438;
    wire N__32437;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32422;
    wire N__32417;
    wire N__32410;
    wire N__32407;
    wire N__32404;
    wire N__32401;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32393;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32379;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32365;
    wire N__32362;
    wire N__32361;
    wire N__32358;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32340;
    wire N__32337;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32323;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32310;
    wire N__32307;
    wire N__32306;
    wire N__32303;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32253;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32232;
    wire N__32231;
    wire N__32228;
    wire N__32223;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32211;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32175;
    wire N__32174;
    wire N__32173;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32163;
    wire N__32160;
    wire N__32155;
    wire N__32150;
    wire N__32147;
    wire N__32144;
    wire N__32143;
    wire N__32142;
    wire N__32141;
    wire N__32140;
    wire N__32139;
    wire N__32136;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32096;
    wire N__32095;
    wire N__32094;
    wire N__32093;
    wire N__32092;
    wire N__32091;
    wire N__32090;
    wire N__32089;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32082;
    wire N__32077;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32057;
    wire N__32046;
    wire N__32037;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32015;
    wire N__32010;
    wire N__32007;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31987;
    wire N__31986;
    wire N__31981;
    wire N__31978;
    wire N__31977;
    wire N__31976;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31945;
    wire N__31942;
    wire N__31941;
    wire N__31940;
    wire N__31939;
    wire N__31934;
    wire N__31929;
    wire N__31928;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31912;
    wire N__31911;
    wire N__31910;
    wire N__31909;
    wire N__31908;
    wire N__31907;
    wire N__31900;
    wire N__31897;
    wire N__31888;
    wire N__31887;
    wire N__31886;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31881;
    wire N__31880;
    wire N__31875;
    wire N__31874;
    wire N__31873;
    wire N__31872;
    wire N__31871;
    wire N__31870;
    wire N__31865;
    wire N__31858;
    wire N__31849;
    wire N__31840;
    wire N__31837;
    wire N__31836;
    wire N__31835;
    wire N__31828;
    wire N__31823;
    wire N__31820;
    wire N__31813;
    wire N__31810;
    wire N__31805;
    wire N__31800;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31739;
    wire N__31736;
    wire N__31731;
    wire N__31730;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31706;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31690;
    wire N__31689;
    wire N__31686;
    wire N__31685;
    wire N__31682;
    wire N__31681;
    wire N__31678;
    wire N__31673;
    wire N__31670;
    wire N__31663;
    wire N__31660;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31648;
    wire N__31647;
    wire N__31644;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31632;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31599;
    wire N__31596;
    wire N__31595;
    wire N__31592;
    wire N__31587;
    wire N__31582;
    wire N__31581;
    wire N__31576;
    wire N__31573;
    wire N__31570;
    wire N__31567;
    wire N__31564;
    wire N__31561;
    wire N__31560;
    wire N__31557;
    wire N__31556;
    wire N__31555;
    wire N__31552;
    wire N__31549;
    wire N__31548;
    wire N__31543;
    wire N__31540;
    wire N__31537;
    wire N__31534;
    wire N__31525;
    wire N__31524;
    wire N__31523;
    wire N__31522;
    wire N__31521;
    wire N__31520;
    wire N__31519;
    wire N__31518;
    wire N__31517;
    wire N__31514;
    wire N__31511;
    wire N__31502;
    wire N__31495;
    wire N__31494;
    wire N__31493;
    wire N__31492;
    wire N__31491;
    wire N__31488;
    wire N__31481;
    wire N__31478;
    wire N__31471;
    wire N__31466;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31411;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31372;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31324;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31251;
    wire N__31250;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31238;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31215;
    wire N__31214;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31177;
    wire N__31176;
    wire N__31173;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31159;
    wire N__31156;
    wire N__31153;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31132;
    wire N__31131;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31085;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31038;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31014;
    wire N__31013;
    wire N__31010;
    wire N__31005;
    wire N__31004;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30988;
    wire N__30987;
    wire N__30986;
    wire N__30985;
    wire N__30982;
    wire N__30981;
    wire N__30980;
    wire N__30979;
    wire N__30978;
    wire N__30977;
    wire N__30976;
    wire N__30975;
    wire N__30974;
    wire N__30973;
    wire N__30970;
    wire N__30961;
    wire N__30960;
    wire N__30959;
    wire N__30958;
    wire N__30957;
    wire N__30956;
    wire N__30953;
    wire N__30952;
    wire N__30951;
    wire N__30950;
    wire N__30945;
    wire N__30938;
    wire N__30933;
    wire N__30928;
    wire N__30927;
    wire N__30924;
    wire N__30917;
    wire N__30916;
    wire N__30913;
    wire N__30912;
    wire N__30909;
    wire N__30902;
    wire N__30899;
    wire N__30892;
    wire N__30887;
    wire N__30884;
    wire N__30877;
    wire N__30862;
    wire N__30861;
    wire N__30860;
    wire N__30859;
    wire N__30858;
    wire N__30857;
    wire N__30856;
    wire N__30855;
    wire N__30854;
    wire N__30853;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30844;
    wire N__30843;
    wire N__30842;
    wire N__30835;
    wire N__30828;
    wire N__30821;
    wire N__30816;
    wire N__30815;
    wire N__30814;
    wire N__30813;
    wire N__30812;
    wire N__30811;
    wire N__30804;
    wire N__30801;
    wire N__30796;
    wire N__30791;
    wire N__30780;
    wire N__30777;
    wire N__30766;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30745;
    wire N__30742;
    wire N__30739;
    wire N__30736;
    wire N__30733;
    wire N__30732;
    wire N__30731;
    wire N__30730;
    wire N__30727;
    wire N__30726;
    wire N__30725;
    wire N__30724;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30711;
    wire N__30710;
    wire N__30709;
    wire N__30708;
    wire N__30707;
    wire N__30702;
    wire N__30701;
    wire N__30700;
    wire N__30699;
    wire N__30698;
    wire N__30697;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30680;
    wire N__30677;
    wire N__30672;
    wire N__30665;
    wire N__30662;
    wire N__30661;
    wire N__30660;
    wire N__30655;
    wire N__30644;
    wire N__30639;
    wire N__30634;
    wire N__30629;
    wire N__30626;
    wire N__30617;
    wire N__30612;
    wire N__30605;
    wire N__30592;
    wire N__30591;
    wire N__30590;
    wire N__30589;
    wire N__30588;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30540;
    wire N__30537;
    wire N__30536;
    wire N__30535;
    wire N__30532;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30516;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30489;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30471;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30438;
    wire N__30437;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30416;
    wire N__30413;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30399;
    wire N__30398;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30366;
    wire N__30365;
    wire N__30360;
    wire N__30357;
    wire N__30352;
    wire N__30349;
    wire N__30348;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30321;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30298;
    wire N__30297;
    wire N__30296;
    wire N__30295;
    wire N__30292;
    wire N__30291;
    wire N__30288;
    wire N__30287;
    wire N__30284;
    wire N__30283;
    wire N__30280;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30246;
    wire N__30243;
    wire N__30242;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30206;
    wire N__30203;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30139;
    wire N__30136;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30087;
    wire N__30086;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30010;
    wire N__30007;
    wire N__30006;
    wire N__30005;
    wire N__30000;
    wire N__29997;
    wire N__29992;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29980;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29923;
    wire N__29922;
    wire N__29921;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29906;
    wire N__29901;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29883;
    wire N__29880;
    wire N__29879;
    wire N__29878;
    wire N__29877;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29863;
    wire N__29856;
    wire N__29851;
    wire N__29846;
    wire N__29839;
    wire N__29838;
    wire N__29837;
    wire N__29836;
    wire N__29833;
    wire N__29832;
    wire N__29829;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29813;
    wire N__29806;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29779;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29771;
    wire N__29766;
    wire N__29761;
    wire N__29758;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29737;
    wire N__29736;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29730;
    wire N__29727;
    wire N__29726;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29713;
    wire N__29710;
    wire N__29707;
    wire N__29706;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29680;
    wire N__29677;
    wire N__29670;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29613;
    wire N__29612;
    wire N__29609;
    wire N__29608;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29594;
    wire N__29591;
    wire N__29590;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29560;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29538;
    wire N__29537;
    wire N__29536;
    wire N__29535;
    wire N__29534;
    wire N__29533;
    wire N__29532;
    wire N__29531;
    wire N__29530;
    wire N__29527;
    wire N__29526;
    wire N__29525;
    wire N__29524;
    wire N__29519;
    wire N__29518;
    wire N__29517;
    wire N__29516;
    wire N__29513;
    wire N__29510;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29499;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29491;
    wire N__29490;
    wire N__29483;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29449;
    wire N__29446;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29426;
    wire N__29417;
    wire N__29410;
    wire N__29401;
    wire N__29400;
    wire N__29399;
    wire N__29398;
    wire N__29397;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29379;
    wire N__29376;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29348;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29334;
    wire N__29331;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29314;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29285;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29223;
    wire N__29220;
    wire N__29219;
    wire N__29218;
    wire N__29217;
    wire N__29216;
    wire N__29215;
    wire N__29212;
    wire N__29209;
    wire N__29204;
    wire N__29201;
    wire N__29200;
    wire N__29199;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29191;
    wire N__29190;
    wire N__29189;
    wire N__29186;
    wire N__29181;
    wire N__29178;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29157;
    wire N__29152;
    wire N__29143;
    wire N__29134;
    wire N__29131;
    wire N__29130;
    wire N__29129;
    wire N__29128;
    wire N__29125;
    wire N__29120;
    wire N__29117;
    wire N__29116;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29102;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29088;
    wire N__29083;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29046;
    wire N__29041;
    wire N__29038;
    wire N__29037;
    wire N__29034;
    wire N__29033;
    wire N__29030;
    wire N__29029;
    wire N__29028;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29015;
    wire N__29012;
    wire N__29009;
    wire N__29006;
    wire N__29005;
    wire N__29002;
    wire N__29001;
    wire N__29000;
    wire N__28997;
    wire N__28994;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28965;
    wire N__28960;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28899;
    wire N__28898;
    wire N__28897;
    wire N__28896;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28886;
    wire N__28883;
    wire N__28882;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28865;
    wire N__28860;
    wire N__28855;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28830;
    wire N__28829;
    wire N__28826;
    wire N__28825;
    wire N__28822;
    wire N__28817;
    wire N__28814;
    wire N__28807;
    wire N__28804;
    wire N__28803;
    wire N__28800;
    wire N__28799;
    wire N__28796;
    wire N__28789;
    wire N__28786;
    wire N__28785;
    wire N__28784;
    wire N__28781;
    wire N__28776;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28759;
    wire N__28758;
    wire N__28757;
    wire N__28756;
    wire N__28755;
    wire N__28754;
    wire N__28751;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28730;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28708;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28506;
    wire N__28503;
    wire N__28502;
    wire N__28499;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28446;
    wire N__28443;
    wire N__28442;
    wire N__28439;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28386;
    wire N__28385;
    wire N__28382;
    wire N__28379;
    wire N__28374;
    wire N__28371;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28142;
    wire N__28139;
    wire N__28136;
    wire N__28133;
    wire N__28126;
    wire N__28125;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28096;
    wire N__28095;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28060;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28035;
    wire N__28030;
    wire N__28027;
    wire N__28026;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28009;
    wire N__28008;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27976;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27937;
    wire N__27934;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27903;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27893;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27877;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27849;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27820;
    wire N__27819;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27790;
    wire N__27787;
    wire N__27786;
    wire N__27781;
    wire N__27778;
    wire N__27775;
    wire N__27772;
    wire N__27769;
    wire N__27766;
    wire N__27763;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27748;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27736;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27723;
    wire N__27722;
    wire N__27721;
    wire N__27720;
    wire N__27719;
    wire N__27718;
    wire N__27715;
    wire N__27714;
    wire N__27711;
    wire N__27710;
    wire N__27707;
    wire N__27702;
    wire N__27701;
    wire N__27700;
    wire N__27695;
    wire N__27692;
    wire N__27689;
    wire N__27688;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27676;
    wire N__27673;
    wire N__27672;
    wire N__27671;
    wire N__27670;
    wire N__27669;
    wire N__27668;
    wire N__27665;
    wire N__27664;
    wire N__27663;
    wire N__27660;
    wire N__27659;
    wire N__27658;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27646;
    wire N__27639;
    wire N__27634;
    wire N__27629;
    wire N__27624;
    wire N__27617;
    wire N__27614;
    wire N__27607;
    wire N__27604;
    wire N__27603;
    wire N__27596;
    wire N__27595;
    wire N__27586;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27569;
    wire N__27564;
    wire N__27553;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27538;
    wire N__27535;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27511;
    wire N__27510;
    wire N__27505;
    wire N__27502;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27472;
    wire N__27469;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27456;
    wire N__27455;
    wire N__27454;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27450;
    wire N__27449;
    wire N__27448;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27438;
    wire N__27437;
    wire N__27430;
    wire N__27421;
    wire N__27420;
    wire N__27419;
    wire N__27418;
    wire N__27415;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27395;
    wire N__27392;
    wire N__27389;
    wire N__27382;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27352;
    wire N__27351;
    wire N__27350;
    wire N__27349;
    wire N__27348;
    wire N__27345;
    wire N__27340;
    wire N__27335;
    wire N__27332;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27252;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27234;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27216;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27177;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27150;
    wire N__27149;
    wire N__27148;
    wire N__27147;
    wire N__27146;
    wire N__27143;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27130;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27109;
    wire N__27108;
    wire N__27105;
    wire N__27104;
    wire N__27103;
    wire N__27102;
    wire N__27101;
    wire N__27100;
    wire N__27097;
    wire N__27096;
    wire N__27093;
    wire N__27092;
    wire N__27089;
    wire N__27088;
    wire N__27085;
    wire N__27082;
    wire N__27079;
    wire N__27078;
    wire N__27075;
    wire N__27070;
    wire N__27065;
    wire N__27064;
    wire N__27063;
    wire N__27060;
    wire N__27059;
    wire N__27058;
    wire N__27055;
    wire N__27054;
    wire N__27051;
    wire N__27034;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27018;
    wire N__27015;
    wire N__27010;
    wire N__26999;
    wire N__26992;
    wire N__26977;
    wire N__26976;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26944;
    wire N__26943;
    wire N__26942;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26904;
    wire N__26899;
    wire N__26896;
    wire N__26887;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26876;
    wire N__26873;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26861;
    wire N__26854;
    wire N__26853;
    wire N__26848;
    wire N__26845;
    wire N__26844;
    wire N__26843;
    wire N__26842;
    wire N__26839;
    wire N__26838;
    wire N__26837;
    wire N__26836;
    wire N__26835;
    wire N__26834;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26812;
    wire N__26809;
    wire N__26808;
    wire N__26801;
    wire N__26800;
    wire N__26799;
    wire N__26798;
    wire N__26795;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26789;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26777;
    wire N__26776;
    wire N__26773;
    wire N__26768;
    wire N__26763;
    wire N__26760;
    wire N__26751;
    wire N__26750;
    wire N__26745;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26726;
    wire N__26723;
    wire N__26718;
    wire N__26713;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26693;
    wire N__26688;
    wire N__26685;
    wire N__26680;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26649;
    wire N__26648;
    wire N__26647;
    wire N__26646;
    wire N__26645;
    wire N__26644;
    wire N__26643;
    wire N__26642;
    wire N__26641;
    wire N__26638;
    wire N__26637;
    wire N__26636;
    wire N__26635;
    wire N__26634;
    wire N__26633;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26616;
    wire N__26613;
    wire N__26612;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26587;
    wire N__26584;
    wire N__26579;
    wire N__26576;
    wire N__26571;
    wire N__26570;
    wire N__26569;
    wire N__26568;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26552;
    wire N__26547;
    wire N__26542;
    wire N__26539;
    wire N__26534;
    wire N__26531;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26508;
    wire N__26505;
    wire N__26496;
    wire N__26489;
    wire N__26482;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26470;
    wire N__26467;
    wire N__26466;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26451;
    wire N__26450;
    wire N__26449;
    wire N__26448;
    wire N__26447;
    wire N__26446;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26438;
    wire N__26437;
    wire N__26436;
    wire N__26435;
    wire N__26434;
    wire N__26433;
    wire N__26432;
    wire N__26427;
    wire N__26426;
    wire N__26425;
    wire N__26422;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26398;
    wire N__26391;
    wire N__26388;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26335;
    wire N__26334;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26328;
    wire N__26327;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26310;
    wire N__26309;
    wire N__26308;
    wire N__26305;
    wire N__26302;
    wire N__26301;
    wire N__26300;
    wire N__26299;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26280;
    wire N__26277;
    wire N__26276;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26233;
    wire N__26228;
    wire N__26221;
    wire N__26206;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26196;
    wire N__26193;
    wire N__26192;
    wire N__26191;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26171;
    wire N__26168;
    wire N__26167;
    wire N__26166;
    wire N__26165;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26153;
    wire N__26148;
    wire N__26145;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26125;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26107;
    wire N__26104;
    wire N__26103;
    wire N__26102;
    wire N__26099;
    wire N__26096;
    wire N__26087;
    wire N__26084;
    wire N__26077;
    wire N__26072;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26004;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25989;
    wire N__25984;
    wire N__25981;
    wire N__25980;
    wire N__25977;
    wire N__25976;
    wire N__25973;
    wire N__25972;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25948;
    wire N__25947;
    wire N__25946;
    wire N__25945;
    wire N__25938;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25916;
    wire N__25909;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25897;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25873;
    wire N__25872;
    wire N__25867;
    wire N__25864;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25859;
    wire N__25858;
    wire N__25857;
    wire N__25854;
    wire N__25853;
    wire N__25844;
    wire N__25841;
    wire N__25840;
    wire N__25839;
    wire N__25838;
    wire N__25837;
    wire N__25836;
    wire N__25835;
    wire N__25834;
    wire N__25831;
    wire N__25830;
    wire N__25827;
    wire N__25826;
    wire N__25825;
    wire N__25824;
    wire N__25823;
    wire N__25820;
    wire N__25819;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25815;
    wire N__25812;
    wire N__25811;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25789;
    wire N__25786;
    wire N__25777;
    wire N__25772;
    wire N__25769;
    wire N__25758;
    wire N__25753;
    wire N__25746;
    wire N__25739;
    wire N__25736;
    wire N__25723;
    wire N__25720;
    wire N__25719;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25704;
    wire N__25699;
    wire N__25696;
    wire N__25693;
    wire N__25690;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25593;
    wire N__25590;
    wire N__25589;
    wire N__25586;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25544;
    wire N__25539;
    wire N__25534;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25518;
    wire N__25517;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25505;
    wire N__25500;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25475;
    wire N__25474;
    wire N__25473;
    wire N__25470;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25372;
    wire N__25369;
    wire N__25366;
    wire N__25365;
    wire N__25364;
    wire N__25357;
    wire N__25354;
    wire N__25353;
    wire N__25352;
    wire N__25351;
    wire N__25348;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25340;
    wire N__25337;
    wire N__25336;
    wire N__25325;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25291;
    wire N__25290;
    wire N__25289;
    wire N__25288;
    wire N__25287;
    wire N__25286;
    wire N__25285;
    wire N__25280;
    wire N__25269;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25239;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25210;
    wire N__25209;
    wire N__25208;
    wire N__25207;
    wire N__25206;
    wire N__25205;
    wire N__25204;
    wire N__25203;
    wire N__25202;
    wire N__25199;
    wire N__25192;
    wire N__25185;
    wire N__25178;
    wire N__25169;
    wire N__25162;
    wire N__25159;
    wire N__25158;
    wire N__25157;
    wire N__25156;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25008;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24984;
    wire N__24979;
    wire N__24976;
    wire N__24973;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24963;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24933;
    wire N__24932;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24924;
    wire N__24921;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24901;
    wire N__24900;
    wire N__24895;
    wire N__24890;
    wire N__24885;
    wire N__24880;
    wire N__24875;
    wire N__24872;
    wire N__24865;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24857;
    wire N__24850;
    wire N__24849;
    wire N__24846;
    wire N__24845;
    wire N__24842;
    wire N__24841;
    wire N__24840;
    wire N__24839;
    wire N__24838;
    wire N__24837;
    wire N__24836;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24815;
    wire N__24810;
    wire N__24805;
    wire N__24802;
    wire N__24797;
    wire N__24794;
    wire N__24787;
    wire N__24784;
    wire N__24783;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24756;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24738;
    wire N__24735;
    wire N__24732;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24720;
    wire N__24717;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24690;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24669;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24657;
    wire N__24654;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24642;
    wire N__24641;
    wire N__24640;
    wire N__24639;
    wire N__24638;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24626;
    wire N__24623;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24607;
    wire N__24606;
    wire N__24605;
    wire N__24604;
    wire N__24601;
    wire N__24596;
    wire N__24593;
    wire N__24588;
    wire N__24587;
    wire N__24586;
    wire N__24583;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24562;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24539;
    wire N__24536;
    wire N__24531;
    wire N__24520;
    wire N__24519;
    wire N__24516;
    wire N__24515;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24511;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24500;
    wire N__24497;
    wire N__24494;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24473;
    wire N__24470;
    wire N__24469;
    wire N__24466;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24429;
    wire N__24426;
    wire N__24415;
    wire N__24410;
    wire N__24405;
    wire N__24400;
    wire N__24397;
    wire N__24396;
    wire N__24395;
    wire N__24394;
    wire N__24393;
    wire N__24392;
    wire N__24391;
    wire N__24390;
    wire N__24389;
    wire N__24388;
    wire N__24387;
    wire N__24376;
    wire N__24371;
    wire N__24370;
    wire N__24367;
    wire N__24366;
    wire N__24365;
    wire N__24362;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24331;
    wire N__24330;
    wire N__24329;
    wire N__24328;
    wire N__24325;
    wire N__24320;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24314;
    wire N__24309;
    wire N__24308;
    wire N__24305;
    wire N__24300;
    wire N__24297;
    wire N__24290;
    wire N__24285;
    wire N__24278;
    wire N__24275;
    wire N__24272;
    wire N__24269;
    wire N__24266;
    wire N__24259;
    wire N__24254;
    wire N__24251;
    wire N__24246;
    wire N__24241;
    wire N__24238;
    wire N__24233;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24213;
    wire N__24212;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24191;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24166;
    wire N__24163;
    wire N__24162;
    wire N__24161;
    wire N__24156;
    wire N__24155;
    wire N__24152;
    wire N__24151;
    wire N__24150;
    wire N__24149;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24133;
    wire N__24132;
    wire N__24129;
    wire N__24128;
    wire N__24127;
    wire N__24126;
    wire N__24125;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24113;
    wire N__24112;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24104;
    wire N__24103;
    wire N__24102;
    wire N__24101;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24086;
    wire N__24083;
    wire N__24076;
    wire N__24073;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24056;
    wire N__24053;
    wire N__24052;
    wire N__24047;
    wire N__24040;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24025;
    wire N__24022;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24000;
    wire N__23995;
    wire N__23992;
    wire N__23991;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23956;
    wire N__23953;
    wire N__23950;
    wire N__23947;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23934;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23919;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23907;
    wire N__23906;
    wire N__23905;
    wire N__23904;
    wire N__23903;
    wire N__23900;
    wire N__23899;
    wire N__23896;
    wire N__23895;
    wire N__23894;
    wire N__23891;
    wire N__23888;
    wire N__23887;
    wire N__23886;
    wire N__23881;
    wire N__23880;
    wire N__23879;
    wire N__23878;
    wire N__23877;
    wire N__23876;
    wire N__23875;
    wire N__23874;
    wire N__23871;
    wire N__23866;
    wire N__23861;
    wire N__23858;
    wire N__23857;
    wire N__23854;
    wire N__23853;
    wire N__23852;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23837;
    wire N__23836;
    wire N__23835;
    wire N__23830;
    wire N__23825;
    wire N__23822;
    wire N__23817;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23793;
    wire N__23792;
    wire N__23789;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23767;
    wire N__23758;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23738;
    wire N__23735;
    wire N__23722;
    wire N__23721;
    wire N__23720;
    wire N__23717;
    wire N__23716;
    wire N__23715;
    wire N__23714;
    wire N__23711;
    wire N__23710;
    wire N__23709;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23703;
    wire N__23702;
    wire N__23701;
    wire N__23700;
    wire N__23699;
    wire N__23698;
    wire N__23697;
    wire N__23696;
    wire N__23695;
    wire N__23694;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23673;
    wire N__23672;
    wire N__23671;
    wire N__23664;
    wire N__23657;
    wire N__23656;
    wire N__23655;
    wire N__23650;
    wire N__23647;
    wire N__23640;
    wire N__23639;
    wire N__23638;
    wire N__23633;
    wire N__23632;
    wire N__23619;
    wire N__23618;
    wire N__23617;
    wire N__23612;
    wire N__23607;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23588;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23573;
    wire N__23568;
    wire N__23563;
    wire N__23560;
    wire N__23555;
    wire N__23552;
    wire N__23533;
    wire N__23532;
    wire N__23531;
    wire N__23528;
    wire N__23525;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23519;
    wire N__23514;
    wire N__23511;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23472;
    wire N__23469;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23452;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23430;
    wire N__23427;
    wire N__23426;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23395;
    wire N__23392;
    wire N__23391;
    wire N__23390;
    wire N__23389;
    wire N__23388;
    wire N__23383;
    wire N__23382;
    wire N__23381;
    wire N__23380;
    wire N__23377;
    wire N__23376;
    wire N__23375;
    wire N__23370;
    wire N__23367;
    wire N__23366;
    wire N__23365;
    wire N__23360;
    wire N__23357;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23305;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23275;
    wire N__23272;
    wire N__23271;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23241;
    wire N__23236;
    wire N__23235;
    wire N__23234;
    wire N__23233;
    wire N__23232;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23226;
    wire N__23221;
    wire N__23216;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23200;
    wire N__23195;
    wire N__23192;
    wire N__23187;
    wire N__23182;
    wire N__23181;
    wire N__23180;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23174;
    wire N__23173;
    wire N__23168;
    wire N__23167;
    wire N__23166;
    wire N__23165;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23157;
    wire N__23154;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23136;
    wire N__23133;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23102;
    wire N__23099;
    wire N__23092;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23076;
    wire N__23071;
    wire N__23068;
    wire N__23067;
    wire N__23066;
    wire N__23065;
    wire N__23062;
    wire N__23061;
    wire N__23060;
    wire N__23059;
    wire N__23058;
    wire N__23057;
    wire N__23056;
    wire N__23055;
    wire N__23054;
    wire N__23053;
    wire N__23052;
    wire N__23051;
    wire N__23048;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23044;
    wire N__23043;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23027;
    wire N__23026;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23012;
    wire N__23005;
    wire N__23002;
    wire N__22997;
    wire N__22992;
    wire N__22991;
    wire N__22988;
    wire N__22987;
    wire N__22986;
    wire N__22983;
    wire N__22976;
    wire N__22971;
    wire N__22968;
    wire N__22961;
    wire N__22954;
    wire N__22947;
    wire N__22944;
    wire N__22937;
    wire N__22930;
    wire N__22925;
    wire N__22922;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22908;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22885;
    wire N__22882;
    wire N__22881;
    wire N__22880;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22857;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22813;
    wire N__22810;
    wire N__22809;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22797;
    wire N__22792;
    wire N__22789;
    wire N__22788;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22770;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22672;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22600;
    wire N__22597;
    wire N__22596;
    wire N__22595;
    wire N__22590;
    wire N__22587;
    wire N__22582;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22558;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22536;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22497;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22398;
    wire N__22397;
    wire N__22394;
    wire N__22393;
    wire N__22390;
    wire N__22383;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22329;
    wire N__22326;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22318;
    wire N__22317;
    wire N__22314;
    wire N__22313;
    wire N__22312;
    wire N__22311;
    wire N__22310;
    wire N__22309;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22278;
    wire N__22273;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22230;
    wire N__22229;
    wire N__22228;
    wire N__22227;
    wire N__22220;
    wire N__22215;
    wire N__22210;
    wire N__22207;
    wire N__22206;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22187;
    wire N__22186;
    wire N__22181;
    wire N__22176;
    wire N__22169;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22119;
    wire N__22116;
    wire N__22115;
    wire N__22114;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22104;
    wire N__22099;
    wire N__22098;
    wire N__22097;
    wire N__22096;
    wire N__22095;
    wire N__22094;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22074;
    wire N__22067;
    wire N__22066;
    wire N__22065;
    wire N__22060;
    wire N__22055;
    wire N__22050;
    wire N__22045;
    wire N__22036;
    wire N__22035;
    wire N__22032;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22021;
    wire N__22018;
    wire N__22013;
    wire N__22010;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__21998;
    wire N__21991;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21979;
    wire N__21978;
    wire N__21977;
    wire N__21974;
    wire N__21969;
    wire N__21966;
    wire N__21959;
    wire N__21956;
    wire N__21951;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21939;
    wire N__21936;
    wire N__21933;
    wire N__21928;
    wire N__21927;
    wire N__21926;
    wire N__21925;
    wire N__21924;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21904;
    wire N__21903;
    wire N__21902;
    wire N__21901;
    wire N__21900;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21876;
    wire N__21875;
    wire N__21874;
    wire N__21871;
    wire N__21870;
    wire N__21869;
    wire N__21858;
    wire N__21857;
    wire N__21854;
    wire N__21853;
    wire N__21850;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21819;
    wire N__21814;
    wire N__21813;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21798;
    wire N__21795;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21754;
    wire N__21751;
    wire N__21750;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21735;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21720;
    wire N__21715;
    wire N__21712;
    wire N__21711;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21699;
    wire N__21694;
    wire N__21691;
    wire N__21690;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21651;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21612;
    wire N__21607;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21599;
    wire N__21594;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21549;
    wire N__21546;
    wire N__21545;
    wire N__21542;
    wire N__21537;
    wire N__21534;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21522;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21472;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21457;
    wire N__21456;
    wire N__21451;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21420;
    wire N__21419;
    wire N__21414;
    wire N__21413;
    wire N__21410;
    wire N__21407;
    wire N__21406;
    wire N__21403;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21391;
    wire N__21388;
    wire N__21379;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21328;
    wire N__21325;
    wire N__21324;
    wire N__21323;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21265;
    wire N__21262;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21243;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21225;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21202;
    wire N__21201;
    wire N__21200;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21177;
    wire N__21174;
    wire N__21169;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21161;
    wire N__21154;
    wire N__21149;
    wire N__21142;
    wire N__21141;
    wire N__21140;
    wire N__21139;
    wire N__21138;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21097;
    wire N__21096;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21061;
    wire N__21058;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21012;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20949;
    wire N__20946;
    wire N__20945;
    wire N__20944;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20929;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20915;
    wire N__20914;
    wire N__20913;
    wire N__20912;
    wire N__20911;
    wire N__20910;
    wire N__20907;
    wire N__20902;
    wire N__20897;
    wire N__20890;
    wire N__20883;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20859;
    wire N__20856;
    wire N__20849;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20820;
    wire N__20809;
    wire N__20800;
    wire N__20799;
    wire N__20798;
    wire N__20797;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20789;
    wire N__20786;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20750;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20707;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20699;
    wire N__20698;
    wire N__20697;
    wire N__20696;
    wire N__20695;
    wire N__20694;
    wire N__20693;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20675;
    wire N__20670;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20611;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20593;
    wire N__20590;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20562;
    wire N__20559;
    wire N__20556;
    wire N__20551;
    wire N__20550;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20535;
    wire N__20530;
    wire N__20527;
    wire N__20524;
    wire N__20521;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20497;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20458;
    wire N__20457;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20439;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20392;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20374;
    wire N__20371;
    wire N__20370;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20350;
    wire N__20347;
    wire N__20346;
    wire N__20343;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20331;
    wire N__20326;
    wire N__20323;
    wire N__20322;
    wire N__20319;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20289;
    wire N__20288;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20260;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20248;
    wire N__20243;
    wire N__20236;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20215;
    wire N__20212;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20202;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20146;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20134;
    wire N__20131;
    wire N__20128;
    wire N__20125;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20083;
    wire N__20082;
    wire N__20081;
    wire N__20078;
    wire N__20073;
    wire N__20070;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20040;
    wire N__20039;
    wire N__20038;
    wire N__20035;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20021;
    wire N__20016;
    wire N__20013;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19989;
    wire N__19988;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19965;
    wire N__19964;
    wire N__19959;
    wire N__19956;
    wire N__19951;
    wire N__19948;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19849;
    wire N__19848;
    wire N__19847;
    wire N__19844;
    wire N__19843;
    wire N__19842;
    wire N__19841;
    wire N__19840;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19815;
    wire N__19814;
    wire N__19813;
    wire N__19808;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19762;
    wire N__19761;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19728;
    wire N__19727;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19715;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19699;
    wire N__19696;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19668;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19624;
    wire N__19623;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19582;
    wire N__19579;
    wire N__19578;
    wire N__19573;
    wire N__19570;
    wire N__19567;
    wire N__19564;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19549;
    wire N__19548;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19536;
    wire N__19535;
    wire N__19534;
    wire N__19533;
    wire N__19532;
    wire N__19531;
    wire N__19530;
    wire N__19527;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19521;
    wire N__19520;
    wire N__19519;
    wire N__19518;
    wire N__19517;
    wire N__19516;
    wire N__19515;
    wire N__19510;
    wire N__19503;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19491;
    wire N__19490;
    wire N__19489;
    wire N__19488;
    wire N__19487;
    wire N__19486;
    wire N__19485;
    wire N__19484;
    wire N__19481;
    wire N__19476;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19458;
    wire N__19455;
    wire N__19450;
    wire N__19447;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19431;
    wire N__19428;
    wire N__19421;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19402;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19384;
    wire N__19379;
    wire N__19374;
    wire N__19363;
    wire N__19362;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19350;
    wire N__19349;
    wire N__19348;
    wire N__19347;
    wire N__19344;
    wire N__19343;
    wire N__19342;
    wire N__19341;
    wire N__19340;
    wire N__19339;
    wire N__19338;
    wire N__19337;
    wire N__19336;
    wire N__19335;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19325;
    wire N__19324;
    wire N__19323;
    wire N__19322;
    wire N__19321;
    wire N__19320;
    wire N__19319;
    wire N__19318;
    wire N__19317;
    wire N__19310;
    wire N__19305;
    wire N__19302;
    wire N__19293;
    wire N__19286;
    wire N__19273;
    wire N__19260;
    wire N__19245;
    wire N__19240;
    wire N__19229;
    wire N__19224;
    wire N__19221;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19174;
    wire N__19173;
    wire N__19168;
    wire N__19165;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19153;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19145;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19092;
    wire N__19089;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19051;
    wire N__19050;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18990;
    wire N__18985;
    wire N__18982;
    wire N__18981;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18969;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18942;
    wire N__18937;
    wire N__18934;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18922;
    wire N__18921;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18853;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18841;
    wire N__18840;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18817;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18741;
    wire N__18740;
    wire N__18737;
    wire N__18736;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18718;
    wire N__18717;
    wire N__18714;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18672;
    wire N__18669;
    wire N__18668;
    wire N__18665;
    wire N__18662;
    wire N__18659;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18636;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18592;
    wire N__18591;
    wire N__18588;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18571;
    wire N__18568;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18556;
    wire N__18555;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18532;
    wire N__18531;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18505;
    wire N__18502;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18450;
    wire N__18447;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18435;
    wire N__18430;
    wire N__18429;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18396;
    wire N__18391;
    wire N__18388;
    wire N__18385;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18360;
    wire N__18357;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18322;
    wire N__18321;
    wire N__18320;
    wire N__18317;
    wire N__18316;
    wire N__18313;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18288;
    wire N__18283;
    wire N__18280;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18258;
    wire N__18257;
    wire N__18256;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18232;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18154;
    wire N__18151;
    wire N__18148;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18111;
    wire N__18108;
    wire N__18107;
    wire N__18106;
    wire N__18103;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18095;
    wire N__18092;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18069;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18051;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18021;
    wire N__18018;
    wire N__18011;
    wire N__18006;
    wire N__18003;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17967;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17946;
    wire N__17943;
    wire N__17938;
    wire N__17933;
    wire N__17926;
    wire N__17923;
    wire N__17922;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17904;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17875;
    wire N__17874;
    wire N__17871;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17842;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17809;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17797;
    wire N__17794;
    wire N__17787;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17775;
    wire N__17772;
    wire N__17767;
    wire N__17764;
    wire N__17763;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17751;
    wire N__17750;
    wire N__17747;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17741;
    wire N__17740;
    wire N__17737;
    wire N__17736;
    wire N__17731;
    wire N__17728;
    wire N__17727;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17685;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17661;
    wire N__17658;
    wire N__17657;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17553;
    wire N__17552;
    wire N__17549;
    wire N__17544;
    wire N__17539;
    wire N__17538;
    wire N__17535;
    wire N__17532;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17493;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17418;
    wire N__17413;
    wire N__17410;
    wire N__17409;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17328;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17256;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17165;
    wire N__17160;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17095;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17083;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire N__17068;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17038;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17026;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17011;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__16999;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16888;
    wire N__16887;
    wire N__16886;
    wire N__16885;
    wire N__16884;
    wire N__16881;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16877;
    wire N__16876;
    wire N__16875;
    wire N__16874;
    wire N__16873;
    wire N__16872;
    wire N__16871;
    wire N__16870;
    wire N__16869;
    wire N__16868;
    wire N__16867;
    wire N__16866;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16852;
    wire N__16845;
    wire N__16838;
    wire N__16831;
    wire N__16816;
    wire N__16809;
    wire N__16798;
    wire N__16795;
    wire N__16794;
    wire N__16791;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16768;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16756;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16741;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16729;
    wire N__16728;
    wire N__16725;
    wire N__16722;
    wire N__16717;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16705;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16690;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16678;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16666;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16654;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16639;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16627;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16615;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16603;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16588;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16576;
    wire N__16573;
    wire N__16572;
    wire N__16569;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16555;
    wire N__16552;
    wire N__16543;
    wire N__16542;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16512;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16489;
    wire N__16486;
    wire N__16485;
    wire N__16480;
    wire N__16477;
    wire N__16474;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16462;
    wire N__16461;
    wire N__16456;
    wire N__16453;
    wire N__16450;
    wire N__16449;
    wire N__16446;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16434;
    wire N__16429;
    wire N__16428;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16407;
    wire N__16406;
    wire N__16403;
    wire N__16398;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16374;
    wire N__16371;
    wire N__16370;
    wire N__16369;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16342;
    wire N__16341;
    wire N__16338;
    wire N__16337;
    wire N__16336;
    wire N__16335;
    wire N__16334;
    wire N__16331;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16317;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16287;
    wire N__16286;
    wire N__16283;
    wire N__16278;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16188;
    wire N__16187;
    wire N__16184;
    wire N__16179;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16056;
    wire N__16055;
    wire N__16054;
    wire N__16053;
    wire N__16046;
    wire N__16045;
    wire N__16044;
    wire N__16043;
    wire N__16040;
    wire N__16039;
    wire N__16038;
    wire N__16037;
    wire N__16036;
    wire N__16035;
    wire N__16034;
    wire N__16031;
    wire N__16030;
    wire N__16029;
    wire N__16028;
    wire N__16027;
    wire N__16026;
    wire N__16025;
    wire N__16024;
    wire N__16023;
    wire N__16020;
    wire N__16009;
    wire N__16004;
    wire N__15999;
    wire N__15992;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15977;
    wire N__15976;
    wire N__15975;
    wire N__15970;
    wire N__15965;
    wire N__15956;
    wire N__15949;
    wire N__15946;
    wire N__15941;
    wire N__15932;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15894;
    wire N__15891;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15886;
    wire N__15885;
    wire N__15884;
    wire N__15883;
    wire N__15882;
    wire N__15881;
    wire N__15878;
    wire N__15873;
    wire N__15870;
    wire N__15859;
    wire N__15856;
    wire N__15845;
    wire N__15838;
    wire N__15829;
    wire N__15826;
    wire N__15823;
    wire N__15820;
    wire N__15817;
    wire N__15814;
    wire N__15811;
    wire N__15810;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15804;
    wire N__15803;
    wire N__15802;
    wire N__15795;
    wire N__15790;
    wire N__15785;
    wire N__15778;
    wire N__15777;
    wire N__15774;
    wire N__15773;
    wire N__15772;
    wire N__15769;
    wire N__15762;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15726;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15711;
    wire N__15710;
    wire N__15709;
    wire N__15702;
    wire N__15699;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15684;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15633;
    wire N__15632;
    wire N__15627;
    wire N__15624;
    wire N__15619;
    wire N__15618;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15600;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15553;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15541;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15523;
    wire N__15520;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15502;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15490;
    wire N__15489;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15456;
    wire N__15453;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15433;
    wire N__15432;
    wire N__15427;
    wire N__15424;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15405;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15390;
    wire N__15389;
    wire N__15386;
    wire N__15383;
    wire N__15380;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15364;
    wire N__15361;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15349;
    wire N__15348;
    wire N__15345;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15325;
    wire N__15322;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15310;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15274;
    wire N__15271;
    wire N__15268;
    wire N__15265;
    wire N__15264;
    wire N__15263;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15238;
    wire N__15237;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15219;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15187;
    wire N__15184;
    wire N__15181;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15139;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15091;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14979;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14959;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14881;
    wire N__14878;
    wire N__14875;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14844;
    wire N__14843;
    wire N__14838;
    wire N__14835;
    wire N__14830;
    wire N__14829;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14814;
    wire N__14813;
    wire N__14810;
    wire N__14805;
    wire N__14802;
    wire N__14797;
    wire N__14796;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14778;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14737;
    wire N__14736;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire VCCG0;
    wire GNDG0;
    wire \b2v_inst16.count_rst_0_cascade_ ;
    wire \b2v_inst16.countZ0Z_11_cascade_ ;
    wire \b2v_inst16.count_4_11 ;
    wire \b2v_inst16.countZ0Z_8_cascade_ ;
    wire \b2v_inst16.count_4_8 ;
    wire \b2v_inst16.count_rst_8_cascade_ ;
    wire \b2v_inst16.countZ0Z_3_cascade_ ;
    wire \b2v_inst16.count_4_3 ;
    wire \b2v_inst16.countZ0Z_9_cascade_ ;
    wire \b2v_inst16.count_rst_14 ;
    wire \b2v_inst16.count_4_9 ;
    wire \b2v_inst16.count_rst_12_cascade_ ;
    wire \b2v_inst16.countZ0Z_7_cascade_ ;
    wire \b2v_inst16.count_4_7 ;
    wire bfn_1_3_0_;
    wire \b2v_inst16.un4_count_1_cry_1 ;
    wire \b2v_inst16.un4_count_1_cry_2_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_2 ;
    wire \b2v_inst16.un4_count_1_cry_3 ;
    wire \b2v_inst16.un4_count_1_cry_4 ;
    wire \b2v_inst16.un4_count_1_cry_5 ;
    wire \b2v_inst16.countZ0Z_7 ;
    wire \b2v_inst16.un4_count_1_cry_6_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_6 ;
    wire \b2v_inst16.un4_count_1_cry_7 ;
    wire \b2v_inst16.un4_count_1_cry_8 ;
    wire \b2v_inst16.countZ0Z_9 ;
    wire \b2v_inst16.un4_count_1_cry_8_THRU_CO ;
    wire bfn_1_4_0_;
    wire \b2v_inst16.un4_count_1_cry_9 ;
    wire \b2v_inst16.un4_count_1_cry_10_THRU_CO ;
    wire \b2v_inst16.un4_count_1_cry_10 ;
    wire \b2v_inst16.un4_count_1_cry_11 ;
    wire \b2v_inst16.un4_count_1_cry_12 ;
    wire \b2v_inst16.un4_count_1_cry_13 ;
    wire \b2v_inst16.un4_count_1_cry_14 ;
    wire \b2v_inst16.delayed_vddq_pwrgd_en ;
    wire \b2v_inst16.delayed_vddq_pwrgdZ0 ;
    wire \b2v_inst16.delayed_vddq_pwrgd_en_cascade_ ;
    wire b2v_inst16_un2_vpp_en_0_i;
    wire \b2v_inst200.count_enZ0 ;
    wire \b2v_inst16.count_rst_7 ;
    wire \b2v_inst16.count_en_cascade_ ;
    wire \b2v_inst16.count_4_2 ;
    wire \b2v_inst11.g3_cascade_ ;
    wire \b2v_inst11.g1_0_1_cascade_ ;
    wire \b2v_inst11.N_7_3_0_cascade_ ;
    wire \b2v_inst11.g2_1_0_0_cascade_ ;
    wire \b2v_inst11.g2_2_0 ;
    wire \b2v_inst11.g2_1_0 ;
    wire \b2v_inst11.g0_12_0 ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ;
    wire \b2v_inst11.N_379_cascade_ ;
    wire SLP_S3n_ibuf_RNIF6NLZ0;
    wire \b2v_inst11.N_379 ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_13 ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2 ;
    wire \b2v_inst11.count_clk_RNIVS8U1Z0Z_14 ;
    wire \b2v_inst11.N_428 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_0 ;
    wire \b2v_inst11.N_175 ;
    wire \b2v_inst11.N_175_cascade_ ;
    wire \b2v_inst11.N_190 ;
    wire \b2v_inst11.N_190_cascade_ ;
    wire \b2v_inst11.un2_count_clk_17_0_o3_0_4 ;
    wire \b2v_inst11.count_clk_en_cascade_ ;
    wire \b2v_inst11.count_clk_0_13 ;
    wire \b2v_inst11.count_clk_0_15 ;
    wire \b2v_inst11.count_clk_0_12 ;
    wire \b2v_inst11.count_clk_0_10 ;
    wire \b2v_inst11.count_clkZ0Z_10_cascade_ ;
    wire \b2v_inst11.un2_count_clk_17_0_o2_4 ;
    wire \b2v_inst11.count_clk_0_11 ;
    wire \b2v_inst11.count_clk_0_4 ;
    wire bfn_1_13_0_;
    wire \b2v_inst20.counter_1_cry_1 ;
    wire \b2v_inst20.counter_1_cry_2 ;
    wire \b2v_inst20.counter_1_cry_3 ;
    wire \b2v_inst20.counter_1_cry_4 ;
    wire \b2v_inst20.counter_1_cry_5 ;
    wire \b2v_inst20.counter_1_cry_6 ;
    wire \b2v_inst20.counter_1_cry_7 ;
    wire \b2v_inst20.counter_1_cry_8 ;
    wire bfn_1_14_0_;
    wire \b2v_inst20.counter_1_cry_9 ;
    wire \b2v_inst20.counter_1_cry_10 ;
    wire \b2v_inst20.counter_1_cry_11 ;
    wire \b2v_inst20.counter_1_cry_12 ;
    wire \b2v_inst20.counter_1_cry_13 ;
    wire \b2v_inst20.counter_1_cry_14 ;
    wire \b2v_inst20.counter_1_cry_15 ;
    wire \b2v_inst20.counter_1_cry_16 ;
    wire bfn_1_15_0_;
    wire \b2v_inst20.counter_1_cry_17 ;
    wire \b2v_inst20.counter_1_cry_18 ;
    wire \b2v_inst20.counter_1_cry_19 ;
    wire \b2v_inst20.counter_1_cry_20 ;
    wire \b2v_inst20.counter_1_cry_21 ;
    wire \b2v_inst20.counter_1_cry_22 ;
    wire \b2v_inst20.counter_1_cry_23 ;
    wire \b2v_inst20.counter_1_cry_24 ;
    wire bfn_1_16_0_;
    wire \b2v_inst20.counter_1_cry_25 ;
    wire \b2v_inst20.counter_1_cry_26 ;
    wire \b2v_inst20.counter_1_cry_27 ;
    wire \b2v_inst20.counter_1_cry_28 ;
    wire \b2v_inst20.counter_1_cry_29 ;
    wire \b2v_inst20.counter_1_cry_30 ;
    wire \b2v_inst16.countZ0Z_0_cascade_ ;
    wire \b2v_inst16.countZ0Z_8 ;
    wire \b2v_inst16.N_416_cascade_ ;
    wire \b2v_inst16.un4_count_1_cry_7_THRU_CO ;
    wire \b2v_inst16.count_rst_13 ;
    wire \b2v_inst16.count_rst_5 ;
    wire \b2v_inst16.un4_count_1_cry_4_THRU_CO ;
    wire \b2v_inst16.count_rst_10_cascade_ ;
    wire \b2v_inst16.count_4_5 ;
    wire \b2v_inst16.countZ0Z_5 ;
    wire \b2v_inst16.count_rst ;
    wire \b2v_inst16.count_4_10 ;
    wire \b2v_inst16.count_rst_11 ;
    wire \b2v_inst16.count_4_6 ;
    wire \b2v_inst16.count_rst_4 ;
    wire \b2v_inst16.count_4_15 ;
    wire \b2v_inst16.count_4_14 ;
    wire \b2v_inst16.count_rst_3 ;
    wire \b2v_inst16.countZ0Z_14 ;
    wire \b2v_inst16.countZ0Z_3 ;
    wire \b2v_inst16.countZ0Z_14_cascade_ ;
    wire \b2v_inst16.countZ0Z_13 ;
    wire \b2v_inst16.count_rst_9_cascade_ ;
    wire \b2v_inst16.countZ0Z_4 ;
    wire \b2v_inst16.un4_count_1_cry_3_THRU_CO ;
    wire \b2v_inst16.countZ0Z_4_cascade_ ;
    wire \b2v_inst16.count_4_4 ;
    wire \b2v_inst16.count_rst_2 ;
    wire \b2v_inst16.count_4_13 ;
    wire \b2v_inst16.un4_count_1_axb_1_cascade_ ;
    wire \b2v_inst16.un4_count_1_axb_1 ;
    wire \b2v_inst16.countZ0Z_6 ;
    wire \b2v_inst16.countZ0Z_12 ;
    wire \b2v_inst16.countZ0Z_10 ;
    wire \b2v_inst16.countZ0Z_2 ;
    wire \b2v_inst16.count_4_1 ;
    wire \b2v_inst16.count_rst_6 ;
    wire \b2v_inst16.countZ0Z_15 ;
    wire \b2v_inst16.countZ0Z_1_cascade_ ;
    wire \b2v_inst16.countZ0Z_11 ;
    wire \b2v_inst16.count_4_i_a3_8_0 ;
    wire \b2v_inst16.count_4_i_a3_10_0 ;
    wire \b2v_inst16.count_4_i_a3_7_0_cascade_ ;
    wire \b2v_inst16.count_4_i_a3_9_0 ;
    wire \b2v_inst16.N_414 ;
    wire \b2v_inst16.countZ0Z_0 ;
    wire \b2v_inst16.N_414_cascade_ ;
    wire \b2v_inst16.count_4_0 ;
    wire \b2v_inst11.count_offZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_off_RNIZ0Z_1 ;
    wire \b2v_inst11.count_off_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_off_0_1 ;
    wire \b2v_inst11.count_off_0_0 ;
    wire \b2v_inst11.count_off_0_10 ;
    wire \b2v_inst16.N_1440 ;
    wire \b2v_inst16.curr_state_RNI3B692Z0Z_0_cascade_ ;
    wire \b2v_inst16.N_416 ;
    wire \b2v_inst16.curr_state_7_0_1_cascade_ ;
    wire \b2v_inst16.curr_state_2_1 ;
    wire \b2v_inst16.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst16.curr_state_2_0 ;
    wire \b2v_inst16.curr_stateZ0Z_1 ;
    wire \b2v_inst16.curr_state_RNI3B692Z0Z_0 ;
    wire \b2v_inst16.N_268 ;
    wire \b2v_inst16.N_268_cascade_ ;
    wire \b2v_inst16.N_26 ;
    wire \b2v_inst11.un1_func_state25_6_0_a3_0_0_cascade_ ;
    wire \b2v_inst11.func_state_RNINPGR_2Z0Z_1_cascade_ ;
    wire \b2v_inst11.g0_20_1 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_ ;
    wire \b2v_inst11.count_clk_RNIVS8U1Z0Z_13 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_329_N ;
    wire \b2v_inst11.un1_func_state25_6_0_1_cascade_ ;
    wire \b2v_inst11.func_state_RNI_1Z0Z_0 ;
    wire N_236_0;
    wire \b2v_inst11.g1_0_0_1 ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_331_N ;
    wire \b2v_inst11.count_clk_en_1 ;
    wire \b2v_inst11.N_328 ;
    wire \b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1 ;
    wire \b2v_inst11.N_340 ;
    wire \b2v_inst11.func_state_1_ss0_i_0_o3_1 ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_1 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz ;
    wire \b2v_inst11.count_off_RNIZ0Z_9_cascade_ ;
    wire \b2v_inst11.func_state_RNI_1Z0Z_1_cascade_ ;
    wire \b2v_inst11.un1_func_state25_4_i_a3_0_1 ;
    wire \b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_clkZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_clk_0_1 ;
    wire \b2v_inst11.count_clk_0_0 ;
    wire \b2v_inst11.count_clk_0_7 ;
    wire \b2v_inst11.N_168_cascade_ ;
    wire \b2v_inst11.func_state_RNICGI84_0_0_cascade_ ;
    wire \b2v_inst11.count_clk_RNI_0Z0Z_0 ;
    wire \b2v_inst11.func_state_RNIVS8U1_0Z0Z_0 ;
    wire \b2v_inst11.count_clk_0_14 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_2 ;
    wire \b2v_inst11.un1_count_clk_1_sqmuxa_0_3 ;
    wire \b2v_inst11.count_clkZ0Z_1 ;
    wire \b2v_inst11.count_clkZ0Z_0 ;
    wire bfn_2_12_0_;
    wire \b2v_inst11.un1_count_clk_2_cry_1 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2 ;
    wire \b2v_inst11.count_clkZ0Z_4 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_3 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5 ;
    wire \b2v_inst11.count_clkZ0Z_7 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_6 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_cZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8 ;
    wire bfn_2_13_0_;
    wire \b2v_inst11.count_clkZ0Z_10 ;
    wire \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_9_cZ0 ;
    wire \b2v_inst11.count_clkZ0Z_11 ;
    wire \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_10_cZ0 ;
    wire \b2v_inst11.count_clkZ0Z_12 ;
    wire \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_11 ;
    wire \b2v_inst11.count_clkZ0Z_13 ;
    wire \b2v_inst11.count_clk_1_13 ;
    wire \b2v_inst11.un1_count_clk_2_cry_12 ;
    wire \b2v_inst11.count_clkZ0Z_14 ;
    wire \b2v_inst11.count_clk_1_14 ;
    wire \b2v_inst11.un1_count_clk_2_cry_13 ;
    wire \b2v_inst11.count_clkZ0Z_15 ;
    wire \b2v_inst11.func_state_RNICGI84_0_0 ;
    wire \b2v_inst11.un1_count_clk_2_cry_14 ;
    wire \b2v_inst11.count_clk_1_15 ;
    wire \b2v_inst20.counterZ0Z_11 ;
    wire \b2v_inst20.counterZ0Z_9 ;
    wire \b2v_inst20.counterZ0Z_10 ;
    wire \b2v_inst20.counterZ0Z_8 ;
    wire \b2v_inst20.counterZ0Z_15 ;
    wire \b2v_inst20.counterZ0Z_14 ;
    wire \b2v_inst20.counterZ0Z_13 ;
    wire \b2v_inst20.counterZ0Z_12 ;
    wire \b2v_inst20.counterZ0Z_19 ;
    wire \b2v_inst20.counterZ0Z_17 ;
    wire \b2v_inst20.counterZ0Z_18 ;
    wire \b2v_inst20.counterZ0Z_16 ;
    wire \b2v_inst20.counterZ0Z_23 ;
    wire \b2v_inst20.counterZ0Z_21 ;
    wire \b2v_inst20.counterZ0Z_22 ;
    wire \b2v_inst20.counterZ0Z_20 ;
    wire VPP_OK_c;
    wire VDDQ_EN_c;
    wire bfn_2_15_0_;
    wire \b2v_inst20.un4_counter_0 ;
    wire \b2v_inst20.un4_counter_2_and ;
    wire \b2v_inst20.un4_counter_1 ;
    wire \b2v_inst20.un4_counter_3_and ;
    wire \b2v_inst20.un4_counter_2 ;
    wire \b2v_inst20.un4_counter_4_and ;
    wire \b2v_inst20.un4_counter_3 ;
    wire \b2v_inst20.un4_counter_5_and ;
    wire \b2v_inst20.un4_counter_4 ;
    wire \b2v_inst20.un4_counter_5 ;
    wire \b2v_inst20.un4_counter_6 ;
    wire b2v_inst20_un4_counter_7;
    wire bfn_2_16_0_;
    wire \b2v_inst20.counterZ0Z_31 ;
    wire \b2v_inst20.counterZ0Z_29 ;
    wire \b2v_inst20.counterZ0Z_30 ;
    wire \b2v_inst20.counterZ0Z_28 ;
    wire \b2v_inst20.un4_counter_7_and ;
    wire \b2v_inst20.counterZ0Z_27 ;
    wire \b2v_inst20.counterZ0Z_25 ;
    wire \b2v_inst20.counterZ0Z_26 ;
    wire \b2v_inst20.counterZ0Z_24 ;
    wire \b2v_inst20.un4_counter_6_and ;
    wire \b2v_inst200.count_3_1 ;
    wire \b2v_inst200.count_3_2 ;
    wire \b2v_inst200.count_3_3 ;
    wire \b2v_inst200.count_3_12 ;
    wire \b2v_inst200.count_3_4 ;
    wire \b2v_inst200.count_3_5 ;
    wire \b2v_inst200.count_3_7 ;
    wire \b2v_inst11.count_off_0_15 ;
    wire \b2v_inst11.count_off_0_13 ;
    wire \b2v_inst11.count_offZ0Z_13_cascade_ ;
    wire \b2v_inst11.count_off_0_8 ;
    wire \b2v_inst11.count_offZ0Z_8_cascade_ ;
    wire \b2v_inst11.count_offZ0Z_0 ;
    wire bfn_4_4_0_;
    wire \b2v_inst11.un3_count_off_1_cry_1 ;
    wire \b2v_inst11.un3_count_off_1_cry_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_3 ;
    wire \b2v_inst11.un3_count_off_1_cry_4 ;
    wire \b2v_inst11.un3_count_off_1_axb_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_5 ;
    wire \b2v_inst11.un3_count_off_1_axb_7 ;
    wire \b2v_inst11.un3_count_off_1_cry_6 ;
    wire \b2v_inst11.count_offZ0Z_8 ;
    wire \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ;
    wire \b2v_inst11.un3_count_off_1_cry_7 ;
    wire \b2v_inst11.un3_count_off_1_cry_8 ;
    wire bfn_4_5_0_;
    wire \b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ;
    wire \b2v_inst11.un3_count_off_1_cry_9 ;
    wire \b2v_inst11.un3_count_off_1_cry_10 ;
    wire \b2v_inst11.un3_count_off_1_cry_11 ;
    wire \b2v_inst11.count_offZ0Z_13 ;
    wire \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ;
    wire \b2v_inst11.un3_count_off_1_cry_12 ;
    wire \b2v_inst11.un3_count_off_1_cry_13 ;
    wire \b2v_inst11.count_offZ0Z_15 ;
    wire \b2v_inst11.un3_count_off_1_cry_14 ;
    wire \b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ;
    wire \b2v_inst11.un3_count_off_1_axb_11 ;
    wire \b2v_inst11.count_off_1_11 ;
    wire \b2v_inst11.count_off_1_11_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ;
    wire \b2v_inst11.count_off_0_12 ;
    wire \b2v_inst11.count_offZ0Z_12 ;
    wire \b2v_inst11.count_offZ0Z_10 ;
    wire \b2v_inst11.un34_clk_100khz_5 ;
    wire \b2v_inst11.un34_clk_100khz_4_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_11 ;
    wire \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ;
    wire \b2v_inst11.count_offZ0Z_11 ;
    wire \b2v_inst11.g4_cascade_ ;
    wire \b2v_inst11.g0_17_N_3L3_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIVGS13Z0Z_7 ;
    wire \b2v_inst11.dutycycleZ1Z_7 ;
    wire \b2v_inst11.dutycycle_RNI24DD8Z0Z_7 ;
    wire \b2v_inst11.dutycycle_RNIVGS13Z0Z_7_cascade_ ;
    wire \b2v_inst11.N_160_i_cascade_ ;
    wire \b2v_inst11.g1_0_sx ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_0_cascade_ ;
    wire \b2v_inst11.func_state_RNI608H1_0Z0Z_1 ;
    wire \b2v_inst11.N_354_cascade_ ;
    wire b2v_inst11_g0_i_m2_i_a6_3_2;
    wire \b2v_inst11.N_159_cascade_ ;
    wire \b2v_inst11.func_state_1_m0_0_1_1_0_cascade_ ;
    wire \b2v_inst11.un1_func_state25_6_0_o_N_313_N ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_sx_cascade_ ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1 ;
    wire \b2v_inst11.func_state_RNI_2Z0Z_1_cascade_ ;
    wire \b2v_inst11.N_337 ;
    wire \b2v_inst11.func_state_1_m2s2_i_0_cascade_ ;
    wire \b2v_inst11.N_338 ;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_6_cascade_ ;
    wire \b2v_inst11.N_231_N ;
    wire \b2v_inst11.N_306_cascade_ ;
    wire \b2v_inst11.func_state_RNI_1Z0Z_1 ;
    wire \b2v_inst11.func_state_1_m2_am_1_1_cascade_ ;
    wire \b2v_inst11.count_off_RNIZ0Z_9 ;
    wire \b2v_inst11.func_state_RNIR5S85Z0Z_1_cascade_ ;
    wire \b2v_inst11.func_state_cascade_ ;
    wire \b2v_inst11.func_stateZ0Z_0 ;
    wire \b2v_inst11.N_160_i ;
    wire \b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ;
    wire \b2v_inst11.func_state_1_m0_0_1_0 ;
    wire \b2v_inst11.func_state_1_m2_1_0_cascade_ ;
    wire \b2v_inst11.N_76 ;
    wire \b2v_inst11.func_state_1_m2_0 ;
    wire func_state_RNIVS8U1_4_1;
    wire \b2v_inst11.func_stateZ0Z_1 ;
    wire \b2v_inst11.count_clk_enZ0Z_0 ;
    wire VCCST_EN_i_0_o3_0_cascade_;
    wire \b2v_inst11.func_state_1_m2_1 ;
    wire func_state_RNI6BE8E_0_1_cascade_;
    wire \b2v_inst11.count_0_7 ;
    wire \b2v_inst11.count_clkZ0Z_3 ;
    wire \b2v_inst11.count_clkZ0Z_6 ;
    wire \b2v_inst11.count_clkZ0Z_8 ;
    wire \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ;
    wire \b2v_inst11.count_clk_0_2 ;
    wire \b2v_inst11.count_clkZ0Z_2 ;
    wire \b2v_inst11.count_clkZ0Z_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ;
    wire \b2v_inst11.count_clk_0_9 ;
    wire \b2v_inst11.count_clkZ0Z_9 ;
    wire \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ;
    wire \b2v_inst11.count_clk_0_3 ;
    wire \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ;
    wire \b2v_inst11.count_clk_0_5 ;
    wire \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ;
    wire \b2v_inst11.count_clk_0_6 ;
    wire \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ;
    wire \b2v_inst11.count_clk_0_8 ;
    wire \b2v_inst11.count_clk_en ;
    wire \b2v_inst20.un4_counter_0_and ;
    wire \b2v_inst11.N_381_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ;
    wire \b2v_inst11.N_381_0 ;
    wire N_15_i_0_a4_0_1;
    wire \b2v_inst20.counter_1_cry_2_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_3 ;
    wire \b2v_inst20.counterZ0Z_0 ;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ;
    wire \b2v_inst20.counter_1_cry_3_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_4 ;
    wire \b2v_inst20.counter_1_cry_4_THRU_CO ;
    wire delayed_vccin_vccinaux_ok_RNI8L1J7_0;
    wire \b2v_inst20.counter_1_cry_1_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_2 ;
    wire bfn_5_1_0_;
    wire \b2v_inst200.countZ0Z_1 ;
    wire \b2v_inst200.count_RNIC03N_5Z0Z_0 ;
    wire \b2v_inst200.un2_count_1_cry_1_cy ;
    wire \b2v_inst200.countZ0Z_2 ;
    wire \b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_1 ;
    wire \b2v_inst200.countZ0Z_3 ;
    wire \b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_2 ;
    wire \b2v_inst200.countZ0Z_4 ;
    wire \b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_3 ;
    wire \b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ;
    wire \b2v_inst200.un2_count_1_cry_4 ;
    wire \b2v_inst200.un2_count_1_cry_5_cZ0 ;
    wire \b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ;
    wire \b2v_inst200.un2_count_1_cry_6 ;
    wire \b2v_inst200.un2_count_1_cry_7 ;
    wire bfn_5_2_0_;
    wire \b2v_inst200.un2_count_1_cry_8 ;
    wire \b2v_inst200.un2_count_1_cry_9 ;
    wire \b2v_inst200.un2_count_1_cry_10 ;
    wire \b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ;
    wire \b2v_inst200.un2_count_1_cry_11 ;
    wire \b2v_inst200.un2_count_1_cry_12 ;
    wire \b2v_inst200.un2_count_1_cry_13 ;
    wire \b2v_inst200.un2_count_1_cry_14 ;
    wire \b2v_inst200.un2_count_1_cry_15 ;
    wire bfn_5_3_0_;
    wire \b2v_inst200.un2_count_1_cry_16 ;
    wire \b2v_inst200.count_0_17 ;
    wire \b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ;
    wire \b2v_inst11.count_off_1_3_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_axb_3 ;
    wire \b2v_inst11.count_offZ0Z_4 ;
    wire \b2v_inst11.count_off_1_3 ;
    wire \b2v_inst11.count_offZ0Z_4_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ;
    wire \b2v_inst11.count_offZ0Z_3 ;
    wire \b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ;
    wire \b2v_inst11.count_off_0_4 ;
    wire \b2v_inst11.count_off_0_14 ;
    wire \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ;
    wire \b2v_inst11.count_offZ0Z_14 ;
    wire \b2v_inst11.count_off_1_2 ;
    wire \b2v_inst11.un3_count_off_1_axb_2 ;
    wire \b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ;
    wire \b2v_inst11.count_offZ0Z_2 ;
    wire \b2v_inst11.count_offZ0Z_5 ;
    wire \b2v_inst11.count_offZ0Z_1 ;
    wire \b2v_inst11.un34_clk_100khz_0 ;
    wire \b2v_inst11.un34_clk_100khz_2 ;
    wire \b2v_inst11.un34_clk_100khz_1_cascade_ ;
    wire \b2v_inst11.un34_clk_100khz_3 ;
    wire \b2v_inst11.un34_clk_100khz_12 ;
    wire \b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ;
    wire \b2v_inst11.count_off_0_5 ;
    wire \b2v_inst11.count_offZ0Z_6 ;
    wire \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ;
    wire \b2v_inst11.count_off_1_9 ;
    wire \b2v_inst11.count_offZ0Z_9 ;
    wire \b2v_inst11.count_off_1_9_cascade_ ;
    wire \b2v_inst11.un3_count_off_1_axb_9 ;
    wire \b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ;
    wire \b2v_inst11.count_off_1_6 ;
    wire \b2v_inst11.count_offZ0Z_7 ;
    wire \b2v_inst11.count_off_enZ0 ;
    wire \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ;
    wire \b2v_inst11.N_125 ;
    wire \b2v_inst11.count_off_1_7 ;
    wire \b2v_inst11.g0_3_0 ;
    wire \b2v_inst11.g2_0 ;
    wire \b2v_inst11.dutycycle_eena_8_cascade_ ;
    wire \b2v_inst11.dutycycle_rst_7 ;
    wire \b2v_inst11.dutycycle_0_3 ;
    wire \b2v_inst11.dutycycle_rst_7_cascade_ ;
    wire \b2v_inst11.dutycycle_eena_8 ;
    wire \b2v_inst11.dutycycleZ0Z_3_cascade_ ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_0_d_0 ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_0_ccf1 ;
    wire \b2v_inst11.un1_clk_100khz_43_and_i_0_c ;
    wire \b2v_inst11.N_307_cascade_ ;
    wire \b2v_inst11.N_234_N ;
    wire \b2v_inst11.N_308 ;
    wire \b2v_inst11.N_234_N_cascade_ ;
    wire \b2v_inst11.func_state_RNI9R6T4Z0Z_1_cascade_ ;
    wire \b2v_inst11.func_state_RNI9R6T4Z0Z_1 ;
    wire \b2v_inst11.dutycycleZ1Z_11 ;
    wire \b2v_inst11.N_159 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ;
    wire \b2v_inst11.N_155_N_cascade_ ;
    wire \b2v_inst11.dutycycle_en_11_cascade_ ;
    wire \b2v_inst11.N_305 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_6 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_6_cascade_ ;
    wire \b2v_inst11.i2_mux_cascade_ ;
    wire \b2v_inst11.N_301 ;
    wire \b2v_inst11.N_382_cascade_ ;
    wire \b2v_inst11.g0_2_0_cascade_ ;
    wire \b2v_inst11.N_430 ;
    wire \b2v_inst11.func_state_RNIRF2E4Z0Z_0 ;
    wire VCCST_EN_i_0_i;
    wire \b2v_inst11.un1_clk_100khz_2_i_o3_sx ;
    wire \b2v_inst11.func_state ;
    wire \b2v_inst11.func_state_RNI_0Z0Z_0 ;
    wire \b2v_inst5.N_2897_i_cascade_ ;
    wire \b2v_inst5.curr_state_0_0 ;
    wire \b2v_inst5.m4_0_cascade_ ;
    wire \b2v_inst11.g2_0_1_cascade_ ;
    wire dutycycle_RNISSAOS1_0_5_cascade_;
    wire \b2v_inst11.dutycycle_RNIZ0Z_5_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_1 ;
    wire \b2v_inst11.N_73_mux_i_i_o7_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIUNGA5Z0Z_5 ;
    wire \b2v_inst11.N_73_mux_i_i_0 ;
    wire \b2v_inst11.N_73_mux_i_i_a7_1_cascade_ ;
    wire g0_0_0;
    wire N_5_0;
    wire b2v_inst11_un1_dutycycle_172_m3_amcf1;
    wire N_73_mux_i_i_a7_4_0_1_cascade_;
    wire N_73_mux_i_i_a7_4_0_cascade_;
    wire \b2v_inst11.N_73_mux_i_i_1 ;
    wire \b2v_inst11.N_73_mux_i_i_2 ;
    wire N_15;
    wire \b2v_inst11.N_73_mux_i_i_1_cascade_ ;
    wire \b2v_inst11.dutycycle_0_5 ;
    wire \b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx ;
    wire RSMRSTn_fast_RNIGMH81_cascade_;
    wire N_7_2;
    wire N_10_0;
    wire \b2v_inst20.tmp_1_rep1_RNI07FZ0Z73 ;
    wire \b2v_inst20.counter_1_cry_5_THRU_CO ;
    wire \b2v_inst20.counterZ0Z_7 ;
    wire \b2v_inst20.counterZ0Z_5 ;
    wire \b2v_inst20.counterZ0Z_6 ;
    wire \b2v_inst20.counterZ0Z_1 ;
    wire \b2v_inst20.un4_counter_1_and ;
    wire SYNTHESIZED_WIRE_1keep_3_fast;
    wire HDA_SDO_ATP_c;
    wire \b2v_inst200.N_205 ;
    wire \b2v_inst200.N_205_cascade_ ;
    wire G_2734_cascade_;
    wire \b2v_inst200.curr_stateZ0Z_2 ;
    wire \b2v_inst200.curr_stateZ0Z_2_cascade_ ;
    wire \b2v_inst200.HDA_SDO_ATP_0 ;
    wire G_2734;
    wire \b2v_inst200.curr_state_0_2 ;
    wire \b2v_inst200.countZ0Z_6 ;
    wire \b2v_inst200.countZ0Z_6_cascade_ ;
    wire \b2v_inst200.countZ0Z_8 ;
    wire \b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ;
    wire \b2v_inst200.count_3_6 ;
    wire \b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0 ;
    wire \b2v_inst200.count_3_8 ;
    wire \b2v_inst200.count_1_0 ;
    wire \b2v_inst200.countZ0Z_0_cascade_ ;
    wire \b2v_inst200.count_3_0 ;
    wire \b2v_inst200.countZ0Z_12 ;
    wire \b2v_inst200.count_3_13 ;
    wire \b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ;
    wire \b2v_inst200.countZ0Z_13 ;
    wire \b2v_inst200.countZ0Z_13_cascade_ ;
    wire \b2v_inst200.countZ0Z_0 ;
    wire \b2v_inst200.countZ0Z_7 ;
    wire \b2v_inst200.countZ0Z_5 ;
    wire \b2v_inst200.un25_clk_100khz_10_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_3 ;
    wire \b2v_inst200.countZ0Z_15 ;
    wire \b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ;
    wire \b2v_inst200.count_3_15 ;
    wire \b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ;
    wire \b2v_inst200.count_3_14 ;
    wire \b2v_inst200.countZ0Z_14 ;
    wire \b2v_inst200.count_0_16 ;
    wire \b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79 ;
    wire \b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29 ;
    wire \b2v_inst200.count_3_11 ;
    wire \b2v_inst200.countZ0Z_11 ;
    wire \b2v_inst200.countZ0Z_17 ;
    wire \b2v_inst200.countZ0Z_11_cascade_ ;
    wire \b2v_inst200.countZ0Z_16 ;
    wire \b2v_inst200.un25_clk_100khz_9 ;
    wire \b2v_inst200.un25_clk_100khz_12 ;
    wire \b2v_inst200.un25_clk_100khz_13_cascade_ ;
    wire \b2v_inst200.un25_clk_100khz_14 ;
    wire \b2v_inst200.count_RNIC03N_6Z0Z_0_cascade_ ;
    wire \b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0 ;
    wire \b2v_inst200.count_3_10 ;
    wire \b2v_inst200.count_RNI_0_0_cascade_ ;
    wire \b2v_inst200.countZ0Z_10 ;
    wire \b2v_inst16.count_rst_1 ;
    wire \b2v_inst16.count_4_12 ;
    wire \b2v_inst16.count_en ;
    wire \b2v_inst16.N_2987_i ;
    wire \b2v_inst11.N_366 ;
    wire bfn_6_6_0_;
    wire \b2v_inst11.mult1_un152_sum_cry_2_c ;
    wire \b2v_inst11.mult1_un152_sum_cry_3_c ;
    wire \b2v_inst11.mult1_un152_sum_cry_4_c ;
    wire \b2v_inst11.mult1_un152_sum_cry_5_c ;
    wire \b2v_inst11.mult1_un152_sum_cry_6_c ;
    wire \b2v_inst11.mult1_un152_sum_cry_7 ;
    wire \b2v_inst11.mult1_un145_sum_i_0_8 ;
    wire VDDQ_OK_c;
    wire VCCST_EN_i_0_o3_0;
    wire \b2v_inst16.N_208_0 ;
    wire \b2v_inst11.N_354 ;
    wire \b2v_inst11.un2_count_clk_17_0_a2_1_3 ;
    wire \b2v_inst11.un2_count_clk_17_0_a2_1_2_cascade_ ;
    wire \b2v_inst11.N_363 ;
    wire \b2v_inst11.N_360 ;
    wire \b2v_inst11.N_363_cascade_ ;
    wire \b2v_inst11.N_365 ;
    wire \b2v_inst11.N_365_cascade_ ;
    wire \b2v_inst11.N_293 ;
    wire \b2v_inst11.un1_dutycycle_53_30_1_0_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_9 ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_11 ;
    wire \b2v_inst11.dutycycle_RNI_7Z0Z_1 ;
    wire bfn_6_9_0_;
    wire \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_2 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_4_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_cZ0 ;
    wire bfn_6_10_0_;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_10_cZ0 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ;
    wire \b2v_inst11.dutycycle_RNIP7P13Z0Z_4 ;
    wire \b2v_inst11.dutycycleZ1Z_4 ;
    wire \b2v_inst11.dutycycle_RNIP7P13Z0Z_4_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_7_cascade_ ;
    wire \b2v_inst11.dutycycle_e_1_4 ;
    wire \b2v_inst11.N_158_N_cascade_ ;
    wire \b2v_inst11.dutycycle_0_6 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQZ0Z6 ;
    wire \b2v_inst11.dutycycle_e_1_6 ;
    wire \b2v_inst11.func_state_RNI_5Z0Z_1 ;
    wire \b2v_inst11.N_186_cascade_ ;
    wire \b2v_inst11.N_426_0 ;
    wire b2v_inst11_g0_i_m2_i_a6_1_1_cascade_;
    wire SLP_S3n_ibuf_RNI9HQHZ0Z3;
    wire \b2v_inst11.dutycycle_RNI_9Z0Z_1 ;
    wire \b2v_inst11.N_165_0 ;
    wire \b2v_inst11.g0_i_m2_i_0_1_cascade_ ;
    wire N_15_i_0_a4_1_0;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_0 ;
    wire \b2v_inst11.N_19_i ;
    wire \b2v_inst11.N_5572_0 ;
    wire \b2v_inst11.N_172 ;
    wire \b2v_inst11.un1_count_off_1_sqmuxa_8_m2_1 ;
    wire \b2v_inst11.dutycycle_eena ;
    wire \b2v_inst11.dutycycleZ1Z_0 ;
    wire \b2v_inst11.dutycycle_1_0_0 ;
    wire \b2v_inst11.dutycycle_eena_cascade_ ;
    wire \b2v_inst11.N_117_f0_1 ;
    wire \b2v_inst11.dutycycle_eena_0_cascade_ ;
    wire \b2v_inst11.dutycycle_cascade_ ;
    wire \b2v_inst11.dutycycle_1_0_1 ;
    wire \b2v_inst11.dutycycle_eena_0 ;
    wire \b2v_inst11.dutycycleZ1Z_1 ;
    wire \b2v_inst5.curr_state_RNIZ0Z_1_cascade_ ;
    wire b2v_inst5_RSMRSTn_latmux;
    wire b2v_inst5_RSMRSTn_fast;
    wire RSMRSTn_0;
    wire \b2v_inst5.N_2897_i ;
    wire \b2v_inst5.curr_stateZ0Z_0 ;
    wire \b2v_inst5.curr_state_RNIZ0Z_1 ;
    wire \b2v_inst5.N_51_cascade_ ;
    wire \b2v_inst11.count_0_9 ;
    wire \b2v_inst11.count_0_10 ;
    wire \b2v_inst11.count_0_11 ;
    wire \b2v_inst11.count_0_2 ;
    wire \b2v_inst200.N_56_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst200.count_RNI_0_0 ;
    wire GPIO_FPGA_SoC_1_c;
    wire N_411_cascade_;
    wire \b2v_inst200.m6_i_0 ;
    wire \b2v_inst200.m6_i_0_cascade_ ;
    wire \b2v_inst200.curr_state_3_0 ;
    wire \b2v_inst200.N_58_cascade_ ;
    wire \b2v_inst200.curr_stateZ0Z_0 ;
    wire \b2v_inst200.curr_stateZ0Z_0_cascade_ ;
    wire N_412;
    wire N_412_cascade_;
    wire \b2v_inst200.curr_stateZ0Z_1 ;
    wire \b2v_inst200.curr_state_3_1 ;
    wire \b2v_inst36.count_2_6 ;
    wire \b2v_inst36.count_2_4 ;
    wire \b2v_inst36.count_2_9 ;
    wire \b2v_inst36.count_2_12 ;
    wire \b2v_inst36.curr_state_RNI8TT2Z0Z_0_cascade_ ;
    wire DSW_PWROK_c;
    wire \b2v_inst36.DSW_PWROK_0 ;
    wire \b2v_inst36.curr_state_0_0 ;
    wire \b2v_inst36.curr_state_7_0_cascade_ ;
    wire \b2v_inst36.curr_stateZ0Z_0 ;
    wire \b2v_inst36.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst36.N_2939_i_cascade_ ;
    wire bfn_7_5_0_;
    wire \b2v_inst11.mult1_un131_sum_cry_2 ;
    wire \b2v_inst11.mult1_un131_sum_cry_3 ;
    wire \b2v_inst11.mult1_un131_sum_cry_4 ;
    wire \b2v_inst11.mult1_un131_sum_cry_5 ;
    wire \b2v_inst11.mult1_un131_sum_cry_6 ;
    wire \b2v_inst11.mult1_un131_sum_cry_7 ;
    wire \b2v_inst11.mult1_un131_sum_axb_7_l_fx ;
    wire bfn_7_6_0_;
    wire \b2v_inst11.mult1_un124_sum_cry_2 ;
    wire \b2v_inst11.mult1_un124_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_3 ;
    wire \b2v_inst11.mult1_un124_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_4 ;
    wire \b2v_inst11.mult1_un124_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un124_sum_cry_5 ;
    wire \b2v_inst11.mult1_un131_sum_axb_8 ;
    wire \b2v_inst11.mult1_un124_sum_cry_6 ;
    wire \b2v_inst11.mult1_un124_sum_cry_7 ;
    wire \b2v_inst11.mult1_un124_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un124_sum_i_0_8 ;
    wire \b2v_inst11.N_382 ;
    wire \b2v_inst11.N_302 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_9 ;
    wire \b2v_inst11.mult1_un124_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un131_sum_axb_4_l_fx ;
    wire \b2v_inst11.g0_13_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_9_cascade_ ;
    wire \b2v_inst200.count_RNIC03N_6Z0Z_0 ;
    wire N_411;
    wire \b2v_inst200.m11_0_a3_0 ;
    wire \b2v_inst5.count_rst_10_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_4_cascade_ ;
    wire \b2v_inst5.count_1_8 ;
    wire \b2v_inst5.count_rst_10 ;
    wire \b2v_inst5.countZ0Z_8_cascade_ ;
    wire \b2v_inst5.count_1_4 ;
    wire \b2v_inst5.un12_clk_100khz_7_cascade_ ;
    wire \b2v_inst11.N_8_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_ ;
    wire \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ;
    wire \b2v_inst11.dutycycle_en_11 ;
    wire \b2v_inst11.dutycycleZ0Z_14 ;
    wire \b2v_inst11.dutycycleZ0Z_12_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_11 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_3 ;
    wire \b2v_inst11.dutycycleZ0Z_8_cascade_ ;
    wire \b2v_inst11.N_153_N_cascade_ ;
    wire \b2v_inst11.N_156_N_cascade_ ;
    wire \b2v_inst11.dutycycle_e_1_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ;
    wire \b2v_inst11.dutycycle_e_1_9_cascade_ ;
    wire \b2v_inst11.dutycycleZ1Z_9 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ;
    wire \b2v_inst11.dutycycle_en_10 ;
    wire \b2v_inst11.dutycycleZ0Z_13 ;
    wire \b2v_inst11.dutycycleZ0Z_5_cascade_ ;
    wire \b2v_inst11.N_326_N ;
    wire \b2v_inst11.N_140_N ;
    wire \b2v_inst11.N_425 ;
    wire \b2v_inst11.N_154_N_cascade_ ;
    wire \b2v_inst11.dutycycle_en_4_cascade_ ;
    wire \b2v_inst11.dutycycle_e_1_8 ;
    wire \b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ;
    wire \b2v_inst11.dutycycle_en_4 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69 ;
    wire \b2v_inst11.dutycycleZ0Z_10 ;
    wire \b2v_inst11.dutycycleZ1Z_8 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49 ;
    wire \b2v_inst11.dutycycle_RNI1KT13Z0Z_8 ;
    wire GPIO_FPGA_SoC_4_c;
    wire N_161;
    wire \b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ;
    wire SLP_S3n_c;
    wire \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIZ0 ;
    wire \b2v_inst11.func_state_RNI_2Z0Z_1 ;
    wire SLP_S4n_c;
    wire \b2v_inst11.g1_0_0_cascade_ ;
    wire \b2v_inst11.N_295 ;
    wire \b2v_inst11.g1 ;
    wire \b2v_inst11.g1_cascade_ ;
    wire \b2v_inst11.g1_0 ;
    wire \b2v_inst11.dutycycleZ0Z_2 ;
    wire RSMRSTn_fast_RNIGMH81;
    wire func_state_RNI6BE8E_0_1;
    wire b2v_inst11_dutycycle_1_0_iv_0_o3_out;
    wire func_state_RNI_4_0;
    wire bfn_7_13_0_;
    wire \b2v_inst11.count_1_2 ;
    wire \b2v_inst11.un1_count_cry_1 ;
    wire \b2v_inst11.un1_count_cry_2 ;
    wire \b2v_inst11.un1_count_cry_3 ;
    wire \b2v_inst11.un1_count_cry_4 ;
    wire \b2v_inst11.un1_count_cry_5 ;
    wire \b2v_inst11.count_1_7 ;
    wire \b2v_inst11.un1_count_cry_6 ;
    wire \b2v_inst11.un1_count_cry_7 ;
    wire \b2v_inst11.un1_count_cry_8 ;
    wire \b2v_inst11.count_1_9 ;
    wire bfn_7_14_0_;
    wire \b2v_inst11.count_1_10 ;
    wire \b2v_inst11.un1_count_cry_9 ;
    wire \b2v_inst11.count_1_11 ;
    wire \b2v_inst11.un1_count_cry_10 ;
    wire \b2v_inst11.un1_count_cry_11 ;
    wire \b2v_inst11.un1_count_cry_12 ;
    wire \b2v_inst11.un1_count_cry_13 ;
    wire \b2v_inst11.un1_count_cry_14 ;
    wire \b2v_inst11.count_1_5 ;
    wire \b2v_inst11.count_0_5 ;
    wire \b2v_inst11.count_1_14 ;
    wire \b2v_inst11.count_0_14 ;
    wire \b2v_inst11.count_1_6 ;
    wire \b2v_inst11.count_0_6 ;
    wire \b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ;
    wire \b2v_inst11.count_0_15 ;
    wire \b2v_inst11.pwm_out_en_cascade_ ;
    wire PWRBTN_LED_c;
    wire \b2v_inst11.pwm_out_1_sqmuxa_0 ;
    wire SYNTHESIZED_WIRE_1keep_3_rep1;
    wire b2v_inst20_un4_counter_7_THRU_CO;
    wire \b2v_inst36.countZ0Z_1_cascade_ ;
    wire \b2v_inst36.un12_clk_100khz_9 ;
    wire \b2v_inst36.un12_clk_100khz_10_cascade_ ;
    wire \b2v_inst36.count_2_0 ;
    wire \b2v_inst36.countZ0Z_0_cascade_ ;
    wire \b2v_inst36.count_rst_13 ;
    wire \b2v_inst36.count_rst_13_cascade_ ;
    wire \b2v_inst36.un2_count_1_axb_1_cascade_ ;
    wire \b2v_inst36.count_2_1 ;
    wire \b2v_inst36.un12_clk_100khz_8 ;
    wire \b2v_inst36.count_rst_14 ;
    wire \b2v_inst36.count_rst_3_cascade_ ;
    wire \b2v_inst36.countZ0Z_11_cascade_ ;
    wire \b2v_inst36.count_2_11 ;
    wire \b2v_inst36.count_rst_12_cascade_ ;
    wire \b2v_inst36.countZ0Z_2_cascade_ ;
    wire \b2v_inst36.count_2_2 ;
    wire \b2v_inst36.curr_state_7_1 ;
    wire \b2v_inst36.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst36.curr_state_0_1 ;
    wire \b2v_inst36.N_2939_i ;
    wire V33DSW_OK_c;
    wire \b2v_inst36.curr_stateZ0Z_1 ;
    wire \b2v_inst36.count_rst_7_cascade_ ;
    wire \b2v_inst36.N_2942_i_cascade_ ;
    wire \b2v_inst200.countZ0Z_9 ;
    wire \b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ;
    wire \b2v_inst200.count_3_9 ;
    wire \b2v_inst200.count_en_g ;
    wire \b2v_inst36.count_2_14 ;
    wire \b2v_inst5.count_1_11 ;
    wire \b2v_inst5.count_1_12 ;
    wire \b2v_inst5.count_1_14 ;
    wire bfn_8_5_0_;
    wire \b2v_inst11.mult1_un138_sum_cry_2 ;
    wire \b2v_inst11.mult1_un131_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_3 ;
    wire \b2v_inst11.mult1_un131_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_4 ;
    wire \b2v_inst11.mult1_un131_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_5 ;
    wire \b2v_inst11.mult1_un131_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un138_sum_cry_6 ;
    wire \b2v_inst11.mult1_un138_sum_axb_8 ;
    wire \b2v_inst11.mult1_un138_sum_cry_7 ;
    wire \b2v_inst11.mult1_un131_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un117_sum_i ;
    wire \b2v_inst11.mult1_un131_sum_i ;
    wire \b2v_inst11.mult1_un131_sum_s_8 ;
    wire \b2v_inst11.mult1_un124_sum_i ;
    wire \b2v_inst11.mult1_un145_sum_i ;
    wire bfn_8_7_0_;
    wire \b2v_inst11.mult1_un117_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_2 ;
    wire \b2v_inst11.mult1_un117_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_3 ;
    wire \b2v_inst11.mult1_un117_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_4 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un117_sum_cry_5 ;
    wire \b2v_inst11.mult1_un124_sum_axb_8 ;
    wire \b2v_inst11.mult1_un117_sum_cry_6 ;
    wire \b2v_inst11.mult1_un117_sum_cry_7 ;
    wire \b2v_inst11.mult1_un117_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un117_sum_i_0_8 ;
    wire \b2v_inst5.curr_stateZ0Z_1 ;
    wire N_413;
    wire \b2v_inst11.mult1_un110_sum_i ;
    wire \b2v_inst5.un12_clk_100khz_13 ;
    wire \b2v_inst11.un1_dutycycle_53_axb_11 ;
    wire \b2v_inst11.i7_mux_cascade_ ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_11_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_3Z0Z_9 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_8_cascade_ ;
    wire \b2v_inst11.N_15_mux ;
    wire \b2v_inst11.i6_mux_i_1 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_11 ;
    wire \b2v_inst11.dutycycle_RNI9R6T4Z0Z_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5 ;
    wire \b2v_inst11.dutycycleZ1Z_12 ;
    wire \b2v_inst11.N_224_iZ0 ;
    wire \b2v_inst11.dutycycleZ0Z_15 ;
    wire func_state_RNIVS8U1_3_1;
    wire \b2v_inst11.dutycycle_en_12 ;
    wire \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ;
    wire \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_3_1 ;
    wire \b2v_inst11.un1_dutycycle_53_50_1_i_i_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_1 ;
    wire \b2v_inst11.un1_dutycycle_53_50_1_i_0_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_1_cascade_ ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_3_cascade_ ;
    wire \b2v_inst11.dutycycleZ0Z_5 ;
    wire \b2v_inst11.m6_0_1 ;
    wire \b2v_inst11.dutycycleZ1Z_6 ;
    wire \b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_0_1 ;
    wire N_18;
    wire \b2v_inst11.g2_0_0 ;
    wire b2v_inst11_un1_dutycycle_164_0;
    wire \b2v_inst5.N_6 ;
    wire b2v_inst11_un1_dutycycle_164_0_cascade_;
    wire \b2v_inst5.N_13 ;
    wire \b2v_inst11.N_3060_i ;
    wire \b2v_inst11.un1_dutycycle_96_0_a3_1 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_7 ;
    wire \b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_5 ;
    wire N_73_mux_i_i_o3_1_1;
    wire \b2v_inst11.dutycycleZ1Z_3 ;
    wire \b2v_inst11.g3_0_1 ;
    wire \b2v_inst11.N_3038_i ;
    wire g3_0_4;
    wire \b2v_inst11.count_1_12 ;
    wire \b2v_inst11.count_0_12 ;
    wire \b2v_inst11.count_1_3 ;
    wire \b2v_inst11.count_0_3 ;
    wire \b2v_inst11.count_1_13 ;
    wire \b2v_inst11.count_0_13 ;
    wire \b2v_inst11.count_1_4 ;
    wire \b2v_inst11.count_0_4 ;
    wire \b2v_inst11.un79_clk_100khzlto15_5_cascade_ ;
    wire \b2v_inst11.un79_clk_100khzlt6 ;
    wire \b2v_inst11.un79_clk_100khzlto15_4_cascade_ ;
    wire \b2v_inst11.un79_clk_100khzlto15_7 ;
    wire \b2v_inst11.count_RNIZ0Z_13_cascade_ ;
    wire \b2v_inst11.countZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_1_1_cascade_ ;
    wire \b2v_inst11.countZ0Z_1_cascade_ ;
    wire \b2v_inst11.count_0_1 ;
    wire \b2v_inst11.count_0_0 ;
    wire b2v_inst11_dutycycle_set_1;
    wire G_146;
    wire N_15_i_0_a4_1;
    wire N_73_mux_i_i_a7_0_0;
    wire \b2v_inst11.count_1_8 ;
    wire \b2v_inst11.count_0_8 ;
    wire \b2v_inst11.g0_2_1 ;
    wire \b2v_inst11.pwm_outZ0 ;
    wire \b2v_inst11.pwm_out_1_sqmuxa ;
    wire \b2v_inst11.curr_state_3_0_cascade_ ;
    wire \b2v_inst11.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst11.count_0_sqmuxa_i ;
    wire \b2v_inst11.count_0_sqmuxa_i_cascade_ ;
    wire \b2v_inst11.count_1_0 ;
    wire \b2v_inst36.un2_count_1_axb_1 ;
    wire \b2v_inst36.countZ0Z_0 ;
    wire bfn_9_1_0_;
    wire \b2v_inst36.un2_count_1_cry_1_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_1 ;
    wire \b2v_inst36.un2_count_1_cry_2 ;
    wire \b2v_inst36.countZ0Z_4 ;
    wire \b2v_inst36.count_rst_10 ;
    wire \b2v_inst36.un2_count_1_cry_3 ;
    wire \b2v_inst36.un2_count_1_cry_4 ;
    wire \b2v_inst36.countZ0Z_6 ;
    wire \b2v_inst36.count_rst_8 ;
    wire \b2v_inst36.un2_count_1_cry_5 ;
    wire \b2v_inst36.un2_count_1_cry_6 ;
    wire \b2v_inst36.un2_count_1_cry_7 ;
    wire \b2v_inst36.un2_count_1_cry_8 ;
    wire \b2v_inst36.countZ0Z_9 ;
    wire \b2v_inst36.count_rst_5 ;
    wire bfn_9_2_0_;
    wire \b2v_inst36.un2_count_1_cry_9 ;
    wire \b2v_inst36.countZ0Z_11 ;
    wire \b2v_inst36.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst36.un2_count_1_cry_10 ;
    wire \b2v_inst36.countZ0Z_12 ;
    wire \b2v_inst36.count_rst_2 ;
    wire \b2v_inst36.un2_count_1_cry_11 ;
    wire \b2v_inst36.un2_count_1_cry_12 ;
    wire \b2v_inst36.countZ0Z_14 ;
    wire \b2v_inst36.count_rst_0 ;
    wire \b2v_inst36.un2_count_1_cry_13 ;
    wire \b2v_inst36.un2_count_1_cry_14 ;
    wire \b2v_inst36.count_rst_6 ;
    wire \b2v_inst36.countZ0Z_8 ;
    wire \b2v_inst36.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst36.countZ0Z_8_cascade_ ;
    wire \b2v_inst36.count_2_8 ;
    wire \b2v_inst36.count_rst_4_cascade_ ;
    wire \b2v_inst36.countZ0Z_10 ;
    wire \b2v_inst36.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst36.countZ0Z_10_cascade_ ;
    wire \b2v_inst36.count_2_10 ;
    wire \b2v_inst36.countZ0Z_13 ;
    wire \b2v_inst36.count_rst_1 ;
    wire \b2v_inst36.count_2_13 ;
    wire \b2v_inst36.count_2_15 ;
    wire \b2v_inst36.count_rst ;
    wire \b2v_inst36.countZ0Z_15 ;
    wire \b2v_inst5.un12_clk_100khz_4 ;
    wire \b2v_inst5.count_1_2 ;
    wire \b2v_inst5.count_RNIZ0Z_1_cascade_ ;
    wire \b2v_inst5.count_1_3 ;
    wire \b2v_inst5.count_RNIZ0Z_1 ;
    wire \b2v_inst5.count_1_1 ;
    wire \b2v_inst5.count_rst_14_cascade_ ;
    wire \b2v_inst5.count_rst_1_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_13_cascade_ ;
    wire \b2v_inst5.count_rst_1 ;
    wire \b2v_inst5.count_1_13 ;
    wire \b2v_inst5.un12_clk_100khz_5 ;
    wire \b2v_inst5.count_rst_6 ;
    wire \b2v_inst5.un12_clk_100khz_8 ;
    wire bfn_9_6_0_;
    wire \b2v_inst11.mult1_un138_sum_i ;
    wire \b2v_inst11.mult1_un145_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_2 ;
    wire \b2v_inst11.mult1_un138_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_3 ;
    wire \b2v_inst11.mult1_un138_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_4 ;
    wire \b2v_inst11.mult1_un138_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un145_sum_cry_5 ;
    wire \b2v_inst11.mult1_un138_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un152_sum_axb_8 ;
    wire \b2v_inst11.mult1_un145_sum_cry_6 ;
    wire \b2v_inst11.mult1_un145_sum_axb_8 ;
    wire \b2v_inst11.mult1_un145_sum_cry_7 ;
    wire \b2v_inst11.mult1_un138_sum_i_0_8 ;
    wire bfn_9_7_0_;
    wire \b2v_inst11.mult1_un103_sum_i ;
    wire \b2v_inst11.mult1_un110_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_2 ;
    wire \b2v_inst11.mult1_un110_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_3 ;
    wire \b2v_inst11.mult1_un110_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_4 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un110_sum_cry_5 ;
    wire \b2v_inst11.mult1_un117_sum_axb_8 ;
    wire \b2v_inst11.mult1_un110_sum_cry_6 ;
    wire \b2v_inst11.mult1_un110_sum_cry_7 ;
    wire \b2v_inst11.mult1_un110_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un110_sum_i_0_8 ;
    wire bfn_9_8_0_;
    wire \b2v_inst11.mult1_un103_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_2 ;
    wire \b2v_inst11.mult1_un103_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_3 ;
    wire \b2v_inst11.mult1_un103_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_4 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un103_sum_cry_5 ;
    wire \b2v_inst11.mult1_un96_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un110_sum_axb_8 ;
    wire \b2v_inst11.mult1_un103_sum_cry_6 ;
    wire \b2v_inst11.mult1_un103_sum_cry_7 ;
    wire \b2v_inst11.mult1_un103_sum_s_8 ;
    wire \b2v_inst11.mult1_un103_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un103_sum_i_0_8 ;
    wire \b2v_inst11.dutycycleZ0Z_3 ;
    wire \b2v_inst11.un1_dutycycle_53_axb_0 ;
    wire bfn_9_9_0_;
    wire \b2v_inst11.dutycycle_RNI_5Z0Z_1 ;
    wire \b2v_inst11.mult1_un138_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_0 ;
    wire \b2v_inst11.mult1_un131_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_1 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_2 ;
    wire \b2v_inst11.mult1_un124_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_2 ;
    wire \b2v_inst11.dutycycle_RNI_4Z0Z_3 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_3 ;
    wire \b2v_inst11.mult1_un117_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_3 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_8 ;
    wire \b2v_inst11.mult1_un110_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_4 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_9 ;
    wire \b2v_inst11.mult1_un103_sum ;
    wire \b2v_inst11.un1_dutycycle_53_cry_5 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_9 ;
    wire \b2v_inst11.dutycycleZ0Z_4 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_6 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_7 ;
    wire \b2v_inst11.dutycycleZ0Z_6 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_11 ;
    wire bfn_9_10_0_;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_12 ;
    wire \b2v_inst11.dutycycleZ0Z_9 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_8 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_9 ;
    wire \b2v_inst11.dutycycle_RNI_0Z0Z_14 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_10 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_11 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_11 ;
    wire \b2v_inst11.dutycycleZ0Z_8 ;
    wire \b2v_inst11.dutycycle_RNI_2Z0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_12 ;
    wire \b2v_inst11.dutycycleZ0Z_12 ;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_13 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_13 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_15 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14 ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15 ;
    wire \b2v_inst11.dutycycle_RNIZ0Z_14 ;
    wire \b2v_inst11.dutycycleZ0Z_11 ;
    wire bfn_9_11_0_;
    wire \b2v_inst11.CO2 ;
    wire \b2v_inst11.dutycycleZ0Z_7 ;
    wire dutycycle_RNISSAOS1_0_5;
    wire \b2v_inst11.dutycycle_RNI_1Z0Z_1 ;
    wire \b2v_inst11.curr_stateZ0Z_0 ;
    wire \b2v_inst11.count_RNIZ0Z_13 ;
    wire \b2v_inst11.curr_state_4_0 ;
    wire \b2v_inst11.CO2_THRU_CO ;
    wire \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ;
    wire bfn_9_13_0_;
    wire \b2v_inst11.mult1_un47_sum_i ;
    wire \b2v_inst11.mult1_un54_sum_cry_2 ;
    wire \b2v_inst11.mult1_un54_sum_cry_3 ;
    wire \b2v_inst11.mult1_un54_sum_cry_4 ;
    wire \b2v_inst11.mult1_un54_sum_cry_5 ;
    wire \b2v_inst11.mult1_un47_sum_s_6 ;
    wire \b2v_inst11.mult1_un47_sum_l_fx_6 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6 ;
    wire \b2v_inst11.mult1_un40_sum_i_5 ;
    wire \b2v_inst11.mult1_un54_sum_cry_7 ;
    wire \b2v_inst11.mult1_un47_sum_l_fx_3 ;
    wire \b2v_inst11.mult1_un47_sum ;
    wire bfn_9_14_0_;
    wire \b2v_inst11.mult1_un47_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un47_sum_cry_2 ;
    wire \b2v_inst11.mult1_un47_sum_s_4_sf ;
    wire \b2v_inst11.mult1_un47_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un47_sum_cry_3 ;
    wire \b2v_inst11.mult1_un40_sum_i_l_ofx_4 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un47_sum_cry_4 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5 ;
    wire \b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ;
    wire \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ;
    wire \b2v_inst11.un1_dutycycle_53_i_29 ;
    wire dutycycle_RNIU8G3G_0_2;
    wire bfn_9_15_0_;
    wire \b2v_inst11.mult1_un152_sum_i ;
    wire \b2v_inst11.mult1_un159_sum_cry_1 ;
    wire \b2v_inst11.mult1_un152_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_2 ;
    wire \b2v_inst11.mult1_un152_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_3 ;
    wire \b2v_inst11.mult1_un152_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_4 ;
    wire \b2v_inst11.mult1_un152_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un159_sum_cry_5 ;
    wire \b2v_inst11.mult1_un159_sum_axb_7 ;
    wire \b2v_inst11.mult1_un159_sum_cry_6 ;
    wire \b2v_inst11.mult1_un152_sum_i_0_8 ;
    wire \b2v_inst5.N_51 ;
    wire \b2v_inst5.curr_state_0_1 ;
    wire CONSTANT_ONE_NET;
    wire \b2v_inst36.countZ0Z_2 ;
    wire \b2v_inst36.un12_clk_100khz_11 ;
    wire \b2v_inst36.count_rst_11_cascade_ ;
    wire \b2v_inst36.countZ0Z_3 ;
    wire \b2v_inst36.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst36.countZ0Z_3_cascade_ ;
    wire \b2v_inst36.count_2_3 ;
    wire \b2v_inst36.count_rst_9_cascade_ ;
    wire \b2v_inst36.countZ0Z_5 ;
    wire \b2v_inst36.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst36.countZ0Z_5_cascade_ ;
    wire \b2v_inst36.count_2_5 ;
    wire \b2v_inst36.countZ0Z_7 ;
    wire \b2v_inst36.N_2942_i ;
    wire \b2v_inst36.N_1_i ;
    wire \b2v_inst36.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst36.count_2_7 ;
    wire \b2v_inst36.count_en ;
    wire \b2v_inst36.count_0_sqmuxa ;
    wire \b2v_inst6.count_0_14 ;
    wire \b2v_inst6.countZ0Z_14_cascade_ ;
    wire \b2v_inst6.count_0_6 ;
    wire \b2v_inst5.countZ0Z_1 ;
    wire bfn_11_3_0_;
    wire \b2v_inst5.un2_count_1_axb_2 ;
    wire \b2v_inst5.count_rst_12 ;
    wire \b2v_inst5.un2_count_1_cry_1 ;
    wire \b2v_inst5.countZ0Z_3 ;
    wire \b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ;
    wire \b2v_inst5.un2_count_1_cry_2 ;
    wire \b2v_inst5.un2_count_1_axb_4 ;
    wire \b2v_inst5.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst5.un2_count_1_cry_3 ;
    wire \b2v_inst5.un2_count_1_cry_4 ;
    wire \b2v_inst5.un2_count_1_cry_5 ;
    wire \b2v_inst5.un2_count_1_cry_6 ;
    wire \b2v_inst5.countZ0Z_8 ;
    wire \b2v_inst5.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst5.un2_count_1_cry_7 ;
    wire \b2v_inst5.un2_count_1_cry_8 ;
    wire bfn_11_4_0_;
    wire \b2v_inst5.un2_count_1_cry_9 ;
    wire \b2v_inst5.count_rst_3 ;
    wire \b2v_inst5.un2_count_1_cry_10 ;
    wire \b2v_inst5.countZ0Z_12 ;
    wire \b2v_inst5.count_rst_2 ;
    wire \b2v_inst5.un2_count_1_cry_11 ;
    wire \b2v_inst5.un2_count_1_axb_13 ;
    wire \b2v_inst5.un2_count_1_cry_12_THRU_CO ;
    wire \b2v_inst5.un2_count_1_cry_12 ;
    wire \b2v_inst5.countZ0Z_14 ;
    wire \b2v_inst5.count_rst_0 ;
    wire \b2v_inst5.un2_count_1_cry_13 ;
    wire \b2v_inst5.countZ0Z_15 ;
    wire \b2v_inst5.un2_count_1_cry_14 ;
    wire \b2v_inst5.count_rst ;
    wire \b2v_inst5.count_1_15 ;
    wire \b2v_inst5.count_rst_5_cascade_ ;
    wire \b2v_inst5.un2_count_1_axb_9 ;
    wire \b2v_inst5.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst5.un2_count_1_axb_9_cascade_ ;
    wire \b2v_inst5.count_1_9 ;
    wire \b2v_inst5.count_rst_5 ;
    wire \b2v_inst5.un12_clk_100khz_6 ;
    wire \b2v_inst5.count_rst_4_cascade_ ;
    wire \b2v_inst5.countZ0Z_10 ;
    wire \b2v_inst5.un2_count_1_cry_9_THRU_CO ;
    wire \b2v_inst5.countZ0Z_10_cascade_ ;
    wire \b2v_inst5.count_1_10 ;
    wire \b2v_inst5.un2_count_1_cry_0 ;
    wire \b2v_inst5.N_1_i ;
    wire \b2v_inst5.count_1_0 ;
    wire \b2v_inst5.un2_count_1_axb_5 ;
    wire \b2v_inst5.count_1_6 ;
    wire \b2v_inst5.count_rst_8 ;
    wire \b2v_inst5.countZ0Z_6 ;
    wire \b2v_inst5.count_rst_9 ;
    wire \b2v_inst5.countZ0Z_6_cascade_ ;
    wire \b2v_inst5.count_1_5 ;
    wire \b2v_inst5.un12_clk_100khz_3 ;
    wire \b2v_inst5.un2_count_1_axb_7 ;
    wire \b2v_inst5.count_0_sqmuxa ;
    wire \b2v_inst5.count_1_7 ;
    wire \b2v_inst5.count_rst_7 ;
    wire \b2v_inst5.countZ0Z_11 ;
    wire \b2v_inst5.curr_state_RNIFLPH1Z0Z_1 ;
    wire \b2v_inst5.un12_clk_100khz_2 ;
    wire \b2v_inst11.mult1_un152_sum_s_8 ;
    wire \b2v_inst11.mult1_un110_sum_s_8 ;
    wire \b2v_inst11.mult1_un117_sum_s_8 ;
    wire \b2v_inst11.mult1_un124_sum_s_8 ;
    wire \b2v_inst11.mult1_un145_sum_s_8 ;
    wire \b2v_inst11.mult1_un138_sum_s_8 ;
    wire \b2v_inst11.countZ0Z_0 ;
    wire \b2v_inst11.un1_count_cry_0_i ;
    wire bfn_11_8_0_;
    wire \b2v_inst11.countZ0Z_1 ;
    wire \b2v_inst11.N_5530_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_0 ;
    wire \b2v_inst11.countZ0Z_2 ;
    wire \b2v_inst11.un85_clk_100khz_2 ;
    wire \b2v_inst11.N_5531_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_1 ;
    wire \b2v_inst11.countZ0Z_3 ;
    wire \b2v_inst11.mult1_un145_sum_i_8 ;
    wire \b2v_inst11.N_5532_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_2 ;
    wire \b2v_inst11.countZ0Z_4 ;
    wire \b2v_inst11.mult1_un138_sum_i_8 ;
    wire \b2v_inst11.N_5533_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_3 ;
    wire \b2v_inst11.countZ0Z_5 ;
    wire \b2v_inst11.mult1_un131_sum_i_8 ;
    wire \b2v_inst11.N_5534_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_4 ;
    wire \b2v_inst11.mult1_un124_sum_i_8 ;
    wire \b2v_inst11.countZ0Z_6 ;
    wire \b2v_inst11.N_5535_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_5 ;
    wire \b2v_inst11.countZ0Z_7 ;
    wire \b2v_inst11.mult1_un117_sum_i_8 ;
    wire \b2v_inst11.N_5536_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_6 ;
    wire \b2v_inst11.un85_clk_100khz_cry_7 ;
    wire \b2v_inst11.countZ0Z_8 ;
    wire \b2v_inst11.mult1_un110_sum_i_8 ;
    wire \b2v_inst11.N_5537_i ;
    wire bfn_11_9_0_;
    wire \b2v_inst11.countZ0Z_9 ;
    wire \b2v_inst11.mult1_un103_sum_i_8 ;
    wire \b2v_inst11.N_5538_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_8 ;
    wire \b2v_inst11.countZ0Z_10 ;
    wire \b2v_inst11.N_5539_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_9 ;
    wire \b2v_inst11.countZ0Z_11 ;
    wire \b2v_inst11.N_5540_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_10 ;
    wire \b2v_inst11.countZ0Z_12 ;
    wire \b2v_inst11.N_5541_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_11 ;
    wire \b2v_inst11.countZ0Z_13 ;
    wire \b2v_inst11.N_5542_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_12 ;
    wire \b2v_inst11.countZ0Z_14 ;
    wire \b2v_inst11.N_5543_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_13 ;
    wire \b2v_inst11.countZ0Z_15 ;
    wire \b2v_inst11.N_5544_i ;
    wire \b2v_inst11.un85_clk_100khz_cry_14 ;
    wire \b2v_inst11.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_11_10_0_;
    wire \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \b2v_inst11.mult1_un89_sum_i_8 ;
    wire \b2v_inst11.un85_clk_100khz_1 ;
    wire \b2v_inst11.mult1_un82_sum_i_8 ;
    wire \b2v_inst11.mult1_un89_sum ;
    wire bfn_11_11_0_;
    wire \b2v_inst11.mult1_un82_sum_i ;
    wire \b2v_inst11.mult1_un89_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6 ;
    wire \b2v_inst11.mult1_un89_sum_cry_7 ;
    wire \b2v_inst11.dutycycle ;
    wire \b2v_inst11.mult1_un54_sum ;
    wire \b2v_inst11.mult1_un61_sum_i_8 ;
    wire \b2v_inst11.mult1_un61_sum ;
    wire bfn_11_13_0_;
    wire \b2v_inst11.mult1_un54_sum_i ;
    wire \b2v_inst11.mult1_un61_sum_cry_2 ;
    wire \b2v_inst11.mult1_un54_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_3 ;
    wire \b2v_inst11.mult1_un54_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_4 ;
    wire \b2v_inst11.mult1_un54_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_5 ;
    wire \b2v_inst11.mult1_un54_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un61_sum_cry_6 ;
    wire \b2v_inst11.mult1_un61_sum_axb_8 ;
    wire \b2v_inst11.mult1_un61_sum_cry_7 ;
    wire \b2v_inst11.mult1_un61_sum_s_8_cascade_ ;
    wire V33S_OK_c;
    wire V5S_OK_c;
    wire VCCIN_EN_c;
    wire \b2v_inst6.N_276_0_cascade_ ;
    wire VR_READY_VCCINAUX_c;
    wire VR_READY_VCCIN_c;
    wire \b2v_inst6.N_192_cascade_ ;
    wire \b2v_inst6.delayed_vccin_vccinaux_ok_0 ;
    wire \b2v_inst6.curr_state_RNIUL1J2Z0Z_0_cascade_ ;
    wire \b2v_inst6.N_276_0 ;
    wire N_15_i_0_a4_1_N_3L3_1;
    wire \b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ;
    wire N_222;
    wire \b2v_inst11.dutycycleZ0Z_0 ;
    wire bfn_11_15_0_;
    wire \b2v_inst11.mult1_un159_sum_i ;
    wire \b2v_inst11.mult1_un166_sum_cry_0 ;
    wire \b2v_inst11.mult1_un159_sum_cry_2_s ;
    wire \b2v_inst11.mult1_un166_sum_cry_1 ;
    wire \b2v_inst11.mult1_un159_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un166_sum_cry_2 ;
    wire \b2v_inst11.mult1_un159_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un159_sum_s_7 ;
    wire \b2v_inst11.mult1_un166_sum_cry_3 ;
    wire \b2v_inst11.mult1_un159_sum_cry_5_s ;
    wire G_2836;
    wire \b2v_inst11.mult1_un166_sum_cry_4 ;
    wire \b2v_inst11.mult1_un166_sum_axb_6 ;
    wire \b2v_inst11.mult1_un166_sum_cry_5 ;
    wire \b2v_inst11.un85_clk_100khz_0 ;
    wire bfn_12_1_0_;
    wire \b2v_inst6.countZ0Z_2 ;
    wire \b2v_inst6.un2_count_1_cry_1 ;
    wire \b2v_inst6.un2_count_1_cry_2 ;
    wire \b2v_inst6.un2_count_1_cry_3 ;
    wire \b2v_inst6.un2_count_1_cry_4 ;
    wire \b2v_inst6.countZ0Z_6 ;
    wire \b2v_inst6.count_rst_8 ;
    wire \b2v_inst6.un2_count_1_cry_5 ;
    wire \b2v_inst6.un2_count_1_cry_6 ;
    wire \b2v_inst6.un2_count_1_cry_7 ;
    wire \b2v_inst6.un2_count_1_cry_8 ;
    wire bfn_12_2_0_;
    wire \b2v_inst6.un2_count_1_cry_9 ;
    wire \b2v_inst6.un2_count_1_cry_10 ;
    wire \b2v_inst6.un2_count_1_cry_11 ;
    wire \b2v_inst6.un2_count_1_cry_12 ;
    wire \b2v_inst6.countZ0Z_14 ;
    wire \b2v_inst6.count_rst_0 ;
    wire \b2v_inst6.un2_count_1_cry_13 ;
    wire \b2v_inst6.un2_count_1_cry_14 ;
    wire \b2v_inst6.count_0_13 ;
    wire \b2v_inst6.count_rst_1 ;
    wire \b2v_inst6.countZ0Z_13 ;
    wire \b2v_inst6.count_0_5 ;
    wire \b2v_inst6.un2_count_1_cry_4_THRU_CO ;
    wire \b2v_inst6.countZ0Z_5_cascade_ ;
    wire \b2v_inst6.count_rst_9 ;
    wire \b2v_inst6.count_rst_5 ;
    wire \b2v_inst6.countZ0Z_9_cascade_ ;
    wire \b2v_inst6.countZ0Z_5 ;
    wire \b2v_inst6.countZ0Z_9 ;
    wire \b2v_inst6.un2_count_1_cry_8_THRU_CO ;
    wire \b2v_inst6.count_0_9 ;
    wire \b2v_inst6.countZ0Z_10 ;
    wire \b2v_inst6.countZ0Z_10_cascade_ ;
    wire \b2v_inst6.count_0_12 ;
    wire \b2v_inst6.count_rst_2 ;
    wire \b2v_inst6.countZ0Z_12 ;
    wire \b2v_inst6.count_rst_10_cascade_ ;
    wire \b2v_inst6.countZ0Z_4 ;
    wire \b2v_inst6.un2_count_1_cry_3_THRU_CO ;
    wire \b2v_inst6.countZ0Z_4_cascade_ ;
    wire \b2v_inst6.count_0_4 ;
    wire \b2v_inst6.count_rst_4 ;
    wire \b2v_inst6.count_0_10 ;
    wire \b2v_inst6.un2_count_1_cry_6_THRU_CO ;
    wire \b2v_inst6.count_0_7 ;
    wire \b2v_inst6.count_rst_7_cascade_ ;
    wire \b2v_inst6.countZ0Z_7 ;
    wire \b2v_inst6.count_rst ;
    wire \b2v_inst6.count_0_15 ;
    wire \b2v_inst6.count_rst_12 ;
    wire \b2v_inst6.count_0_2 ;
    wire \b2v_inst6.count_rst_6 ;
    wire \b2v_inst6.countZ0Z_8 ;
    wire \b2v_inst6.countZ0Z_8_cascade_ ;
    wire \b2v_inst6.un2_count_1_cry_7_THRU_CO ;
    wire \b2v_inst6.count_0_8 ;
    wire \b2v_inst6.count_rst_11_cascade_ ;
    wire \b2v_inst6.countZ0Z_3 ;
    wire \b2v_inst6.un2_count_1_cry_2_THRU_CO ;
    wire \b2v_inst6.countZ0Z_3_cascade_ ;
    wire \b2v_inst6.count_0_3 ;
    wire \b2v_inst6.un2_count_1_cry_10_THRU_CO ;
    wire \b2v_inst6.N_394_cascade_ ;
    wire \b2v_inst6.count_0_11 ;
    wire \b2v_inst6.count_rst_3_cascade_ ;
    wire \b2v_inst6.un2_count_1_axb_1 ;
    wire \b2v_inst6.un2_count_1_axb_1_cascade_ ;
    wire V1P8A_OK_c;
    wire V33A_OK_c;
    wire V5A_OK_c;
    wire VCCST_CPU_OK_c;
    wire N_1661;
    wire \b2v_inst6.count_0_1 ;
    wire \b2v_inst6.count_RNI_0_1 ;
    wire \b2v_inst6.countZ0Z_15 ;
    wire \b2v_inst6.countZ0Z_1_cascade_ ;
    wire \b2v_inst6.countZ0Z_11 ;
    wire \b2v_inst6.count_1_i_a3_8_0 ;
    wire \b2v_inst6.count_1_i_a3_9_0 ;
    wire \b2v_inst6.count_1_i_a3_7_0_cascade_ ;
    wire \b2v_inst6.count_1_i_a3_10_0 ;
    wire \b2v_inst6.N_389 ;
    wire \b2v_inst6.N_389_cascade_ ;
    wire \b2v_inst11.mult1_un75_sum_i_8 ;
    wire \b2v_inst11.mult1_un96_sum_i_8 ;
    wire \b2v_inst11.mult1_un96_sum_i ;
    wire \b2v_inst11.mult1_un68_sum_i_8 ;
    wire \b2v_inst6.count_en ;
    wire \b2v_inst6.count_RNIM2CM2Z0Z_0 ;
    wire \b2v_inst6.count_en_cascade_ ;
    wire \b2v_inst6.count_0_0 ;
    wire \b2v_inst6.countZ0Z_0 ;
    wire \b2v_inst11.mult1_un96_sum ;
    wire bfn_12_10_0_;
    wire \b2v_inst11.mult1_un89_sum_i ;
    wire \b2v_inst11.mult1_un96_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_2 ;
    wire \b2v_inst11.mult1_un89_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_3 ;
    wire \b2v_inst11.mult1_un89_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_4 ;
    wire \b2v_inst11.mult1_un89_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un96_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un103_sum_axb_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_6 ;
    wire \b2v_inst11.mult1_un96_sum_axb_8 ;
    wire \b2v_inst11.mult1_un96_sum_cry_7 ;
    wire \b2v_inst11.mult1_un96_sum_s_8 ;
    wire \b2v_inst11.mult1_un89_sum_s_8 ;
    wire \b2v_inst11.mult1_un89_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un82_sum ;
    wire bfn_12_11_0_;
    wire \b2v_inst11.mult1_un75_sum_i ;
    wire \b2v_inst11.mult1_un82_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_2 ;
    wire \b2v_inst11.mult1_un82_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_3 ;
    wire \b2v_inst11.mult1_un82_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_4 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un82_sum_cry_5 ;
    wire \b2v_inst11.mult1_un89_sum_axb_8 ;
    wire \b2v_inst11.mult1_un82_sum_cry_6 ;
    wire \b2v_inst11.mult1_un82_sum_cry_7 ;
    wire \b2v_inst11.mult1_un82_sum_s_8 ;
    wire \b2v_inst11.mult1_un82_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un82_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un75_sum ;
    wire bfn_12_12_0_;
    wire \b2v_inst11.mult1_un68_sum_i ;
    wire \b2v_inst11.mult1_un75_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_2 ;
    wire \b2v_inst11.mult1_un75_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_3 ;
    wire \b2v_inst11.mult1_un75_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_4 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un75_sum_cry_5 ;
    wire \b2v_inst11.mult1_un68_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un82_sum_axb_8 ;
    wire \b2v_inst11.mult1_un75_sum_cry_6 ;
    wire \b2v_inst11.mult1_un75_sum_cry_7 ;
    wire \b2v_inst11.mult1_un75_sum_s_8 ;
    wire \b2v_inst11.mult1_un75_sum_s_8_cascade_ ;
    wire \b2v_inst11.mult1_un75_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un68_sum ;
    wire bfn_12_13_0_;
    wire \b2v_inst11.mult1_un61_sum_i ;
    wire \b2v_inst11.mult1_un68_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_2 ;
    wire \b2v_inst11.mult1_un61_sum_cry_3_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_3 ;
    wire \b2v_inst11.mult1_un61_sum_cry_4_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_4 ;
    wire \b2v_inst11.mult1_un61_sum_s_8 ;
    wire \b2v_inst11.mult1_un61_sum_cry_5_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un68_sum_cry_5 ;
    wire \b2v_inst11.mult1_un61_sum_cry_6_s ;
    wire \b2v_inst11.mult1_un61_sum_i_0_8 ;
    wire \b2v_inst11.mult1_un75_sum_axb_8 ;
    wire \b2v_inst11.mult1_un68_sum_cry_6 ;
    wire \b2v_inst11.mult1_un68_sum_axb_8 ;
    wire \b2v_inst11.mult1_un68_sum_cry_7 ;
    wire \b2v_inst11.mult1_un68_sum_s_8 ;
    wire \b2v_inst11.mult1_un54_sum_s_8 ;
    wire \b2v_inst11.mult1_un54_sum_i_8 ;
    wire \b2v_inst6.N_192 ;
    wire \b2v_inst6.curr_stateZ0Z_0_cascade_ ;
    wire \b2v_inst6.count_0_sqmuxa ;
    wire \b2v_inst6.curr_state_1_0 ;
    wire SYNTHESIZED_WIRE_1keep_3;
    wire \b2v_inst6.curr_stateZ0Z_0 ;
    wire \b2v_inst6.curr_stateZ0Z_1_cascade_ ;
    wire \b2v_inst6.curr_state_RNIUL1J2Z0Z_0 ;
    wire \b2v_inst6.curr_state_7_0 ;
    wire \b2v_inst6.N_2937_i ;
    wire \b2v_inst6.curr_stateZ0Z_1 ;
    wire \b2v_inst6.N_394 ;
    wire \b2v_inst6.m6_i_a3 ;
    wire \b2v_inst6.N_241 ;
    wire \b2v_inst6.m6_i_a3_cascade_ ;
    wire \b2v_inst6.curr_state_1_1 ;
    wire FPGA_OSC_0_c_g;
    wire N_606_g;
    wire _gnd_net_;

    PRE_IO_GBUF FPGA_OSC_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__37127),
            .GLOBALBUFFEROUTPUT(FPGA_OSC_0_c_g));
    IO_PAD FPGA_OSC_ibuf_gb_io_iopad (
            .OE(N__37129),
            .DIN(N__37128),
            .DOUT(N__37127),
            .PACKAGEPIN(FPGA_OSC));
    defparam FPGA_OSC_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam FPGA_OSC_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO FPGA_OSC_ibuf_gb_io_preio (
            .PADOEN(N__37129),
            .PADOUT(N__37128),
            .PADIN(N__37127),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V1P8A_OK_ibuf_iopad (
            .OE(N__37118),
            .DIN(N__37117),
            .DOUT(N__37116),
            .PACKAGEPIN(V1P8A_OK));
    defparam V1P8A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V1P8A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V1P8A_OK_ibuf_preio (
            .PADOEN(N__37118),
            .PADOUT(N__37117),
            .PADIN(N__37116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V1P8A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5A_OK_ibuf_iopad (
            .OE(N__37109),
            .DIN(N__37108),
            .DOUT(N__37107),
            .PACKAGEPIN(V5A_OK));
    defparam V5A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V5A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V5A_OK_ibuf_preio (
            .PADOEN(N__37109),
            .PADOUT(N__37108),
            .PADIN(N__37107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCH_PWROK_obuf_iopad (
            .OE(N__37100),
            .DIN(N__37099),
            .DOUT(N__37098),
            .PACKAGEPIN(PCH_PWROK));
    defparam PCH_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCH_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCH_PWROK_obuf_preio (
            .PADOEN(N__37100),
            .PADOUT(N__37099),
            .PADIN(N__37098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18636),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCIN_EN_obuf_iopad (
            .OE(N__37091),
            .DIN(N__37090),
            .DOUT(N__37089),
            .PACKAGEPIN(VCCIN_EN));
    defparam VCCIN_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCIN_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCIN_EN_obuf_preio (
            .PADOEN(N__37091),
            .PADOUT(N__37090),
            .PADIN(N__37089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33399),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33S_OK_ibuf_iopad (
            .OE(N__37082),
            .DIN(N__37081),
            .DOUT(N__37080),
            .PACKAGEPIN(V33S_OK));
    defparam V33S_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33S_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33S_OK_ibuf_preio (
            .PADOEN(N__37082),
            .PADOUT(N__37081),
            .PADIN(N__37080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33S_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5S_ENn_obuf_iopad (
            .OE(N__37073),
            .DIN(N__37072),
            .DOUT(N__37071),
            .PACKAGEPIN(V5S_ENn));
    defparam V5S_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V5S_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V5S_ENn_obuf_preio (
            .PADOEN(N__37073),
            .PADOUT(N__37072),
            .PADIN(N__37071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33801),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_S4n_ibuf_iopad (
            .OE(N__37064),
            .DIN(N__37063),
            .DOUT(N__37062),
            .PACKAGEPIN(SLP_S4n));
    defparam SLP_S4n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_S4n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_S4n_ibuf_preio (
            .PADOEN(N__37064),
            .PADOUT(N__37063),
            .PADIN(N__37062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SLP_S4n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VR_READY_VCCINAUX_ibuf_iopad (
            .OE(N__37055),
            .DIN(N__37054),
            .DOUT(N__37053),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam VR_READY_VCCINAUX_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VR_READY_VCCINAUX_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VR_READY_VCCINAUX_ibuf_preio (
            .PADOEN(N__37055),
            .PADOUT(N__37054),
            .PADIN(N__37053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VR_READY_VCCINAUX_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_S3n_ibuf_iopad (
            .OE(N__37046),
            .DIN(N__37045),
            .DOUT(N__37044),
            .PACKAGEPIN(SLP_S3n));
    defparam SLP_S3n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_S3n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_S3n_ibuf_preio (
            .PADOEN(N__37046),
            .PADOUT(N__37045),
            .PADIN(N__37044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SLP_S3n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_PWRGD_obuf_iopad (
            .OE(N__37037),
            .DIN(N__37036),
            .DOUT(N__37035),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam VCCST_PWRGD_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_PWRGD_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCST_PWRGD_obuf_preio (
            .PADOEN(N__37037),
            .PADOUT(N__37036),
            .PADIN(N__37035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18640),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD HDA_SDO_ATP_obuf_iopad (
            .OE(N__37028),
            .DIN(N__37027),
            .DOUT(N__37026),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam HDA_SDO_ATP_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HDA_SDO_ATP_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HDA_SDO_ATP_obuf_preio (
            .PADOEN(N__37028),
            .PADOUT(N__37027),
            .PADIN(N__37026),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20227),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_EN_obuf_iopad (
            .OE(N__37019),
            .DIN(N__37018),
            .DOUT(N__37017),
            .PACKAGEPIN(VCCST_EN));
    defparam VCCST_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCST_EN_obuf_preio (
            .PADOEN(N__37019),
            .PADOUT(N__37018),
            .PADIN(N__37017),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19873),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VPP_OK_ibuf_iopad (
            .OE(N__37010),
            .DIN(N__37009),
            .DOUT(N__37008),
            .PACKAGEPIN(VPP_OK));
    defparam VPP_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VPP_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VPP_OK_ibuf_preio (
            .PADOEN(N__37010),
            .PADOUT(N__37009),
            .PADIN(N__37008),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VPP_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO_FPGA_SoC_1_ibuf_iopad (
            .OE(N__37001),
            .DIN(N__37000),
            .DOUT(N__36999),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam GPIO_FPGA_SoC_1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO_FPGA_SoC_1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO GPIO_FPGA_SoC_1_ibuf_preio (
            .PADOEN(N__37001),
            .PADOUT(N__37000),
            .PADIN(N__36999),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(GPIO_FPGA_SoC_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_CPU_OK_ibuf_iopad (
            .OE(N__36992),
            .DIN(N__36991),
            .DOUT(N__36990),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam VCCST_CPU_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_CPU_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VCCST_CPU_OK_ibuf_preio (
            .PADOEN(N__36992),
            .PADOUT(N__36991),
            .PADIN(N__36990),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VCCST_CPU_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD GPIO_FPGA_SoC_4_ibuf_iopad (
            .OE(N__36983),
            .DIN(N__36982),
            .DOUT(N__36981),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam GPIO_FPGA_SoC_4_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam GPIO_FPGA_SoC_4_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO GPIO_FPGA_SoC_4_ibuf_preio (
            .PADOEN(N__36983),
            .PADOUT(N__36982),
            .PADIN(N__36981),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(GPIO_FPGA_SoC_4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VPP_EN_obuf_iopad (
            .OE(N__36974),
            .DIN(N__36973),
            .DOUT(N__36972),
            .PACKAGEPIN(VPP_EN));
    defparam VPP_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VPP_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VPP_EN_obuf_preio (
            .PADOEN(N__36974),
            .PADOUT(N__36973),
            .PADIN(N__36972),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14902),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWRBTN_LED_obuf_iopad (
            .OE(N__36965),
            .DIN(N__36964),
            .DOUT(N__36963),
            .PACKAGEPIN(PWRBTN_LED));
    defparam PWRBTN_LED_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWRBTN_LED_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PWRBTN_LED_obuf_preio (
            .PADOEN(N__36965),
            .PADOUT(N__36964),
            .PADIN(N__36963),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24946),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33S_ENn_obuf_iopad (
            .OE(N__36956),
            .DIN(N__36955),
            .DOUT(N__36954),
            .PACKAGEPIN(V33S_ENn));
    defparam V33S_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V33S_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V33S_ENn_obuf_preio (
            .PADOEN(N__36956),
            .PADOUT(N__36955),
            .PADIN(N__36954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33792),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RSMRSTn_obuf_iopad (
            .OE(N__36947),
            .DIN(N__36946),
            .DOUT(N__36945),
            .PACKAGEPIN(RSMRSTn));
    defparam RSMRSTn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RSMRSTn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RSMRSTn_obuf_preio (
            .PADOEN(N__36947),
            .PADOUT(N__36946),
            .PADIN(N__36945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23911),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V1P8A_EN_obuf_iopad (
            .OE(N__36938),
            .DIN(N__36937),
            .DOUT(N__36936),
            .PACKAGEPIN(V1P8A_EN));
    defparam V1P8A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V1P8A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V1P8A_EN_obuf_preio (
            .PADOEN(N__36938),
            .PADOUT(N__36937),
            .PADIN(N__36936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VDDQ_OK_ibuf_iopad (
            .OE(N__36929),
            .DIN(N__36928),
            .DOUT(N__36927),
            .PACKAGEPIN(VDDQ_OK));
    defparam VDDQ_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VDDQ_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VDDQ_OK_ibuf_preio (
            .PADOEN(N__36929),
            .PADOUT(N__36928),
            .PADIN(N__36927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VDDQ_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DSW_PWROK_obuf_iopad (
            .OE(N__36920),
            .DIN(N__36919),
            .DOUT(N__36918),
            .PACKAGEPIN(DSW_PWROK));
    defparam DSW_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DSW_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DSW_PWROK_obuf_preio (
            .PADOEN(N__36920),
            .PADOUT(N__36919),
            .PADIN(N__36918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22351),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SYS_PWROK_obuf_iopad (
            .OE(N__36911),
            .DIN(N__36910),
            .DOUT(N__36909),
            .PACKAGEPIN(SYS_PWROK));
    defparam SYS_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SYS_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SYS_PWROK_obuf_preio (
            .PADOEN(N__36911),
            .PADOUT(N__36910),
            .PADIN(N__36909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18635),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33DSW_OK_ibuf_iopad (
            .OE(N__36902),
            .DIN(N__36901),
            .DOUT(N__36900),
            .PACKAGEPIN(V33DSW_OK));
    defparam V33DSW_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33DSW_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33DSW_OK_ibuf_preio (
            .PADOEN(N__36902),
            .PADOUT(N__36901),
            .PADIN(N__36900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33DSW_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VR_READY_VCCIN_ibuf_iopad (
            .OE(N__36893),
            .DIN(N__36892),
            .DOUT(N__36891),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam VR_READY_VCCIN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VR_READY_VCCIN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VR_READY_VCCIN_ibuf_preio (
            .PADOEN(N__36893),
            .PADOUT(N__36892),
            .PADIN(N__36891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VR_READY_VCCIN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VDDQ_EN_obuf_iopad (
            .OE(N__36884),
            .DIN(N__36883),
            .DOUT(N__36882),
            .PACKAGEPIN(VDDQ_EN));
    defparam VDDQ_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VDDQ_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VDDQ_EN_obuf_preio (
            .PADOEN(N__36884),
            .PADOUT(N__36883),
            .PADIN(N__36882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16966),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5A_EN_obuf_iopad (
            .OE(N__36875),
            .DIN(N__36874),
            .DOUT(N__36873),
            .PACKAGEPIN(V5A_EN));
    defparam V5A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V5A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V5A_EN_obuf_preio (
            .PADOEN(N__36875),
            .PADOUT(N__36874),
            .PADIN(N__36873),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__30442),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCINAUX_EN_obuf_iopad (
            .OE(N__36866),
            .DIN(N__36865),
            .DOUT(N__36864),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam VCCINAUX_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCINAUX_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCINAUX_EN_obuf_preio (
            .PADOEN(N__36866),
            .PADOUT(N__36865),
            .PADIN(N__36864),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33403),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33A_ENn_obuf_iopad (
            .OE(N__36857),
            .DIN(N__36856),
            .DOUT(N__36855),
            .PACKAGEPIN(V33A_ENn));
    defparam V33A_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V33A_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V33A_ENn_obuf_preio (
            .PADOEN(N__36857),
            .PADOUT(N__36856),
            .PADIN(N__36855),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5S_OK_ibuf_iopad (
            .OE(N__36848),
            .DIN(N__36847),
            .DOUT(N__36846),
            .PACKAGEPIN(V5S_OK));
    defparam V5S_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V5S_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V5S_OK_ibuf_preio (
            .PADOEN(N__36848),
            .PADOUT(N__36847),
            .PADIN(N__36846),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5S_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33A_OK_ibuf_iopad (
            .OE(N__36839),
            .DIN(N__36838),
            .DOUT(N__36837),
            .PACKAGEPIN(V33A_OK));
    defparam V33A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33A_OK_ibuf_preio (
            .PADOEN(N__36839),
            .PADOUT(N__36838),
            .PADIN(N__36837),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__8612 (
            .O(N__36820),
            .I(N__36814));
    InMux I__8611 (
            .O(N__36819),
            .I(N__36807));
    InMux I__8610 (
            .O(N__36818),
            .I(N__36807));
    InMux I__8609 (
            .O(N__36817),
            .I(N__36807));
    LocalMux I__8608 (
            .O(N__36814),
            .I(\b2v_inst6.N_2937_i ));
    LocalMux I__8607 (
            .O(N__36807),
            .I(\b2v_inst6.N_2937_i ));
    InMux I__8606 (
            .O(N__36802),
            .I(N__36793));
    InMux I__8605 (
            .O(N__36801),
            .I(N__36793));
    InMux I__8604 (
            .O(N__36800),
            .I(N__36793));
    LocalMux I__8603 (
            .O(N__36793),
            .I(\b2v_inst6.curr_stateZ0Z_1 ));
    CascadeMux I__8602 (
            .O(N__36790),
            .I(N__36784));
    CascadeMux I__8601 (
            .O(N__36789),
            .I(N__36778));
    CascadeMux I__8600 (
            .O(N__36788),
            .I(N__36775));
    InMux I__8599 (
            .O(N__36787),
            .I(N__36765));
    InMux I__8598 (
            .O(N__36784),
            .I(N__36765));
    InMux I__8597 (
            .O(N__36783),
            .I(N__36762));
    InMux I__8596 (
            .O(N__36782),
            .I(N__36753));
    InMux I__8595 (
            .O(N__36781),
            .I(N__36753));
    InMux I__8594 (
            .O(N__36778),
            .I(N__36742));
    InMux I__8593 (
            .O(N__36775),
            .I(N__36742));
    InMux I__8592 (
            .O(N__36774),
            .I(N__36742));
    InMux I__8591 (
            .O(N__36773),
            .I(N__36742));
    InMux I__8590 (
            .O(N__36772),
            .I(N__36742));
    InMux I__8589 (
            .O(N__36771),
            .I(N__36737));
    InMux I__8588 (
            .O(N__36770),
            .I(N__36737));
    LocalMux I__8587 (
            .O(N__36765),
            .I(N__36732));
    LocalMux I__8586 (
            .O(N__36762),
            .I(N__36732));
    InMux I__8585 (
            .O(N__36761),
            .I(N__36727));
    InMux I__8584 (
            .O(N__36760),
            .I(N__36727));
    InMux I__8583 (
            .O(N__36759),
            .I(N__36722));
    InMux I__8582 (
            .O(N__36758),
            .I(N__36722));
    LocalMux I__8581 (
            .O(N__36753),
            .I(N__36713));
    LocalMux I__8580 (
            .O(N__36742),
            .I(N__36713));
    LocalMux I__8579 (
            .O(N__36737),
            .I(N__36713));
    Span12Mux_s8_v I__8578 (
            .O(N__36732),
            .I(N__36713));
    LocalMux I__8577 (
            .O(N__36727),
            .I(\b2v_inst6.N_394 ));
    LocalMux I__8576 (
            .O(N__36722),
            .I(\b2v_inst6.N_394 ));
    Odrv12 I__8575 (
            .O(N__36713),
            .I(\b2v_inst6.N_394 ));
    InMux I__8574 (
            .O(N__36706),
            .I(N__36703));
    LocalMux I__8573 (
            .O(N__36703),
            .I(\b2v_inst6.m6_i_a3 ));
    CascadeMux I__8572 (
            .O(N__36700),
            .I(N__36696));
    InMux I__8571 (
            .O(N__36699),
            .I(N__36693));
    InMux I__8570 (
            .O(N__36696),
            .I(N__36689));
    LocalMux I__8569 (
            .O(N__36693),
            .I(N__36686));
    InMux I__8568 (
            .O(N__36692),
            .I(N__36683));
    LocalMux I__8567 (
            .O(N__36689),
            .I(N__36678));
    Span4Mux_v I__8566 (
            .O(N__36686),
            .I(N__36678));
    LocalMux I__8565 (
            .O(N__36683),
            .I(\b2v_inst6.N_241 ));
    Odrv4 I__8564 (
            .O(N__36678),
            .I(\b2v_inst6.N_241 ));
    CascadeMux I__8563 (
            .O(N__36673),
            .I(\b2v_inst6.m6_i_a3_cascade_ ));
    InMux I__8562 (
            .O(N__36670),
            .I(N__36667));
    LocalMux I__8561 (
            .O(N__36667),
            .I(\b2v_inst6.curr_state_1_1 ));
    ClkMux I__8560 (
            .O(N__36664),
            .I(N__36415));
    ClkMux I__8559 (
            .O(N__36663),
            .I(N__36415));
    ClkMux I__8558 (
            .O(N__36662),
            .I(N__36415));
    ClkMux I__8557 (
            .O(N__36661),
            .I(N__36415));
    ClkMux I__8556 (
            .O(N__36660),
            .I(N__36415));
    ClkMux I__8555 (
            .O(N__36659),
            .I(N__36415));
    ClkMux I__8554 (
            .O(N__36658),
            .I(N__36415));
    ClkMux I__8553 (
            .O(N__36657),
            .I(N__36415));
    ClkMux I__8552 (
            .O(N__36656),
            .I(N__36415));
    ClkMux I__8551 (
            .O(N__36655),
            .I(N__36415));
    ClkMux I__8550 (
            .O(N__36654),
            .I(N__36415));
    ClkMux I__8549 (
            .O(N__36653),
            .I(N__36415));
    ClkMux I__8548 (
            .O(N__36652),
            .I(N__36415));
    ClkMux I__8547 (
            .O(N__36651),
            .I(N__36415));
    ClkMux I__8546 (
            .O(N__36650),
            .I(N__36415));
    ClkMux I__8545 (
            .O(N__36649),
            .I(N__36415));
    ClkMux I__8544 (
            .O(N__36648),
            .I(N__36415));
    ClkMux I__8543 (
            .O(N__36647),
            .I(N__36415));
    ClkMux I__8542 (
            .O(N__36646),
            .I(N__36415));
    ClkMux I__8541 (
            .O(N__36645),
            .I(N__36415));
    ClkMux I__8540 (
            .O(N__36644),
            .I(N__36415));
    ClkMux I__8539 (
            .O(N__36643),
            .I(N__36415));
    ClkMux I__8538 (
            .O(N__36642),
            .I(N__36415));
    ClkMux I__8537 (
            .O(N__36641),
            .I(N__36415));
    ClkMux I__8536 (
            .O(N__36640),
            .I(N__36415));
    ClkMux I__8535 (
            .O(N__36639),
            .I(N__36415));
    ClkMux I__8534 (
            .O(N__36638),
            .I(N__36415));
    ClkMux I__8533 (
            .O(N__36637),
            .I(N__36415));
    ClkMux I__8532 (
            .O(N__36636),
            .I(N__36415));
    ClkMux I__8531 (
            .O(N__36635),
            .I(N__36415));
    ClkMux I__8530 (
            .O(N__36634),
            .I(N__36415));
    ClkMux I__8529 (
            .O(N__36633),
            .I(N__36415));
    ClkMux I__8528 (
            .O(N__36632),
            .I(N__36415));
    ClkMux I__8527 (
            .O(N__36631),
            .I(N__36415));
    ClkMux I__8526 (
            .O(N__36630),
            .I(N__36415));
    ClkMux I__8525 (
            .O(N__36629),
            .I(N__36415));
    ClkMux I__8524 (
            .O(N__36628),
            .I(N__36415));
    ClkMux I__8523 (
            .O(N__36627),
            .I(N__36415));
    ClkMux I__8522 (
            .O(N__36626),
            .I(N__36415));
    ClkMux I__8521 (
            .O(N__36625),
            .I(N__36415));
    ClkMux I__8520 (
            .O(N__36624),
            .I(N__36415));
    ClkMux I__8519 (
            .O(N__36623),
            .I(N__36415));
    ClkMux I__8518 (
            .O(N__36622),
            .I(N__36415));
    ClkMux I__8517 (
            .O(N__36621),
            .I(N__36415));
    ClkMux I__8516 (
            .O(N__36620),
            .I(N__36415));
    ClkMux I__8515 (
            .O(N__36619),
            .I(N__36415));
    ClkMux I__8514 (
            .O(N__36618),
            .I(N__36415));
    ClkMux I__8513 (
            .O(N__36617),
            .I(N__36415));
    ClkMux I__8512 (
            .O(N__36616),
            .I(N__36415));
    ClkMux I__8511 (
            .O(N__36615),
            .I(N__36415));
    ClkMux I__8510 (
            .O(N__36614),
            .I(N__36415));
    ClkMux I__8509 (
            .O(N__36613),
            .I(N__36415));
    ClkMux I__8508 (
            .O(N__36612),
            .I(N__36415));
    ClkMux I__8507 (
            .O(N__36611),
            .I(N__36415));
    ClkMux I__8506 (
            .O(N__36610),
            .I(N__36415));
    ClkMux I__8505 (
            .O(N__36609),
            .I(N__36415));
    ClkMux I__8504 (
            .O(N__36608),
            .I(N__36415));
    ClkMux I__8503 (
            .O(N__36607),
            .I(N__36415));
    ClkMux I__8502 (
            .O(N__36606),
            .I(N__36415));
    ClkMux I__8501 (
            .O(N__36605),
            .I(N__36415));
    ClkMux I__8500 (
            .O(N__36604),
            .I(N__36415));
    ClkMux I__8499 (
            .O(N__36603),
            .I(N__36415));
    ClkMux I__8498 (
            .O(N__36602),
            .I(N__36415));
    ClkMux I__8497 (
            .O(N__36601),
            .I(N__36415));
    ClkMux I__8496 (
            .O(N__36600),
            .I(N__36415));
    ClkMux I__8495 (
            .O(N__36599),
            .I(N__36415));
    ClkMux I__8494 (
            .O(N__36598),
            .I(N__36415));
    ClkMux I__8493 (
            .O(N__36597),
            .I(N__36415));
    ClkMux I__8492 (
            .O(N__36596),
            .I(N__36415));
    ClkMux I__8491 (
            .O(N__36595),
            .I(N__36415));
    ClkMux I__8490 (
            .O(N__36594),
            .I(N__36415));
    ClkMux I__8489 (
            .O(N__36593),
            .I(N__36415));
    ClkMux I__8488 (
            .O(N__36592),
            .I(N__36415));
    ClkMux I__8487 (
            .O(N__36591),
            .I(N__36415));
    ClkMux I__8486 (
            .O(N__36590),
            .I(N__36415));
    ClkMux I__8485 (
            .O(N__36589),
            .I(N__36415));
    ClkMux I__8484 (
            .O(N__36588),
            .I(N__36415));
    ClkMux I__8483 (
            .O(N__36587),
            .I(N__36415));
    ClkMux I__8482 (
            .O(N__36586),
            .I(N__36415));
    ClkMux I__8481 (
            .O(N__36585),
            .I(N__36415));
    ClkMux I__8480 (
            .O(N__36584),
            .I(N__36415));
    ClkMux I__8479 (
            .O(N__36583),
            .I(N__36415));
    ClkMux I__8478 (
            .O(N__36582),
            .I(N__36415));
    GlobalMux I__8477 (
            .O(N__36415),
            .I(N__36412));
    gio2CtrlBuf I__8476 (
            .O(N__36412),
            .I(FPGA_OSC_0_c_g));
    InMux I__8475 (
            .O(N__36409),
            .I(N__36397));
    InMux I__8474 (
            .O(N__36408),
            .I(N__36394));
    InMux I__8473 (
            .O(N__36407),
            .I(N__36391));
    InMux I__8472 (
            .O(N__36406),
            .I(N__36384));
    InMux I__8471 (
            .O(N__36405),
            .I(N__36384));
    InMux I__8470 (
            .O(N__36404),
            .I(N__36384));
    InMux I__8469 (
            .O(N__36403),
            .I(N__36381));
    InMux I__8468 (
            .O(N__36402),
            .I(N__36376));
    InMux I__8467 (
            .O(N__36401),
            .I(N__36376));
    InMux I__8466 (
            .O(N__36400),
            .I(N__36373));
    LocalMux I__8465 (
            .O(N__36397),
            .I(N__36370));
    LocalMux I__8464 (
            .O(N__36394),
            .I(N__36352));
    LocalMux I__8463 (
            .O(N__36391),
            .I(N__36349));
    LocalMux I__8462 (
            .O(N__36384),
            .I(N__36346));
    LocalMux I__8461 (
            .O(N__36381),
            .I(N__36343));
    LocalMux I__8460 (
            .O(N__36376),
            .I(N__36340));
    LocalMux I__8459 (
            .O(N__36373),
            .I(N__36337));
    Glb2LocalMux I__8458 (
            .O(N__36370),
            .I(N__36292));
    CEMux I__8457 (
            .O(N__36369),
            .I(N__36292));
    CEMux I__8456 (
            .O(N__36368),
            .I(N__36292));
    CEMux I__8455 (
            .O(N__36367),
            .I(N__36292));
    CEMux I__8454 (
            .O(N__36366),
            .I(N__36292));
    CEMux I__8453 (
            .O(N__36365),
            .I(N__36292));
    CEMux I__8452 (
            .O(N__36364),
            .I(N__36292));
    CEMux I__8451 (
            .O(N__36363),
            .I(N__36292));
    CEMux I__8450 (
            .O(N__36362),
            .I(N__36292));
    CEMux I__8449 (
            .O(N__36361),
            .I(N__36292));
    CEMux I__8448 (
            .O(N__36360),
            .I(N__36292));
    CEMux I__8447 (
            .O(N__36359),
            .I(N__36292));
    CEMux I__8446 (
            .O(N__36358),
            .I(N__36292));
    CEMux I__8445 (
            .O(N__36357),
            .I(N__36292));
    CEMux I__8444 (
            .O(N__36356),
            .I(N__36292));
    CEMux I__8443 (
            .O(N__36355),
            .I(N__36292));
    Glb2LocalMux I__8442 (
            .O(N__36352),
            .I(N__36292));
    Glb2LocalMux I__8441 (
            .O(N__36349),
            .I(N__36292));
    Glb2LocalMux I__8440 (
            .O(N__36346),
            .I(N__36292));
    Glb2LocalMux I__8439 (
            .O(N__36343),
            .I(N__36292));
    Glb2LocalMux I__8438 (
            .O(N__36340),
            .I(N__36292));
    Glb2LocalMux I__8437 (
            .O(N__36337),
            .I(N__36292));
    GlobalMux I__8436 (
            .O(N__36292),
            .I(N__36289));
    gio2CtrlBuf I__8435 (
            .O(N__36289),
            .I(N_606_g));
    InMux I__8434 (
            .O(N__36286),
            .I(\b2v_inst11.mult1_un68_sum_cry_5 ));
    InMux I__8433 (
            .O(N__36283),
            .I(N__36280));
    LocalMux I__8432 (
            .O(N__36280),
            .I(N__36277));
    Odrv4 I__8431 (
            .O(N__36277),
            .I(\b2v_inst11.mult1_un61_sum_cry_6_s ));
    CascadeMux I__8430 (
            .O(N__36274),
            .I(N__36270));
    CascadeMux I__8429 (
            .O(N__36273),
            .I(N__36266));
    InMux I__8428 (
            .O(N__36270),
            .I(N__36259));
    InMux I__8427 (
            .O(N__36269),
            .I(N__36259));
    InMux I__8426 (
            .O(N__36266),
            .I(N__36259));
    LocalMux I__8425 (
            .O(N__36259),
            .I(\b2v_inst11.mult1_un61_sum_i_0_8 ));
    CascadeMux I__8424 (
            .O(N__36256),
            .I(N__36253));
    InMux I__8423 (
            .O(N__36253),
            .I(N__36250));
    LocalMux I__8422 (
            .O(N__36250),
            .I(\b2v_inst11.mult1_un75_sum_axb_8 ));
    InMux I__8421 (
            .O(N__36247),
            .I(\b2v_inst11.mult1_un68_sum_cry_6 ));
    CascadeMux I__8420 (
            .O(N__36244),
            .I(N__36241));
    InMux I__8419 (
            .O(N__36241),
            .I(N__36238));
    LocalMux I__8418 (
            .O(N__36238),
            .I(\b2v_inst11.mult1_un68_sum_axb_8 ));
    InMux I__8417 (
            .O(N__36235),
            .I(\b2v_inst11.mult1_un68_sum_cry_7 ));
    InMux I__8416 (
            .O(N__36232),
            .I(N__36227));
    CascadeMux I__8415 (
            .O(N__36231),
            .I(N__36223));
    InMux I__8414 (
            .O(N__36230),
            .I(N__36219));
    LocalMux I__8413 (
            .O(N__36227),
            .I(N__36216));
    InMux I__8412 (
            .O(N__36226),
            .I(N__36211));
    InMux I__8411 (
            .O(N__36223),
            .I(N__36211));
    InMux I__8410 (
            .O(N__36222),
            .I(N__36208));
    LocalMux I__8409 (
            .O(N__36219),
            .I(N__36205));
    Odrv12 I__8408 (
            .O(N__36216),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__8407 (
            .O(N__36211),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    LocalMux I__8406 (
            .O(N__36208),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    Odrv4 I__8405 (
            .O(N__36205),
            .I(\b2v_inst11.mult1_un68_sum_s_8 ));
    CascadeMux I__8404 (
            .O(N__36196),
            .I(N__36191));
    InMux I__8403 (
            .O(N__36195),
            .I(N__36188));
    InMux I__8402 (
            .O(N__36194),
            .I(N__36182));
    InMux I__8401 (
            .O(N__36191),
            .I(N__36182));
    LocalMux I__8400 (
            .O(N__36188),
            .I(N__36179));
    InMux I__8399 (
            .O(N__36187),
            .I(N__36176));
    LocalMux I__8398 (
            .O(N__36182),
            .I(N__36171));
    Span4Mux_s0_h I__8397 (
            .O(N__36179),
            .I(N__36171));
    LocalMux I__8396 (
            .O(N__36176),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    Odrv4 I__8395 (
            .O(N__36171),
            .I(\b2v_inst11.mult1_un54_sum_s_8 ));
    CascadeMux I__8394 (
            .O(N__36166),
            .I(N__36162));
    CascadeMux I__8393 (
            .O(N__36165),
            .I(N__36158));
    InMux I__8392 (
            .O(N__36162),
            .I(N__36151));
    InMux I__8391 (
            .O(N__36161),
            .I(N__36151));
    InMux I__8390 (
            .O(N__36158),
            .I(N__36151));
    LocalMux I__8389 (
            .O(N__36151),
            .I(\b2v_inst11.mult1_un54_sum_i_8 ));
    InMux I__8388 (
            .O(N__36148),
            .I(N__36141));
    InMux I__8387 (
            .O(N__36147),
            .I(N__36141));
    InMux I__8386 (
            .O(N__36146),
            .I(N__36138));
    LocalMux I__8385 (
            .O(N__36141),
            .I(\b2v_inst6.N_192 ));
    LocalMux I__8384 (
            .O(N__36138),
            .I(\b2v_inst6.N_192 ));
    CascadeMux I__8383 (
            .O(N__36133),
            .I(\b2v_inst6.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__8382 (
            .O(N__36130),
            .I(N__36125));
    SRMux I__8381 (
            .O(N__36129),
            .I(N__36121));
    SRMux I__8380 (
            .O(N__36128),
            .I(N__36115));
    InMux I__8379 (
            .O(N__36125),
            .I(N__36107));
    InMux I__8378 (
            .O(N__36124),
            .I(N__36107));
    LocalMux I__8377 (
            .O(N__36121),
            .I(N__36104));
    InMux I__8376 (
            .O(N__36120),
            .I(N__36099));
    SRMux I__8375 (
            .O(N__36119),
            .I(N__36099));
    SRMux I__8374 (
            .O(N__36118),
            .I(N__36096));
    LocalMux I__8373 (
            .O(N__36115),
            .I(N__36093));
    SRMux I__8372 (
            .O(N__36114),
            .I(N__36090));
    InMux I__8371 (
            .O(N__36113),
            .I(N__36077));
    InMux I__8370 (
            .O(N__36112),
            .I(N__36077));
    LocalMux I__8369 (
            .O(N__36107),
            .I(N__36067));
    Span4Mux_s1_v I__8368 (
            .O(N__36104),
            .I(N__36067));
    LocalMux I__8367 (
            .O(N__36099),
            .I(N__36067));
    LocalMux I__8366 (
            .O(N__36096),
            .I(N__36067));
    Span4Mux_v I__8365 (
            .O(N__36093),
            .I(N__36062));
    LocalMux I__8364 (
            .O(N__36090),
            .I(N__36062));
    InMux I__8363 (
            .O(N__36089),
            .I(N__36057));
    InMux I__8362 (
            .O(N__36088),
            .I(N__36057));
    InMux I__8361 (
            .O(N__36087),
            .I(N__36050));
    InMux I__8360 (
            .O(N__36086),
            .I(N__36050));
    InMux I__8359 (
            .O(N__36085),
            .I(N__36050));
    InMux I__8358 (
            .O(N__36084),
            .I(N__36043));
    InMux I__8357 (
            .O(N__36083),
            .I(N__36043));
    InMux I__8356 (
            .O(N__36082),
            .I(N__36043));
    LocalMux I__8355 (
            .O(N__36077),
            .I(N__36040));
    CascadeMux I__8354 (
            .O(N__36076),
            .I(N__36033));
    Span4Mux_v I__8353 (
            .O(N__36067),
            .I(N__36018));
    Span4Mux_v I__8352 (
            .O(N__36062),
            .I(N__36018));
    LocalMux I__8351 (
            .O(N__36057),
            .I(N__36009));
    LocalMux I__8350 (
            .O(N__36050),
            .I(N__36009));
    LocalMux I__8349 (
            .O(N__36043),
            .I(N__36009));
    Sp12to4 I__8348 (
            .O(N__36040),
            .I(N__36009));
    InMux I__8347 (
            .O(N__36039),
            .I(N__36004));
    InMux I__8346 (
            .O(N__36038),
            .I(N__36004));
    InMux I__8345 (
            .O(N__36037),
            .I(N__36001));
    SRMux I__8344 (
            .O(N__36036),
            .I(N__35996));
    InMux I__8343 (
            .O(N__36033),
            .I(N__35996));
    InMux I__8342 (
            .O(N__36032),
            .I(N__35991));
    InMux I__8341 (
            .O(N__36031),
            .I(N__35991));
    InMux I__8340 (
            .O(N__36030),
            .I(N__35984));
    InMux I__8339 (
            .O(N__36029),
            .I(N__35984));
    InMux I__8338 (
            .O(N__36028),
            .I(N__35984));
    InMux I__8337 (
            .O(N__36027),
            .I(N__35975));
    InMux I__8336 (
            .O(N__36026),
            .I(N__35975));
    InMux I__8335 (
            .O(N__36025),
            .I(N__35975));
    InMux I__8334 (
            .O(N__36024),
            .I(N__35975));
    InMux I__8333 (
            .O(N__36023),
            .I(N__35972));
    Span4Mux_v I__8332 (
            .O(N__36018),
            .I(N__35969));
    Span12Mux_s10_v I__8331 (
            .O(N__36009),
            .I(N__35966));
    LocalMux I__8330 (
            .O(N__36004),
            .I(N__35951));
    LocalMux I__8329 (
            .O(N__36001),
            .I(N__35951));
    LocalMux I__8328 (
            .O(N__35996),
            .I(N__35951));
    LocalMux I__8327 (
            .O(N__35991),
            .I(N__35951));
    LocalMux I__8326 (
            .O(N__35984),
            .I(N__35951));
    LocalMux I__8325 (
            .O(N__35975),
            .I(N__35951));
    LocalMux I__8324 (
            .O(N__35972),
            .I(N__35951));
    Odrv4 I__8323 (
            .O(N__35969),
            .I(\b2v_inst6.count_0_sqmuxa ));
    Odrv12 I__8322 (
            .O(N__35966),
            .I(\b2v_inst6.count_0_sqmuxa ));
    Odrv12 I__8321 (
            .O(N__35951),
            .I(\b2v_inst6.count_0_sqmuxa ));
    InMux I__8320 (
            .O(N__35944),
            .I(N__35941));
    LocalMux I__8319 (
            .O(N__35941),
            .I(\b2v_inst6.curr_state_1_0 ));
    CascadeMux I__8318 (
            .O(N__35938),
            .I(N__35935));
    InMux I__8317 (
            .O(N__35935),
            .I(N__35926));
    CascadeMux I__8316 (
            .O(N__35934),
            .I(N__35919));
    InMux I__8315 (
            .O(N__35933),
            .I(N__35910));
    InMux I__8314 (
            .O(N__35932),
            .I(N__35910));
    InMux I__8313 (
            .O(N__35931),
            .I(N__35905));
    InMux I__8312 (
            .O(N__35930),
            .I(N__35905));
    CascadeMux I__8311 (
            .O(N__35929),
            .I(N__35893));
    LocalMux I__8310 (
            .O(N__35926),
            .I(N__35888));
    InMux I__8309 (
            .O(N__35925),
            .I(N__35880));
    InMux I__8308 (
            .O(N__35924),
            .I(N__35880));
    InMux I__8307 (
            .O(N__35923),
            .I(N__35871));
    InMux I__8306 (
            .O(N__35922),
            .I(N__35871));
    InMux I__8305 (
            .O(N__35919),
            .I(N__35871));
    InMux I__8304 (
            .O(N__35918),
            .I(N__35871));
    InMux I__8303 (
            .O(N__35917),
            .I(N__35867));
    InMux I__8302 (
            .O(N__35916),
            .I(N__35862));
    InMux I__8301 (
            .O(N__35915),
            .I(N__35862));
    LocalMux I__8300 (
            .O(N__35910),
            .I(N__35854));
    LocalMux I__8299 (
            .O(N__35905),
            .I(N__35854));
    InMux I__8298 (
            .O(N__35904),
            .I(N__35847));
    InMux I__8297 (
            .O(N__35903),
            .I(N__35847));
    InMux I__8296 (
            .O(N__35902),
            .I(N__35847));
    InMux I__8295 (
            .O(N__35901),
            .I(N__35844));
    InMux I__8294 (
            .O(N__35900),
            .I(N__35837));
    InMux I__8293 (
            .O(N__35899),
            .I(N__35837));
    InMux I__8292 (
            .O(N__35898),
            .I(N__35837));
    InMux I__8291 (
            .O(N__35897),
            .I(N__35834));
    InMux I__8290 (
            .O(N__35896),
            .I(N__35831));
    InMux I__8289 (
            .O(N__35893),
            .I(N__35828));
    InMux I__8288 (
            .O(N__35892),
            .I(N__35821));
    InMux I__8287 (
            .O(N__35891),
            .I(N__35821));
    Span4Mux_v I__8286 (
            .O(N__35888),
            .I(N__35816));
    InMux I__8285 (
            .O(N__35887),
            .I(N__35807));
    InMux I__8284 (
            .O(N__35886),
            .I(N__35802));
    InMux I__8283 (
            .O(N__35885),
            .I(N__35802));
    LocalMux I__8282 (
            .O(N__35880),
            .I(N__35797));
    LocalMux I__8281 (
            .O(N__35871),
            .I(N__35797));
    InMux I__8280 (
            .O(N__35870),
            .I(N__35794));
    LocalMux I__8279 (
            .O(N__35867),
            .I(N__35789));
    LocalMux I__8278 (
            .O(N__35862),
            .I(N__35789));
    InMux I__8277 (
            .O(N__35861),
            .I(N__35782));
    InMux I__8276 (
            .O(N__35860),
            .I(N__35782));
    InMux I__8275 (
            .O(N__35859),
            .I(N__35782));
    Span12Mux_s9_h I__8274 (
            .O(N__35854),
            .I(N__35779));
    LocalMux I__8273 (
            .O(N__35847),
            .I(N__35776));
    LocalMux I__8272 (
            .O(N__35844),
            .I(N__35769));
    LocalMux I__8271 (
            .O(N__35837),
            .I(N__35769));
    LocalMux I__8270 (
            .O(N__35834),
            .I(N__35764));
    LocalMux I__8269 (
            .O(N__35831),
            .I(N__35764));
    LocalMux I__8268 (
            .O(N__35828),
            .I(N__35761));
    InMux I__8267 (
            .O(N__35827),
            .I(N__35758));
    InMux I__8266 (
            .O(N__35826),
            .I(N__35755));
    LocalMux I__8265 (
            .O(N__35821),
            .I(N__35752));
    InMux I__8264 (
            .O(N__35820),
            .I(N__35749));
    InMux I__8263 (
            .O(N__35819),
            .I(N__35746));
    Span4Mux_v I__8262 (
            .O(N__35816),
            .I(N__35741));
    InMux I__8261 (
            .O(N__35815),
            .I(N__35736));
    InMux I__8260 (
            .O(N__35814),
            .I(N__35736));
    InMux I__8259 (
            .O(N__35813),
            .I(N__35731));
    InMux I__8258 (
            .O(N__35812),
            .I(N__35731));
    InMux I__8257 (
            .O(N__35811),
            .I(N__35726));
    InMux I__8256 (
            .O(N__35810),
            .I(N__35726));
    LocalMux I__8255 (
            .O(N__35807),
            .I(N__35715));
    LocalMux I__8254 (
            .O(N__35802),
            .I(N__35715));
    Span4Mux_v I__8253 (
            .O(N__35797),
            .I(N__35715));
    LocalMux I__8252 (
            .O(N__35794),
            .I(N__35715));
    Span4Mux_s1_v I__8251 (
            .O(N__35789),
            .I(N__35715));
    LocalMux I__8250 (
            .O(N__35782),
            .I(N__35710));
    Span12Mux_v I__8249 (
            .O(N__35779),
            .I(N__35710));
    Span12Mux_s4_h I__8248 (
            .O(N__35776),
            .I(N__35707));
    InMux I__8247 (
            .O(N__35775),
            .I(N__35702));
    InMux I__8246 (
            .O(N__35774),
            .I(N__35702));
    Span12Mux_s7_h I__8245 (
            .O(N__35769),
            .I(N__35699));
    Span4Mux_v I__8244 (
            .O(N__35764),
            .I(N__35684));
    Span4Mux_h I__8243 (
            .O(N__35761),
            .I(N__35684));
    LocalMux I__8242 (
            .O(N__35758),
            .I(N__35684));
    LocalMux I__8241 (
            .O(N__35755),
            .I(N__35684));
    Span4Mux_h I__8240 (
            .O(N__35752),
            .I(N__35684));
    LocalMux I__8239 (
            .O(N__35749),
            .I(N__35684));
    LocalMux I__8238 (
            .O(N__35746),
            .I(N__35684));
    InMux I__8237 (
            .O(N__35745),
            .I(N__35679));
    InMux I__8236 (
            .O(N__35744),
            .I(N__35679));
    Odrv4 I__8235 (
            .O(N__35741),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__8234 (
            .O(N__35736),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__8233 (
            .O(N__35731),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__8232 (
            .O(N__35726),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__8231 (
            .O(N__35715),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv12 I__8230 (
            .O(N__35710),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv12 I__8229 (
            .O(N__35707),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__8228 (
            .O(N__35702),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv12 I__8227 (
            .O(N__35699),
            .I(SYNTHESIZED_WIRE_1keep_3));
    Odrv4 I__8226 (
            .O(N__35684),
            .I(SYNTHESIZED_WIRE_1keep_3));
    LocalMux I__8225 (
            .O(N__35679),
            .I(SYNTHESIZED_WIRE_1keep_3));
    InMux I__8224 (
            .O(N__35656),
            .I(N__35647));
    InMux I__8223 (
            .O(N__35655),
            .I(N__35647));
    InMux I__8222 (
            .O(N__35654),
            .I(N__35640));
    InMux I__8221 (
            .O(N__35653),
            .I(N__35640));
    InMux I__8220 (
            .O(N__35652),
            .I(N__35640));
    LocalMux I__8219 (
            .O(N__35647),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    LocalMux I__8218 (
            .O(N__35640),
            .I(\b2v_inst6.curr_stateZ0Z_0 ));
    CascadeMux I__8217 (
            .O(N__35635),
            .I(\b2v_inst6.curr_stateZ0Z_1_cascade_ ));
    InMux I__8216 (
            .O(N__35632),
            .I(N__35627));
    InMux I__8215 (
            .O(N__35631),
            .I(N__35622));
    InMux I__8214 (
            .O(N__35630),
            .I(N__35622));
    LocalMux I__8213 (
            .O(N__35627),
            .I(\b2v_inst6.curr_state_RNIUL1J2Z0Z_0 ));
    LocalMux I__8212 (
            .O(N__35622),
            .I(\b2v_inst6.curr_state_RNIUL1J2Z0Z_0 ));
    InMux I__8211 (
            .O(N__35617),
            .I(N__35614));
    LocalMux I__8210 (
            .O(N__35614),
            .I(\b2v_inst6.curr_state_7_0 ));
    InMux I__8209 (
            .O(N__35611),
            .I(\b2v_inst11.mult1_un75_sum_cry_5 ));
    CascadeMux I__8208 (
            .O(N__35608),
            .I(N__35604));
    CascadeMux I__8207 (
            .O(N__35607),
            .I(N__35600));
    InMux I__8206 (
            .O(N__35604),
            .I(N__35593));
    InMux I__8205 (
            .O(N__35603),
            .I(N__35593));
    InMux I__8204 (
            .O(N__35600),
            .I(N__35593));
    LocalMux I__8203 (
            .O(N__35593),
            .I(\b2v_inst11.mult1_un68_sum_i_0_8 ));
    CascadeMux I__8202 (
            .O(N__35590),
            .I(N__35587));
    InMux I__8201 (
            .O(N__35587),
            .I(N__35584));
    LocalMux I__8200 (
            .O(N__35584),
            .I(\b2v_inst11.mult1_un82_sum_axb_8 ));
    InMux I__8199 (
            .O(N__35581),
            .I(\b2v_inst11.mult1_un75_sum_cry_6 ));
    InMux I__8198 (
            .O(N__35578),
            .I(\b2v_inst11.mult1_un75_sum_cry_7 ));
    InMux I__8197 (
            .O(N__35575),
            .I(N__35571));
    CascadeMux I__8196 (
            .O(N__35574),
            .I(N__35567));
    LocalMux I__8195 (
            .O(N__35571),
            .I(N__35563));
    InMux I__8194 (
            .O(N__35570),
            .I(N__35558));
    InMux I__8193 (
            .O(N__35567),
            .I(N__35558));
    InMux I__8192 (
            .O(N__35566),
            .I(N__35555));
    Odrv12 I__8191 (
            .O(N__35563),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__8190 (
            .O(N__35558),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    LocalMux I__8189 (
            .O(N__35555),
            .I(\b2v_inst11.mult1_un75_sum_s_8 ));
    CascadeMux I__8188 (
            .O(N__35548),
            .I(\b2v_inst11.mult1_un75_sum_s_8_cascade_ ));
    CascadeMux I__8187 (
            .O(N__35545),
            .I(N__35541));
    CascadeMux I__8186 (
            .O(N__35544),
            .I(N__35537));
    InMux I__8185 (
            .O(N__35541),
            .I(N__35530));
    InMux I__8184 (
            .O(N__35540),
            .I(N__35530));
    InMux I__8183 (
            .O(N__35537),
            .I(N__35530));
    LocalMux I__8182 (
            .O(N__35530),
            .I(\b2v_inst11.mult1_un75_sum_i_0_8 ));
    InMux I__8181 (
            .O(N__35527),
            .I(N__35523));
    InMux I__8180 (
            .O(N__35526),
            .I(N__35520));
    LocalMux I__8179 (
            .O(N__35523),
            .I(N__35517));
    LocalMux I__8178 (
            .O(N__35520),
            .I(N__35514));
    Span4Mux_v I__8177 (
            .O(N__35517),
            .I(N__35511));
    Span4Mux_s2_h I__8176 (
            .O(N__35514),
            .I(N__35508));
    Odrv4 I__8175 (
            .O(N__35511),
            .I(\b2v_inst11.mult1_un68_sum ));
    Odrv4 I__8174 (
            .O(N__35508),
            .I(\b2v_inst11.mult1_un68_sum ));
    InMux I__8173 (
            .O(N__35503),
            .I(N__35500));
    LocalMux I__8172 (
            .O(N__35500),
            .I(\b2v_inst11.mult1_un61_sum_i ));
    CascadeMux I__8171 (
            .O(N__35497),
            .I(N__35494));
    InMux I__8170 (
            .O(N__35494),
            .I(N__35491));
    LocalMux I__8169 (
            .O(N__35491),
            .I(\b2v_inst11.mult1_un68_sum_cry_3_s ));
    InMux I__8168 (
            .O(N__35488),
            .I(\b2v_inst11.mult1_un68_sum_cry_2 ));
    CascadeMux I__8167 (
            .O(N__35485),
            .I(N__35482));
    InMux I__8166 (
            .O(N__35482),
            .I(N__35479));
    LocalMux I__8165 (
            .O(N__35479),
            .I(\b2v_inst11.mult1_un61_sum_cry_3_s ));
    InMux I__8164 (
            .O(N__35476),
            .I(N__35473));
    LocalMux I__8163 (
            .O(N__35473),
            .I(\b2v_inst11.mult1_un68_sum_cry_4_s ));
    InMux I__8162 (
            .O(N__35470),
            .I(\b2v_inst11.mult1_un68_sum_cry_3 ));
    InMux I__8161 (
            .O(N__35467),
            .I(N__35464));
    LocalMux I__8160 (
            .O(N__35464),
            .I(\b2v_inst11.mult1_un61_sum_cry_4_s ));
    CascadeMux I__8159 (
            .O(N__35461),
            .I(N__35458));
    InMux I__8158 (
            .O(N__35458),
            .I(N__35455));
    LocalMux I__8157 (
            .O(N__35455),
            .I(\b2v_inst11.mult1_un68_sum_cry_5_s ));
    InMux I__8156 (
            .O(N__35452),
            .I(\b2v_inst11.mult1_un68_sum_cry_4 ));
    CascadeMux I__8155 (
            .O(N__35449),
            .I(N__35444));
    InMux I__8154 (
            .O(N__35448),
            .I(N__35440));
    InMux I__8153 (
            .O(N__35447),
            .I(N__35435));
    InMux I__8152 (
            .O(N__35444),
            .I(N__35435));
    InMux I__8151 (
            .O(N__35443),
            .I(N__35432));
    LocalMux I__8150 (
            .O(N__35440),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__8149 (
            .O(N__35435),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    LocalMux I__8148 (
            .O(N__35432),
            .I(\b2v_inst11.mult1_un61_sum_s_8 ));
    CascadeMux I__8147 (
            .O(N__35425),
            .I(N__35422));
    InMux I__8146 (
            .O(N__35422),
            .I(N__35419));
    LocalMux I__8145 (
            .O(N__35419),
            .I(\b2v_inst11.mult1_un61_sum_cry_5_s ));
    InMux I__8144 (
            .O(N__35416),
            .I(N__35413));
    LocalMux I__8143 (
            .O(N__35413),
            .I(\b2v_inst11.mult1_un68_sum_cry_6_s ));
    InMux I__8142 (
            .O(N__35410),
            .I(N__35407));
    LocalMux I__8141 (
            .O(N__35407),
            .I(N__35404));
    Odrv4 I__8140 (
            .O(N__35404),
            .I(\b2v_inst11.mult1_un82_sum_cry_6_s ));
    InMux I__8139 (
            .O(N__35401),
            .I(\b2v_inst11.mult1_un82_sum_cry_5 ));
    CascadeMux I__8138 (
            .O(N__35398),
            .I(N__35395));
    InMux I__8137 (
            .O(N__35395),
            .I(N__35392));
    LocalMux I__8136 (
            .O(N__35392),
            .I(\b2v_inst11.mult1_un89_sum_axb_8 ));
    InMux I__8135 (
            .O(N__35389),
            .I(\b2v_inst11.mult1_un82_sum_cry_6 ));
    InMux I__8134 (
            .O(N__35386),
            .I(\b2v_inst11.mult1_un82_sum_cry_7 ));
    CascadeMux I__8133 (
            .O(N__35383),
            .I(N__35378));
    InMux I__8132 (
            .O(N__35382),
            .I(N__35374));
    InMux I__8131 (
            .O(N__35381),
            .I(N__35369));
    InMux I__8130 (
            .O(N__35378),
            .I(N__35369));
    InMux I__8129 (
            .O(N__35377),
            .I(N__35366));
    LocalMux I__8128 (
            .O(N__35374),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__8127 (
            .O(N__35369),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    LocalMux I__8126 (
            .O(N__35366),
            .I(\b2v_inst11.mult1_un82_sum_s_8 ));
    CascadeMux I__8125 (
            .O(N__35359),
            .I(\b2v_inst11.mult1_un82_sum_s_8_cascade_ ));
    CascadeMux I__8124 (
            .O(N__35356),
            .I(N__35352));
    CascadeMux I__8123 (
            .O(N__35355),
            .I(N__35348));
    InMux I__8122 (
            .O(N__35352),
            .I(N__35341));
    InMux I__8121 (
            .O(N__35351),
            .I(N__35341));
    InMux I__8120 (
            .O(N__35348),
            .I(N__35341));
    LocalMux I__8119 (
            .O(N__35341),
            .I(\b2v_inst11.mult1_un82_sum_i_0_8 ));
    InMux I__8118 (
            .O(N__35338),
            .I(N__35334));
    InMux I__8117 (
            .O(N__35337),
            .I(N__35331));
    LocalMux I__8116 (
            .O(N__35334),
            .I(N__35328));
    LocalMux I__8115 (
            .O(N__35331),
            .I(N__35323));
    Span4Mux_v I__8114 (
            .O(N__35328),
            .I(N__35323));
    Odrv4 I__8113 (
            .O(N__35323),
            .I(\b2v_inst11.mult1_un75_sum ));
    InMux I__8112 (
            .O(N__35320),
            .I(N__35317));
    LocalMux I__8111 (
            .O(N__35317),
            .I(\b2v_inst11.mult1_un68_sum_i ));
    CascadeMux I__8110 (
            .O(N__35314),
            .I(N__35311));
    InMux I__8109 (
            .O(N__35311),
            .I(N__35308));
    LocalMux I__8108 (
            .O(N__35308),
            .I(\b2v_inst11.mult1_un75_sum_cry_3_s ));
    InMux I__8107 (
            .O(N__35305),
            .I(\b2v_inst11.mult1_un75_sum_cry_2 ));
    InMux I__8106 (
            .O(N__35302),
            .I(N__35299));
    LocalMux I__8105 (
            .O(N__35299),
            .I(\b2v_inst11.mult1_un75_sum_cry_4_s ));
    InMux I__8104 (
            .O(N__35296),
            .I(\b2v_inst11.mult1_un75_sum_cry_3 ));
    CascadeMux I__8103 (
            .O(N__35293),
            .I(N__35290));
    InMux I__8102 (
            .O(N__35290),
            .I(N__35287));
    LocalMux I__8101 (
            .O(N__35287),
            .I(\b2v_inst11.mult1_un75_sum_cry_5_s ));
    InMux I__8100 (
            .O(N__35284),
            .I(\b2v_inst11.mult1_un75_sum_cry_4 ));
    InMux I__8099 (
            .O(N__35281),
            .I(N__35278));
    LocalMux I__8098 (
            .O(N__35278),
            .I(\b2v_inst11.mult1_un75_sum_cry_6_s ));
    InMux I__8097 (
            .O(N__35275),
            .I(N__35272));
    LocalMux I__8096 (
            .O(N__35272),
            .I(\b2v_inst11.mult1_un89_sum_cry_5_s ));
    InMux I__8095 (
            .O(N__35269),
            .I(N__35266));
    LocalMux I__8094 (
            .O(N__35266),
            .I(N__35263));
    Span4Mux_h I__8093 (
            .O(N__35263),
            .I(N__35260));
    Odrv4 I__8092 (
            .O(N__35260),
            .I(\b2v_inst11.mult1_un96_sum_cry_6_s ));
    InMux I__8091 (
            .O(N__35257),
            .I(\b2v_inst11.mult1_un96_sum_cry_5 ));
    InMux I__8090 (
            .O(N__35254),
            .I(N__35251));
    LocalMux I__8089 (
            .O(N__35251),
            .I(\b2v_inst11.mult1_un89_sum_cry_6_s ));
    CascadeMux I__8088 (
            .O(N__35248),
            .I(N__35245));
    InMux I__8087 (
            .O(N__35245),
            .I(N__35242));
    LocalMux I__8086 (
            .O(N__35242),
            .I(N__35239));
    Span4Mux_h I__8085 (
            .O(N__35239),
            .I(N__35236));
    Odrv4 I__8084 (
            .O(N__35236),
            .I(\b2v_inst11.mult1_un103_sum_axb_8 ));
    InMux I__8083 (
            .O(N__35233),
            .I(\b2v_inst11.mult1_un96_sum_cry_6 ));
    CascadeMux I__8082 (
            .O(N__35230),
            .I(N__35227));
    InMux I__8081 (
            .O(N__35227),
            .I(N__35224));
    LocalMux I__8080 (
            .O(N__35224),
            .I(\b2v_inst11.mult1_un96_sum_axb_8 ));
    InMux I__8079 (
            .O(N__35221),
            .I(\b2v_inst11.mult1_un96_sum_cry_7 ));
    CascadeMux I__8078 (
            .O(N__35218),
            .I(N__35214));
    InMux I__8077 (
            .O(N__35217),
            .I(N__35208));
    InMux I__8076 (
            .O(N__35214),
            .I(N__35208));
    InMux I__8075 (
            .O(N__35213),
            .I(N__35205));
    LocalMux I__8074 (
            .O(N__35208),
            .I(N__35198));
    LocalMux I__8073 (
            .O(N__35205),
            .I(N__35198));
    InMux I__8072 (
            .O(N__35204),
            .I(N__35195));
    InMux I__8071 (
            .O(N__35203),
            .I(N__35192));
    Span4Mux_h I__8070 (
            .O(N__35198),
            .I(N__35189));
    LocalMux I__8069 (
            .O(N__35195),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    LocalMux I__8068 (
            .O(N__35192),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    Odrv4 I__8067 (
            .O(N__35189),
            .I(\b2v_inst11.mult1_un96_sum_s_8 ));
    CascadeMux I__8066 (
            .O(N__35182),
            .I(N__35177));
    InMux I__8065 (
            .O(N__35181),
            .I(N__35172));
    InMux I__8064 (
            .O(N__35180),
            .I(N__35169));
    InMux I__8063 (
            .O(N__35177),
            .I(N__35162));
    InMux I__8062 (
            .O(N__35176),
            .I(N__35162));
    InMux I__8061 (
            .O(N__35175),
            .I(N__35162));
    LocalMux I__8060 (
            .O(N__35172),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__8059 (
            .O(N__35169),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    LocalMux I__8058 (
            .O(N__35162),
            .I(\b2v_inst11.mult1_un89_sum_s_8 ));
    CascadeMux I__8057 (
            .O(N__35155),
            .I(N__35151));
    CascadeMux I__8056 (
            .O(N__35154),
            .I(N__35147));
    InMux I__8055 (
            .O(N__35151),
            .I(N__35140));
    InMux I__8054 (
            .O(N__35150),
            .I(N__35140));
    InMux I__8053 (
            .O(N__35147),
            .I(N__35140));
    LocalMux I__8052 (
            .O(N__35140),
            .I(\b2v_inst11.mult1_un89_sum_i_0_8 ));
    InMux I__8051 (
            .O(N__35137),
            .I(N__35133));
    InMux I__8050 (
            .O(N__35136),
            .I(N__35130));
    LocalMux I__8049 (
            .O(N__35133),
            .I(N__35127));
    LocalMux I__8048 (
            .O(N__35130),
            .I(N__35124));
    Span4Mux_s3_h I__8047 (
            .O(N__35127),
            .I(N__35121));
    Odrv4 I__8046 (
            .O(N__35124),
            .I(\b2v_inst11.mult1_un82_sum ));
    Odrv4 I__8045 (
            .O(N__35121),
            .I(\b2v_inst11.mult1_un82_sum ));
    InMux I__8044 (
            .O(N__35116),
            .I(N__35113));
    LocalMux I__8043 (
            .O(N__35113),
            .I(\b2v_inst11.mult1_un75_sum_i ));
    CascadeMux I__8042 (
            .O(N__35110),
            .I(N__35107));
    InMux I__8041 (
            .O(N__35107),
            .I(N__35104));
    LocalMux I__8040 (
            .O(N__35104),
            .I(\b2v_inst11.mult1_un82_sum_cry_3_s ));
    InMux I__8039 (
            .O(N__35101),
            .I(\b2v_inst11.mult1_un82_sum_cry_2 ));
    InMux I__8038 (
            .O(N__35098),
            .I(N__35095));
    LocalMux I__8037 (
            .O(N__35095),
            .I(\b2v_inst11.mult1_un82_sum_cry_4_s ));
    InMux I__8036 (
            .O(N__35092),
            .I(\b2v_inst11.mult1_un82_sum_cry_3 ));
    CascadeMux I__8035 (
            .O(N__35089),
            .I(N__35086));
    InMux I__8034 (
            .O(N__35086),
            .I(N__35083));
    LocalMux I__8033 (
            .O(N__35083),
            .I(\b2v_inst11.mult1_un82_sum_cry_5_s ));
    InMux I__8032 (
            .O(N__35080),
            .I(\b2v_inst11.mult1_un82_sum_cry_4 ));
    InMux I__8031 (
            .O(N__35077),
            .I(N__35074));
    LocalMux I__8030 (
            .O(N__35074),
            .I(N__35071));
    Span4Mux_h I__8029 (
            .O(N__35071),
            .I(N__35068));
    Odrv4 I__8028 (
            .O(N__35068),
            .I(\b2v_inst11.mult1_un96_sum_i ));
    InMux I__8027 (
            .O(N__35065),
            .I(N__35062));
    LocalMux I__8026 (
            .O(N__35062),
            .I(\b2v_inst11.mult1_un68_sum_i_8 ));
    CEMux I__8025 (
            .O(N__35059),
            .I(N__35054));
    CEMux I__8024 (
            .O(N__35058),
            .I(N__35050));
    CascadeMux I__8023 (
            .O(N__35057),
            .I(N__35047));
    LocalMux I__8022 (
            .O(N__35054),
            .I(N__35035));
    CEMux I__8021 (
            .O(N__35053),
            .I(N__35032));
    LocalMux I__8020 (
            .O(N__35050),
            .I(N__35029));
    InMux I__8019 (
            .O(N__35047),
            .I(N__35024));
    CEMux I__8018 (
            .O(N__35046),
            .I(N__35024));
    InMux I__8017 (
            .O(N__35045),
            .I(N__35011));
    CEMux I__8016 (
            .O(N__35044),
            .I(N__35011));
    InMux I__8015 (
            .O(N__35043),
            .I(N__35008));
    InMux I__8014 (
            .O(N__35042),
            .I(N__35003));
    InMux I__8013 (
            .O(N__35041),
            .I(N__35003));
    InMux I__8012 (
            .O(N__35040),
            .I(N__34996));
    InMux I__8011 (
            .O(N__35039),
            .I(N__34996));
    InMux I__8010 (
            .O(N__35038),
            .I(N__34996));
    Span4Mux_s2_v I__8009 (
            .O(N__35035),
            .I(N__34990));
    LocalMux I__8008 (
            .O(N__35032),
            .I(N__34990));
    Span4Mux_s3_v I__8007 (
            .O(N__35029),
            .I(N__34987));
    LocalMux I__8006 (
            .O(N__35024),
            .I(N__34984));
    InMux I__8005 (
            .O(N__35023),
            .I(N__34981));
    InMux I__8004 (
            .O(N__35022),
            .I(N__34978));
    InMux I__8003 (
            .O(N__35021),
            .I(N__34971));
    InMux I__8002 (
            .O(N__35020),
            .I(N__34971));
    InMux I__8001 (
            .O(N__35019),
            .I(N__34971));
    CEMux I__8000 (
            .O(N__35018),
            .I(N__34964));
    InMux I__7999 (
            .O(N__35017),
            .I(N__34964));
    InMux I__7998 (
            .O(N__35016),
            .I(N__34964));
    LocalMux I__7997 (
            .O(N__35011),
            .I(N__34955));
    LocalMux I__7996 (
            .O(N__35008),
            .I(N__34955));
    LocalMux I__7995 (
            .O(N__35003),
            .I(N__34955));
    LocalMux I__7994 (
            .O(N__34996),
            .I(N__34955));
    CascadeMux I__7993 (
            .O(N__34995),
            .I(N__34952));
    Span4Mux_v I__7992 (
            .O(N__34990),
            .I(N__34949));
    Span4Mux_v I__7991 (
            .O(N__34987),
            .I(N__34944));
    Span4Mux_s0_h I__7990 (
            .O(N__34984),
            .I(N__34944));
    LocalMux I__7989 (
            .O(N__34981),
            .I(N__34933));
    LocalMux I__7988 (
            .O(N__34978),
            .I(N__34933));
    LocalMux I__7987 (
            .O(N__34971),
            .I(N__34933));
    LocalMux I__7986 (
            .O(N__34964),
            .I(N__34933));
    Sp12to4 I__7985 (
            .O(N__34955),
            .I(N__34933));
    InMux I__7984 (
            .O(N__34952),
            .I(N__34930));
    Odrv4 I__7983 (
            .O(N__34949),
            .I(\b2v_inst6.count_en ));
    Odrv4 I__7982 (
            .O(N__34944),
            .I(\b2v_inst6.count_en ));
    Odrv12 I__7981 (
            .O(N__34933),
            .I(\b2v_inst6.count_en ));
    LocalMux I__7980 (
            .O(N__34930),
            .I(\b2v_inst6.count_en ));
    InMux I__7979 (
            .O(N__34921),
            .I(N__34918));
    LocalMux I__7978 (
            .O(N__34918),
            .I(N__34915));
    Span4Mux_v I__7977 (
            .O(N__34915),
            .I(N__34912));
    Odrv4 I__7976 (
            .O(N__34912),
            .I(\b2v_inst6.count_RNIM2CM2Z0Z_0 ));
    CascadeMux I__7975 (
            .O(N__34909),
            .I(\b2v_inst6.count_en_cascade_ ));
    InMux I__7974 (
            .O(N__34906),
            .I(N__34903));
    LocalMux I__7973 (
            .O(N__34903),
            .I(\b2v_inst6.count_0_0 ));
    InMux I__7972 (
            .O(N__34900),
            .I(N__34896));
    CascadeMux I__7971 (
            .O(N__34899),
            .I(N__34893));
    LocalMux I__7970 (
            .O(N__34896),
            .I(N__34889));
    InMux I__7969 (
            .O(N__34893),
            .I(N__34884));
    InMux I__7968 (
            .O(N__34892),
            .I(N__34884));
    Span12Mux_s3_v I__7967 (
            .O(N__34889),
            .I(N__34879));
    LocalMux I__7966 (
            .O(N__34884),
            .I(N__34876));
    InMux I__7965 (
            .O(N__34883),
            .I(N__34871));
    InMux I__7964 (
            .O(N__34882),
            .I(N__34871));
    Odrv12 I__7963 (
            .O(N__34879),
            .I(\b2v_inst6.countZ0Z_0 ));
    Odrv4 I__7962 (
            .O(N__34876),
            .I(\b2v_inst6.countZ0Z_0 ));
    LocalMux I__7961 (
            .O(N__34871),
            .I(\b2v_inst6.countZ0Z_0 ));
    InMux I__7960 (
            .O(N__34864),
            .I(N__34860));
    InMux I__7959 (
            .O(N__34863),
            .I(N__34857));
    LocalMux I__7958 (
            .O(N__34860),
            .I(N__34854));
    LocalMux I__7957 (
            .O(N__34857),
            .I(N__34851));
    Span4Mux_s2_h I__7956 (
            .O(N__34854),
            .I(N__34848));
    Odrv12 I__7955 (
            .O(N__34851),
            .I(\b2v_inst11.mult1_un96_sum ));
    Odrv4 I__7954 (
            .O(N__34848),
            .I(\b2v_inst11.mult1_un96_sum ));
    InMux I__7953 (
            .O(N__34843),
            .I(N__34840));
    LocalMux I__7952 (
            .O(N__34840),
            .I(\b2v_inst11.mult1_un89_sum_i ));
    CascadeMux I__7951 (
            .O(N__34837),
            .I(N__34834));
    InMux I__7950 (
            .O(N__34834),
            .I(N__34831));
    LocalMux I__7949 (
            .O(N__34831),
            .I(N__34828));
    Span4Mux_h I__7948 (
            .O(N__34828),
            .I(N__34825));
    Odrv4 I__7947 (
            .O(N__34825),
            .I(\b2v_inst11.mult1_un96_sum_cry_3_s ));
    InMux I__7946 (
            .O(N__34822),
            .I(\b2v_inst11.mult1_un96_sum_cry_2 ));
    CascadeMux I__7945 (
            .O(N__34819),
            .I(N__34816));
    InMux I__7944 (
            .O(N__34816),
            .I(N__34813));
    LocalMux I__7943 (
            .O(N__34813),
            .I(\b2v_inst11.mult1_un89_sum_cry_3_s ));
    InMux I__7942 (
            .O(N__34810),
            .I(N__34807));
    LocalMux I__7941 (
            .O(N__34807),
            .I(N__34804));
    Span4Mux_v I__7940 (
            .O(N__34804),
            .I(N__34801));
    Odrv4 I__7939 (
            .O(N__34801),
            .I(\b2v_inst11.mult1_un96_sum_cry_4_s ));
    InMux I__7938 (
            .O(N__34798),
            .I(\b2v_inst11.mult1_un96_sum_cry_3 ));
    CascadeMux I__7937 (
            .O(N__34795),
            .I(N__34792));
    InMux I__7936 (
            .O(N__34792),
            .I(N__34789));
    LocalMux I__7935 (
            .O(N__34789),
            .I(\b2v_inst11.mult1_un89_sum_cry_4_s ));
    CascadeMux I__7934 (
            .O(N__34786),
            .I(N__34783));
    InMux I__7933 (
            .O(N__34783),
            .I(N__34780));
    LocalMux I__7932 (
            .O(N__34780),
            .I(N__34777));
    Span4Mux_v I__7931 (
            .O(N__34777),
            .I(N__34774));
    Odrv4 I__7930 (
            .O(N__34774),
            .I(\b2v_inst11.mult1_un96_sum_cry_5_s ));
    InMux I__7929 (
            .O(N__34771),
            .I(\b2v_inst11.mult1_un96_sum_cry_4 ));
    CascadeMux I__7928 (
            .O(N__34768),
            .I(\b2v_inst6.un2_count_1_axb_1_cascade_ ));
    InMux I__7927 (
            .O(N__34765),
            .I(N__34762));
    LocalMux I__7926 (
            .O(N__34762),
            .I(N__34759));
    IoSpan4Mux I__7925 (
            .O(N__34759),
            .I(N__34756));
    Odrv4 I__7924 (
            .O(N__34756),
            .I(V1P8A_OK_c));
    InMux I__7923 (
            .O(N__34753),
            .I(N__34750));
    LocalMux I__7922 (
            .O(N__34750),
            .I(N__34747));
    Span4Mux_v I__7921 (
            .O(N__34747),
            .I(N__34744));
    Span4Mux_v I__7920 (
            .O(N__34744),
            .I(N__34741));
    Odrv4 I__7919 (
            .O(N__34741),
            .I(V33A_OK_c));
    CascadeMux I__7918 (
            .O(N__34738),
            .I(N__34735));
    InMux I__7917 (
            .O(N__34735),
            .I(N__34732));
    LocalMux I__7916 (
            .O(N__34732),
            .I(V5A_OK_c));
    InMux I__7915 (
            .O(N__34729),
            .I(N__34726));
    LocalMux I__7914 (
            .O(N__34726),
            .I(VCCST_CPU_OK_c));
    CascadeMux I__7913 (
            .O(N__34723),
            .I(N__34718));
    CascadeMux I__7912 (
            .O(N__34722),
            .I(N__34713));
    InMux I__7911 (
            .O(N__34721),
            .I(N__34702));
    InMux I__7910 (
            .O(N__34718),
            .I(N__34702));
    InMux I__7909 (
            .O(N__34717),
            .I(N__34702));
    InMux I__7908 (
            .O(N__34716),
            .I(N__34702));
    InMux I__7907 (
            .O(N__34713),
            .I(N__34697));
    InMux I__7906 (
            .O(N__34712),
            .I(N__34697));
    InMux I__7905 (
            .O(N__34711),
            .I(N__34694));
    LocalMux I__7904 (
            .O(N__34702),
            .I(N__34689));
    LocalMux I__7903 (
            .O(N__34697),
            .I(N__34689));
    LocalMux I__7902 (
            .O(N__34694),
            .I(N__34686));
    Span12Mux_s8_v I__7901 (
            .O(N__34689),
            .I(N__34683));
    Span4Mux_v I__7900 (
            .O(N__34686),
            .I(N__34680));
    Odrv12 I__7899 (
            .O(N__34683),
            .I(N_1661));
    Odrv4 I__7898 (
            .O(N__34680),
            .I(N_1661));
    InMux I__7897 (
            .O(N__34675),
            .I(N__34669));
    InMux I__7896 (
            .O(N__34674),
            .I(N__34669));
    LocalMux I__7895 (
            .O(N__34669),
            .I(\b2v_inst6.count_0_1 ));
    CascadeMux I__7894 (
            .O(N__34666),
            .I(N__34663));
    InMux I__7893 (
            .O(N__34663),
            .I(N__34654));
    InMux I__7892 (
            .O(N__34662),
            .I(N__34654));
    InMux I__7891 (
            .O(N__34661),
            .I(N__34654));
    LocalMux I__7890 (
            .O(N__34654),
            .I(\b2v_inst6.count_RNI_0_1 ));
    InMux I__7889 (
            .O(N__34651),
            .I(N__34648));
    LocalMux I__7888 (
            .O(N__34648),
            .I(N__34645));
    Span4Mux_s3_v I__7887 (
            .O(N__34645),
            .I(N__34641));
    InMux I__7886 (
            .O(N__34644),
            .I(N__34638));
    Span4Mux_s0_h I__7885 (
            .O(N__34641),
            .I(N__34633));
    LocalMux I__7884 (
            .O(N__34638),
            .I(N__34633));
    Odrv4 I__7883 (
            .O(N__34633),
            .I(\b2v_inst6.countZ0Z_15 ));
    CascadeMux I__7882 (
            .O(N__34630),
            .I(\b2v_inst6.countZ0Z_1_cascade_ ));
    InMux I__7881 (
            .O(N__34627),
            .I(N__34621));
    InMux I__7880 (
            .O(N__34626),
            .I(N__34618));
    InMux I__7879 (
            .O(N__34625),
            .I(N__34615));
    InMux I__7878 (
            .O(N__34624),
            .I(N__34612));
    LocalMux I__7877 (
            .O(N__34621),
            .I(N__34607));
    LocalMux I__7876 (
            .O(N__34618),
            .I(N__34607));
    LocalMux I__7875 (
            .O(N__34615),
            .I(\b2v_inst6.countZ0Z_11 ));
    LocalMux I__7874 (
            .O(N__34612),
            .I(\b2v_inst6.countZ0Z_11 ));
    Odrv12 I__7873 (
            .O(N__34607),
            .I(\b2v_inst6.countZ0Z_11 ));
    InMux I__7872 (
            .O(N__34600),
            .I(N__34597));
    LocalMux I__7871 (
            .O(N__34597),
            .I(N__34594));
    Span4Mux_v I__7870 (
            .O(N__34594),
            .I(N__34591));
    Odrv4 I__7869 (
            .O(N__34591),
            .I(\b2v_inst6.count_1_i_a3_8_0 ));
    InMux I__7868 (
            .O(N__34588),
            .I(N__34585));
    LocalMux I__7867 (
            .O(N__34585),
            .I(N__34582));
    Odrv12 I__7866 (
            .O(N__34582),
            .I(\b2v_inst6.count_1_i_a3_9_0 ));
    CascadeMux I__7865 (
            .O(N__34579),
            .I(\b2v_inst6.count_1_i_a3_7_0_cascade_ ));
    InMux I__7864 (
            .O(N__34576),
            .I(N__34573));
    LocalMux I__7863 (
            .O(N__34573),
            .I(N__34570));
    Span4Mux_v I__7862 (
            .O(N__34570),
            .I(N__34567));
    Odrv4 I__7861 (
            .O(N__34567),
            .I(\b2v_inst6.count_1_i_a3_10_0 ));
    InMux I__7860 (
            .O(N__34564),
            .I(N__34558));
    InMux I__7859 (
            .O(N__34563),
            .I(N__34558));
    LocalMux I__7858 (
            .O(N__34558),
            .I(\b2v_inst6.N_389 ));
    CascadeMux I__7857 (
            .O(N__34555),
            .I(\b2v_inst6.N_389_cascade_ ));
    InMux I__7856 (
            .O(N__34552),
            .I(N__34549));
    LocalMux I__7855 (
            .O(N__34549),
            .I(\b2v_inst11.mult1_un75_sum_i_8 ));
    InMux I__7854 (
            .O(N__34546),
            .I(N__34543));
    LocalMux I__7853 (
            .O(N__34543),
            .I(\b2v_inst11.mult1_un96_sum_i_8 ));
    CascadeMux I__7852 (
            .O(N__34540),
            .I(\b2v_inst6.count_rst_11_cascade_ ));
    CascadeMux I__7851 (
            .O(N__34537),
            .I(N__34532));
    InMux I__7850 (
            .O(N__34536),
            .I(N__34529));
    InMux I__7849 (
            .O(N__34535),
            .I(N__34526));
    InMux I__7848 (
            .O(N__34532),
            .I(N__34523));
    LocalMux I__7847 (
            .O(N__34529),
            .I(N__34518));
    LocalMux I__7846 (
            .O(N__34526),
            .I(N__34518));
    LocalMux I__7845 (
            .O(N__34523),
            .I(\b2v_inst6.countZ0Z_3 ));
    Odrv12 I__7844 (
            .O(N__34518),
            .I(\b2v_inst6.countZ0Z_3 ));
    InMux I__7843 (
            .O(N__34513),
            .I(N__34507));
    InMux I__7842 (
            .O(N__34512),
            .I(N__34507));
    LocalMux I__7841 (
            .O(N__34507),
            .I(N__34504));
    Odrv12 I__7840 (
            .O(N__34504),
            .I(\b2v_inst6.un2_count_1_cry_2_THRU_CO ));
    CascadeMux I__7839 (
            .O(N__34501),
            .I(\b2v_inst6.countZ0Z_3_cascade_ ));
    InMux I__7838 (
            .O(N__34498),
            .I(N__34495));
    LocalMux I__7837 (
            .O(N__34495),
            .I(\b2v_inst6.count_0_3 ));
    CascadeMux I__7836 (
            .O(N__34492),
            .I(N__34489));
    InMux I__7835 (
            .O(N__34489),
            .I(N__34485));
    InMux I__7834 (
            .O(N__34488),
            .I(N__34482));
    LocalMux I__7833 (
            .O(N__34485),
            .I(N__34477));
    LocalMux I__7832 (
            .O(N__34482),
            .I(N__34477));
    Span4Mux_v I__7831 (
            .O(N__34477),
            .I(N__34474));
    Odrv4 I__7830 (
            .O(N__34474),
            .I(\b2v_inst6.un2_count_1_cry_10_THRU_CO ));
    CascadeMux I__7829 (
            .O(N__34471),
            .I(\b2v_inst6.N_394_cascade_ ));
    InMux I__7828 (
            .O(N__34468),
            .I(N__34465));
    LocalMux I__7827 (
            .O(N__34465),
            .I(\b2v_inst6.count_0_11 ));
    CascadeMux I__7826 (
            .O(N__34462),
            .I(\b2v_inst6.count_rst_3_cascade_ ));
    CascadeMux I__7825 (
            .O(N__34459),
            .I(N__34456));
    InMux I__7824 (
            .O(N__34456),
            .I(N__34453));
    LocalMux I__7823 (
            .O(N__34453),
            .I(N__34450));
    Span4Mux_s3_v I__7822 (
            .O(N__34450),
            .I(N__34447));
    Odrv4 I__7821 (
            .O(N__34447),
            .I(\b2v_inst6.un2_count_1_axb_1 ));
    InMux I__7820 (
            .O(N__34444),
            .I(N__34441));
    LocalMux I__7819 (
            .O(N__34441),
            .I(\b2v_inst6.count_0_10 ));
    InMux I__7818 (
            .O(N__34438),
            .I(N__34434));
    InMux I__7817 (
            .O(N__34437),
            .I(N__34431));
    LocalMux I__7816 (
            .O(N__34434),
            .I(N__34426));
    LocalMux I__7815 (
            .O(N__34431),
            .I(N__34426));
    Odrv12 I__7814 (
            .O(N__34426),
            .I(\b2v_inst6.un2_count_1_cry_6_THRU_CO ));
    InMux I__7813 (
            .O(N__34423),
            .I(N__34420));
    LocalMux I__7812 (
            .O(N__34420),
            .I(N__34417));
    Odrv4 I__7811 (
            .O(N__34417),
            .I(\b2v_inst6.count_0_7 ));
    CascadeMux I__7810 (
            .O(N__34414),
            .I(\b2v_inst6.count_rst_7_cascade_ ));
    InMux I__7809 (
            .O(N__34411),
            .I(N__34403));
    InMux I__7808 (
            .O(N__34410),
            .I(N__34403));
    InMux I__7807 (
            .O(N__34409),
            .I(N__34400));
    InMux I__7806 (
            .O(N__34408),
            .I(N__34397));
    LocalMux I__7805 (
            .O(N__34403),
            .I(N__34392));
    LocalMux I__7804 (
            .O(N__34400),
            .I(N__34392));
    LocalMux I__7803 (
            .O(N__34397),
            .I(\b2v_inst6.countZ0Z_7 ));
    Odrv12 I__7802 (
            .O(N__34392),
            .I(\b2v_inst6.countZ0Z_7 ));
    InMux I__7801 (
            .O(N__34387),
            .I(N__34381));
    InMux I__7800 (
            .O(N__34386),
            .I(N__34381));
    LocalMux I__7799 (
            .O(N__34381),
            .I(N__34378));
    Odrv4 I__7798 (
            .O(N__34378),
            .I(\b2v_inst6.count_rst ));
    InMux I__7797 (
            .O(N__34375),
            .I(N__34372));
    LocalMux I__7796 (
            .O(N__34372),
            .I(\b2v_inst6.count_0_15 ));
    InMux I__7795 (
            .O(N__34369),
            .I(N__34366));
    LocalMux I__7794 (
            .O(N__34366),
            .I(N__34363));
    Span4Mux_v I__7793 (
            .O(N__34363),
            .I(N__34359));
    InMux I__7792 (
            .O(N__34362),
            .I(N__34356));
    Odrv4 I__7791 (
            .O(N__34359),
            .I(\b2v_inst6.count_rst_12 ));
    LocalMux I__7790 (
            .O(N__34356),
            .I(\b2v_inst6.count_rst_12 ));
    InMux I__7789 (
            .O(N__34351),
            .I(N__34348));
    LocalMux I__7788 (
            .O(N__34348),
            .I(N__34345));
    Span4Mux_s1_v I__7787 (
            .O(N__34345),
            .I(N__34342));
    Odrv4 I__7786 (
            .O(N__34342),
            .I(\b2v_inst6.count_0_2 ));
    InMux I__7785 (
            .O(N__34339),
            .I(N__34336));
    LocalMux I__7784 (
            .O(N__34336),
            .I(\b2v_inst6.count_rst_6 ));
    InMux I__7783 (
            .O(N__34333),
            .I(N__34328));
    CascadeMux I__7782 (
            .O(N__34332),
            .I(N__34325));
    InMux I__7781 (
            .O(N__34331),
            .I(N__34322));
    LocalMux I__7780 (
            .O(N__34328),
            .I(N__34319));
    InMux I__7779 (
            .O(N__34325),
            .I(N__34316));
    LocalMux I__7778 (
            .O(N__34322),
            .I(N__34311));
    Span4Mux_s1_v I__7777 (
            .O(N__34319),
            .I(N__34311));
    LocalMux I__7776 (
            .O(N__34316),
            .I(\b2v_inst6.countZ0Z_8 ));
    Odrv4 I__7775 (
            .O(N__34311),
            .I(\b2v_inst6.countZ0Z_8 ));
    CascadeMux I__7774 (
            .O(N__34306),
            .I(\b2v_inst6.countZ0Z_8_cascade_ ));
    InMux I__7773 (
            .O(N__34303),
            .I(N__34299));
    InMux I__7772 (
            .O(N__34302),
            .I(N__34296));
    LocalMux I__7771 (
            .O(N__34299),
            .I(N__34291));
    LocalMux I__7770 (
            .O(N__34296),
            .I(N__34291));
    Span4Mux_v I__7769 (
            .O(N__34291),
            .I(N__34288));
    Odrv4 I__7768 (
            .O(N__34288),
            .I(\b2v_inst6.un2_count_1_cry_7_THRU_CO ));
    InMux I__7767 (
            .O(N__34285),
            .I(N__34282));
    LocalMux I__7766 (
            .O(N__34282),
            .I(\b2v_inst6.count_0_8 ));
    InMux I__7765 (
            .O(N__34279),
            .I(N__34276));
    LocalMux I__7764 (
            .O(N__34276),
            .I(N__34273));
    Odrv12 I__7763 (
            .O(N__34273),
            .I(\b2v_inst6.countZ0Z_10 ));
    CascadeMux I__7762 (
            .O(N__34270),
            .I(\b2v_inst6.countZ0Z_10_cascade_ ));
    InMux I__7761 (
            .O(N__34267),
            .I(N__34264));
    LocalMux I__7760 (
            .O(N__34264),
            .I(\b2v_inst6.count_0_12 ));
    InMux I__7759 (
            .O(N__34261),
            .I(N__34255));
    InMux I__7758 (
            .O(N__34260),
            .I(N__34255));
    LocalMux I__7757 (
            .O(N__34255),
            .I(N__34252));
    Odrv4 I__7756 (
            .O(N__34252),
            .I(\b2v_inst6.count_rst_2 ));
    CascadeMux I__7755 (
            .O(N__34249),
            .I(N__34246));
    InMux I__7754 (
            .O(N__34246),
            .I(N__34242));
    InMux I__7753 (
            .O(N__34245),
            .I(N__34239));
    LocalMux I__7752 (
            .O(N__34242),
            .I(N__34236));
    LocalMux I__7751 (
            .O(N__34239),
            .I(\b2v_inst6.countZ0Z_12 ));
    Odrv4 I__7750 (
            .O(N__34236),
            .I(\b2v_inst6.countZ0Z_12 ));
    CascadeMux I__7749 (
            .O(N__34231),
            .I(\b2v_inst6.count_rst_10_cascade_ ));
    CascadeMux I__7748 (
            .O(N__34228),
            .I(N__34224));
    InMux I__7747 (
            .O(N__34227),
            .I(N__34220));
    InMux I__7746 (
            .O(N__34224),
            .I(N__34217));
    InMux I__7745 (
            .O(N__34223),
            .I(N__34214));
    LocalMux I__7744 (
            .O(N__34220),
            .I(N__34211));
    LocalMux I__7743 (
            .O(N__34217),
            .I(\b2v_inst6.countZ0Z_4 ));
    LocalMux I__7742 (
            .O(N__34214),
            .I(\b2v_inst6.countZ0Z_4 ));
    Odrv12 I__7741 (
            .O(N__34211),
            .I(\b2v_inst6.countZ0Z_4 ));
    InMux I__7740 (
            .O(N__34204),
            .I(N__34198));
    InMux I__7739 (
            .O(N__34203),
            .I(N__34198));
    LocalMux I__7738 (
            .O(N__34198),
            .I(N__34195));
    Odrv12 I__7737 (
            .O(N__34195),
            .I(\b2v_inst6.un2_count_1_cry_3_THRU_CO ));
    CascadeMux I__7736 (
            .O(N__34192),
            .I(\b2v_inst6.countZ0Z_4_cascade_ ));
    InMux I__7735 (
            .O(N__34189),
            .I(N__34186));
    LocalMux I__7734 (
            .O(N__34186),
            .I(\b2v_inst6.count_0_4 ));
    InMux I__7733 (
            .O(N__34183),
            .I(N__34177));
    InMux I__7732 (
            .O(N__34182),
            .I(N__34177));
    LocalMux I__7731 (
            .O(N__34177),
            .I(N__34174));
    Odrv4 I__7730 (
            .O(N__34174),
            .I(\b2v_inst6.count_rst_4 ));
    InMux I__7729 (
            .O(N__34171),
            .I(\b2v_inst6.un2_count_1_cry_14 ));
    InMux I__7728 (
            .O(N__34168),
            .I(N__34165));
    LocalMux I__7727 (
            .O(N__34165),
            .I(N__34162));
    Odrv4 I__7726 (
            .O(N__34162),
            .I(\b2v_inst6.count_0_13 ));
    InMux I__7725 (
            .O(N__34159),
            .I(N__34155));
    InMux I__7724 (
            .O(N__34158),
            .I(N__34152));
    LocalMux I__7723 (
            .O(N__34155),
            .I(\b2v_inst6.count_rst_1 ));
    LocalMux I__7722 (
            .O(N__34152),
            .I(\b2v_inst6.count_rst_1 ));
    InMux I__7721 (
            .O(N__34147),
            .I(N__34144));
    LocalMux I__7720 (
            .O(N__34144),
            .I(N__34140));
    InMux I__7719 (
            .O(N__34143),
            .I(N__34137));
    Odrv4 I__7718 (
            .O(N__34140),
            .I(\b2v_inst6.countZ0Z_13 ));
    LocalMux I__7717 (
            .O(N__34137),
            .I(\b2v_inst6.countZ0Z_13 ));
    InMux I__7716 (
            .O(N__34132),
            .I(N__34129));
    LocalMux I__7715 (
            .O(N__34129),
            .I(\b2v_inst6.count_0_5 ));
    InMux I__7714 (
            .O(N__34126),
            .I(N__34120));
    InMux I__7713 (
            .O(N__34125),
            .I(N__34120));
    LocalMux I__7712 (
            .O(N__34120),
            .I(N__34117));
    Odrv12 I__7711 (
            .O(N__34117),
            .I(\b2v_inst6.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__7710 (
            .O(N__34114),
            .I(\b2v_inst6.countZ0Z_5_cascade_ ));
    InMux I__7709 (
            .O(N__34111),
            .I(N__34108));
    LocalMux I__7708 (
            .O(N__34108),
            .I(\b2v_inst6.count_rst_9 ));
    InMux I__7707 (
            .O(N__34105),
            .I(N__34102));
    LocalMux I__7706 (
            .O(N__34102),
            .I(\b2v_inst6.count_rst_5 ));
    CascadeMux I__7705 (
            .O(N__34099),
            .I(\b2v_inst6.countZ0Z_9_cascade_ ));
    InMux I__7704 (
            .O(N__34096),
            .I(N__34091));
    InMux I__7703 (
            .O(N__34095),
            .I(N__34086));
    InMux I__7702 (
            .O(N__34094),
            .I(N__34086));
    LocalMux I__7701 (
            .O(N__34091),
            .I(N__34083));
    LocalMux I__7700 (
            .O(N__34086),
            .I(\b2v_inst6.countZ0Z_5 ));
    Odrv4 I__7699 (
            .O(N__34083),
            .I(\b2v_inst6.countZ0Z_5 ));
    CascadeMux I__7698 (
            .O(N__34078),
            .I(N__34075));
    InMux I__7697 (
            .O(N__34075),
            .I(N__34068));
    InMux I__7696 (
            .O(N__34074),
            .I(N__34068));
    InMux I__7695 (
            .O(N__34073),
            .I(N__34065));
    LocalMux I__7694 (
            .O(N__34068),
            .I(\b2v_inst6.countZ0Z_9 ));
    LocalMux I__7693 (
            .O(N__34065),
            .I(\b2v_inst6.countZ0Z_9 ));
    InMux I__7692 (
            .O(N__34060),
            .I(N__34054));
    InMux I__7691 (
            .O(N__34059),
            .I(N__34054));
    LocalMux I__7690 (
            .O(N__34054),
            .I(\b2v_inst6.un2_count_1_cry_8_THRU_CO ));
    InMux I__7689 (
            .O(N__34051),
            .I(N__34048));
    LocalMux I__7688 (
            .O(N__34048),
            .I(\b2v_inst6.count_0_9 ));
    CascadeMux I__7687 (
            .O(N__34045),
            .I(N__34041));
    InMux I__7686 (
            .O(N__34044),
            .I(N__34038));
    InMux I__7685 (
            .O(N__34041),
            .I(N__34035));
    LocalMux I__7684 (
            .O(N__34038),
            .I(\b2v_inst6.countZ0Z_6 ));
    LocalMux I__7683 (
            .O(N__34035),
            .I(\b2v_inst6.countZ0Z_6 ));
    InMux I__7682 (
            .O(N__34030),
            .I(N__34024));
    InMux I__7681 (
            .O(N__34029),
            .I(N__34024));
    LocalMux I__7680 (
            .O(N__34024),
            .I(\b2v_inst6.count_rst_8 ));
    InMux I__7679 (
            .O(N__34021),
            .I(\b2v_inst6.un2_count_1_cry_5 ));
    InMux I__7678 (
            .O(N__34018),
            .I(\b2v_inst6.un2_count_1_cry_6 ));
    InMux I__7677 (
            .O(N__34015),
            .I(\b2v_inst6.un2_count_1_cry_7 ));
    InMux I__7676 (
            .O(N__34012),
            .I(bfn_12_2_0_));
    InMux I__7675 (
            .O(N__34009),
            .I(\b2v_inst6.un2_count_1_cry_9 ));
    InMux I__7674 (
            .O(N__34006),
            .I(\b2v_inst6.un2_count_1_cry_10 ));
    InMux I__7673 (
            .O(N__34003),
            .I(\b2v_inst6.un2_count_1_cry_11 ));
    InMux I__7672 (
            .O(N__34000),
            .I(\b2v_inst6.un2_count_1_cry_12 ));
    InMux I__7671 (
            .O(N__33997),
            .I(N__33994));
    LocalMux I__7670 (
            .O(N__33994),
            .I(\b2v_inst6.countZ0Z_14 ));
    InMux I__7669 (
            .O(N__33991),
            .I(N__33985));
    InMux I__7668 (
            .O(N__33990),
            .I(N__33985));
    LocalMux I__7667 (
            .O(N__33985),
            .I(\b2v_inst6.count_rst_0 ));
    InMux I__7666 (
            .O(N__33982),
            .I(\b2v_inst6.un2_count_1_cry_13 ));
    InMux I__7665 (
            .O(N__33979),
            .I(N__33976));
    LocalMux I__7664 (
            .O(N__33976),
            .I(N__33973));
    Odrv4 I__7663 (
            .O(N__33973),
            .I(\b2v_inst11.mult1_un159_sum_cry_4_s ));
    InMux I__7662 (
            .O(N__33970),
            .I(N__33967));
    LocalMux I__7661 (
            .O(N__33967),
            .I(N__33962));
    CascadeMux I__7660 (
            .O(N__33966),
            .I(N__33959));
    CascadeMux I__7659 (
            .O(N__33965),
            .I(N__33956));
    Span4Mux_v I__7658 (
            .O(N__33962),
            .I(N__33951));
    InMux I__7657 (
            .O(N__33959),
            .I(N__33948));
    InMux I__7656 (
            .O(N__33956),
            .I(N__33943));
    InMux I__7655 (
            .O(N__33955),
            .I(N__33943));
    InMux I__7654 (
            .O(N__33954),
            .I(N__33940));
    Span4Mux_v I__7653 (
            .O(N__33951),
            .I(N__33931));
    LocalMux I__7652 (
            .O(N__33948),
            .I(N__33931));
    LocalMux I__7651 (
            .O(N__33943),
            .I(N__33931));
    LocalMux I__7650 (
            .O(N__33940),
            .I(N__33931));
    Odrv4 I__7649 (
            .O(N__33931),
            .I(\b2v_inst11.mult1_un159_sum_s_7 ));
    InMux I__7648 (
            .O(N__33928),
            .I(N__33925));
    LocalMux I__7647 (
            .O(N__33925),
            .I(N__33922));
    Odrv4 I__7646 (
            .O(N__33922),
            .I(\b2v_inst11.mult1_un159_sum_cry_5_s ));
    CascadeMux I__7645 (
            .O(N__33919),
            .I(N__33915));
    CascadeMux I__7644 (
            .O(N__33918),
            .I(N__33911));
    InMux I__7643 (
            .O(N__33915),
            .I(N__33904));
    InMux I__7642 (
            .O(N__33914),
            .I(N__33904));
    InMux I__7641 (
            .O(N__33911),
            .I(N__33904));
    LocalMux I__7640 (
            .O(N__33904),
            .I(G_2836));
    InMux I__7639 (
            .O(N__33901),
            .I(N__33898));
    LocalMux I__7638 (
            .O(N__33898),
            .I(N__33895));
    Odrv12 I__7637 (
            .O(N__33895),
            .I(\b2v_inst11.mult1_un166_sum_axb_6 ));
    InMux I__7636 (
            .O(N__33892),
            .I(\b2v_inst11.mult1_un166_sum_cry_5 ));
    CascadeMux I__7635 (
            .O(N__33889),
            .I(N__33886));
    InMux I__7634 (
            .O(N__33886),
            .I(N__33883));
    LocalMux I__7633 (
            .O(N__33883),
            .I(N__33880));
    Span4Mux_v I__7632 (
            .O(N__33880),
            .I(N__33877));
    Span4Mux_v I__7631 (
            .O(N__33877),
            .I(N__33874));
    Odrv4 I__7630 (
            .O(N__33874),
            .I(\b2v_inst11.un85_clk_100khz_0 ));
    InMux I__7629 (
            .O(N__33871),
            .I(N__33867));
    InMux I__7628 (
            .O(N__33870),
            .I(N__33864));
    LocalMux I__7627 (
            .O(N__33867),
            .I(\b2v_inst6.countZ0Z_2 ));
    LocalMux I__7626 (
            .O(N__33864),
            .I(\b2v_inst6.countZ0Z_2 ));
    InMux I__7625 (
            .O(N__33859),
            .I(\b2v_inst6.un2_count_1_cry_1 ));
    InMux I__7624 (
            .O(N__33856),
            .I(\b2v_inst6.un2_count_1_cry_2 ));
    InMux I__7623 (
            .O(N__33853),
            .I(\b2v_inst6.un2_count_1_cry_3 ));
    InMux I__7622 (
            .O(N__33850),
            .I(\b2v_inst6.un2_count_1_cry_4 ));
    CascadeMux I__7621 (
            .O(N__33847),
            .I(\b2v_inst6.N_276_0_cascade_ ));
    InMux I__7620 (
            .O(N__33844),
            .I(N__33841));
    LocalMux I__7619 (
            .O(N__33841),
            .I(N__33838));
    Span4Mux_v I__7618 (
            .O(N__33838),
            .I(N__33835));
    Odrv4 I__7617 (
            .O(N__33835),
            .I(VR_READY_VCCINAUX_c));
    InMux I__7616 (
            .O(N__33832),
            .I(N__33829));
    LocalMux I__7615 (
            .O(N__33829),
            .I(N__33826));
    Odrv4 I__7614 (
            .O(N__33826),
            .I(VR_READY_VCCIN_c));
    CascadeMux I__7613 (
            .O(N__33823),
            .I(\b2v_inst6.N_192_cascade_ ));
    InMux I__7612 (
            .O(N__33820),
            .I(N__33814));
    InMux I__7611 (
            .O(N__33819),
            .I(N__33814));
    LocalMux I__7610 (
            .O(N__33814),
            .I(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ));
    CascadeMux I__7609 (
            .O(N__33811),
            .I(\b2v_inst6.curr_state_RNIUL1J2Z0Z_0_cascade_ ));
    InMux I__7608 (
            .O(N__33808),
            .I(N__33805));
    LocalMux I__7607 (
            .O(N__33805),
            .I(\b2v_inst6.N_276_0 ));
    CascadeMux I__7606 (
            .O(N__33802),
            .I(N__33798));
    IoInMux I__7605 (
            .O(N__33801),
            .I(N__33793));
    InMux I__7604 (
            .O(N__33798),
            .I(N__33785));
    InMux I__7603 (
            .O(N__33797),
            .I(N__33785));
    InMux I__7602 (
            .O(N__33796),
            .I(N__33785));
    LocalMux I__7601 (
            .O(N__33793),
            .I(N__33777));
    IoInMux I__7600 (
            .O(N__33792),
            .I(N__33774));
    LocalMux I__7599 (
            .O(N__33785),
            .I(N__33771));
    InMux I__7598 (
            .O(N__33784),
            .I(N__33768));
    InMux I__7597 (
            .O(N__33783),
            .I(N__33765));
    InMux I__7596 (
            .O(N__33782),
            .I(N__33762));
    InMux I__7595 (
            .O(N__33781),
            .I(N__33759));
    CascadeMux I__7594 (
            .O(N__33780),
            .I(N__33756));
    IoSpan4Mux I__7593 (
            .O(N__33777),
            .I(N__33749));
    LocalMux I__7592 (
            .O(N__33774),
            .I(N__33749));
    Span4Mux_v I__7591 (
            .O(N__33771),
            .I(N__33746));
    LocalMux I__7590 (
            .O(N__33768),
            .I(N__33743));
    LocalMux I__7589 (
            .O(N__33765),
            .I(N__33738));
    LocalMux I__7588 (
            .O(N__33762),
            .I(N__33738));
    LocalMux I__7587 (
            .O(N__33759),
            .I(N__33735));
    InMux I__7586 (
            .O(N__33756),
            .I(N__33730));
    InMux I__7585 (
            .O(N__33755),
            .I(N__33730));
    CascadeMux I__7584 (
            .O(N__33754),
            .I(N__33726));
    Span4Mux_s3_h I__7583 (
            .O(N__33749),
            .I(N__33720));
    Span4Mux_h I__7582 (
            .O(N__33746),
            .I(N__33720));
    Span4Mux_v I__7581 (
            .O(N__33743),
            .I(N__33715));
    Span4Mux_h I__7580 (
            .O(N__33738),
            .I(N__33715));
    Span4Mux_h I__7579 (
            .O(N__33735),
            .I(N__33710));
    LocalMux I__7578 (
            .O(N__33730),
            .I(N__33710));
    InMux I__7577 (
            .O(N__33729),
            .I(N__33705));
    InMux I__7576 (
            .O(N__33726),
            .I(N__33705));
    InMux I__7575 (
            .O(N__33725),
            .I(N__33702));
    Odrv4 I__7574 (
            .O(N__33720),
            .I(N_15_i_0_a4_1_N_3L3_1));
    Odrv4 I__7573 (
            .O(N__33715),
            .I(N_15_i_0_a4_1_N_3L3_1));
    Odrv4 I__7572 (
            .O(N__33710),
            .I(N_15_i_0_a4_1_N_3L3_1));
    LocalMux I__7571 (
            .O(N__33705),
            .I(N_15_i_0_a4_1_N_3L3_1));
    LocalMux I__7570 (
            .O(N__33702),
            .I(N_15_i_0_a4_1_N_3L3_1));
    CascadeMux I__7569 (
            .O(N__33691),
            .I(\b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ));
    InMux I__7568 (
            .O(N__33688),
            .I(N__33680));
    InMux I__7567 (
            .O(N__33687),
            .I(N__33675));
    InMux I__7566 (
            .O(N__33686),
            .I(N__33675));
    InMux I__7565 (
            .O(N__33685),
            .I(N__33668));
    InMux I__7564 (
            .O(N__33684),
            .I(N__33668));
    InMux I__7563 (
            .O(N__33683),
            .I(N__33668));
    LocalMux I__7562 (
            .O(N__33680),
            .I(N__33665));
    LocalMux I__7561 (
            .O(N__33675),
            .I(N__33662));
    LocalMux I__7560 (
            .O(N__33668),
            .I(N__33659));
    Span4Mux_s2_v I__7559 (
            .O(N__33665),
            .I(N__33656));
    Span4Mux_s2_v I__7558 (
            .O(N__33662),
            .I(N__33653));
    Span4Mux_s1_v I__7557 (
            .O(N__33659),
            .I(N__33650));
    Span4Mux_h I__7556 (
            .O(N__33656),
            .I(N__33647));
    Span4Mux_h I__7555 (
            .O(N__33653),
            .I(N__33644));
    Span4Mux_h I__7554 (
            .O(N__33650),
            .I(N__33641));
    Odrv4 I__7553 (
            .O(N__33647),
            .I(N_222));
    Odrv4 I__7552 (
            .O(N__33644),
            .I(N_222));
    Odrv4 I__7551 (
            .O(N__33641),
            .I(N_222));
    CascadeMux I__7550 (
            .O(N__33634),
            .I(N__33630));
    CascadeMux I__7549 (
            .O(N__33633),
            .I(N__33625));
    InMux I__7548 (
            .O(N__33630),
            .I(N__33622));
    InMux I__7547 (
            .O(N__33629),
            .I(N__33618));
    InMux I__7546 (
            .O(N__33628),
            .I(N__33614));
    InMux I__7545 (
            .O(N__33625),
            .I(N__33610));
    LocalMux I__7544 (
            .O(N__33622),
            .I(N__33607));
    InMux I__7543 (
            .O(N__33621),
            .I(N__33604));
    LocalMux I__7542 (
            .O(N__33618),
            .I(N__33601));
    CascadeMux I__7541 (
            .O(N__33617),
            .I(N__33598));
    LocalMux I__7540 (
            .O(N__33614),
            .I(N__33592));
    InMux I__7539 (
            .O(N__33613),
            .I(N__33589));
    LocalMux I__7538 (
            .O(N__33610),
            .I(N__33583));
    Span4Mux_h I__7537 (
            .O(N__33607),
            .I(N__33580));
    LocalMux I__7536 (
            .O(N__33604),
            .I(N__33577));
    Span4Mux_h I__7535 (
            .O(N__33601),
            .I(N__33574));
    InMux I__7534 (
            .O(N__33598),
            .I(N__33571));
    InMux I__7533 (
            .O(N__33597),
            .I(N__33566));
    InMux I__7532 (
            .O(N__33596),
            .I(N__33566));
    InMux I__7531 (
            .O(N__33595),
            .I(N__33563));
    Span12Mux_s6_h I__7530 (
            .O(N__33592),
            .I(N__33558));
    LocalMux I__7529 (
            .O(N__33589),
            .I(N__33558));
    InMux I__7528 (
            .O(N__33588),
            .I(N__33551));
    InMux I__7527 (
            .O(N__33587),
            .I(N__33551));
    InMux I__7526 (
            .O(N__33586),
            .I(N__33551));
    Span4Mux_h I__7525 (
            .O(N__33583),
            .I(N__33544));
    Span4Mux_h I__7524 (
            .O(N__33580),
            .I(N__33544));
    Span4Mux_h I__7523 (
            .O(N__33577),
            .I(N__33544));
    Odrv4 I__7522 (
            .O(N__33574),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__7521 (
            .O(N__33571),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__7520 (
            .O(N__33566),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__7519 (
            .O(N__33563),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv12 I__7518 (
            .O(N__33558),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    LocalMux I__7517 (
            .O(N__33551),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    Odrv4 I__7516 (
            .O(N__33544),
            .I(\b2v_inst11.dutycycleZ0Z_0 ));
    InMux I__7515 (
            .O(N__33529),
            .I(N__33526));
    LocalMux I__7514 (
            .O(N__33526),
            .I(N__33523));
    Odrv12 I__7513 (
            .O(N__33523),
            .I(\b2v_inst11.mult1_un159_sum_i ));
    CascadeMux I__7512 (
            .O(N__33520),
            .I(N__33517));
    InMux I__7511 (
            .O(N__33517),
            .I(N__33514));
    LocalMux I__7510 (
            .O(N__33514),
            .I(N__33511));
    Odrv4 I__7509 (
            .O(N__33511),
            .I(\b2v_inst11.mult1_un159_sum_cry_2_s ));
    InMux I__7508 (
            .O(N__33508),
            .I(N__33505));
    LocalMux I__7507 (
            .O(N__33505),
            .I(N__33502));
    Odrv12 I__7506 (
            .O(N__33502),
            .I(\b2v_inst11.mult1_un159_sum_cry_3_s ));
    CascadeMux I__7505 (
            .O(N__33499),
            .I(N__33496));
    InMux I__7504 (
            .O(N__33496),
            .I(N__33493));
    LocalMux I__7503 (
            .O(N__33493),
            .I(N__33490));
    Span4Mux_s1_h I__7502 (
            .O(N__33490),
            .I(N__33487));
    Odrv4 I__7501 (
            .O(N__33487),
            .I(\b2v_inst11.mult1_un54_sum_cry_3_s ));
    InMux I__7500 (
            .O(N__33484),
            .I(\b2v_inst11.mult1_un61_sum_cry_3 ));
    InMux I__7499 (
            .O(N__33481),
            .I(N__33478));
    LocalMux I__7498 (
            .O(N__33478),
            .I(N__33475));
    Odrv4 I__7497 (
            .O(N__33475),
            .I(\b2v_inst11.mult1_un54_sum_cry_4_s ));
    InMux I__7496 (
            .O(N__33472),
            .I(\b2v_inst11.mult1_un61_sum_cry_4 ));
    CascadeMux I__7495 (
            .O(N__33469),
            .I(N__33466));
    InMux I__7494 (
            .O(N__33466),
            .I(N__33463));
    LocalMux I__7493 (
            .O(N__33463),
            .I(N__33460));
    Odrv4 I__7492 (
            .O(N__33460),
            .I(\b2v_inst11.mult1_un54_sum_cry_5_s ));
    InMux I__7491 (
            .O(N__33457),
            .I(\b2v_inst11.mult1_un61_sum_cry_5 ));
    InMux I__7490 (
            .O(N__33454),
            .I(N__33451));
    LocalMux I__7489 (
            .O(N__33451),
            .I(N__33448));
    Odrv4 I__7488 (
            .O(N__33448),
            .I(\b2v_inst11.mult1_un54_sum_cry_6_s ));
    InMux I__7487 (
            .O(N__33445),
            .I(\b2v_inst11.mult1_un61_sum_cry_6 ));
    CascadeMux I__7486 (
            .O(N__33442),
            .I(N__33439));
    InMux I__7485 (
            .O(N__33439),
            .I(N__33436));
    LocalMux I__7484 (
            .O(N__33436),
            .I(N__33433));
    Odrv4 I__7483 (
            .O(N__33433),
            .I(\b2v_inst11.mult1_un61_sum_axb_8 ));
    InMux I__7482 (
            .O(N__33430),
            .I(\b2v_inst11.mult1_un61_sum_cry_7 ));
    CascadeMux I__7481 (
            .O(N__33427),
            .I(\b2v_inst11.mult1_un61_sum_s_8_cascade_ ));
    InMux I__7480 (
            .O(N__33424),
            .I(N__33421));
    LocalMux I__7479 (
            .O(N__33421),
            .I(N__33418));
    IoSpan4Mux I__7478 (
            .O(N__33418),
            .I(N__33415));
    Odrv4 I__7477 (
            .O(N__33415),
            .I(V33S_OK_c));
    InMux I__7476 (
            .O(N__33412),
            .I(N__33409));
    LocalMux I__7475 (
            .O(N__33409),
            .I(N__33406));
    Odrv4 I__7474 (
            .O(N__33406),
            .I(V5S_OK_c));
    IoInMux I__7473 (
            .O(N__33403),
            .I(N__33400));
    LocalMux I__7472 (
            .O(N__33400),
            .I(N__33396));
    IoInMux I__7471 (
            .O(N__33399),
            .I(N__33393));
    Span4Mux_s2_h I__7470 (
            .O(N__33396),
            .I(N__33390));
    LocalMux I__7469 (
            .O(N__33393),
            .I(N__33387));
    Span4Mux_v I__7468 (
            .O(N__33390),
            .I(N__33384));
    Span12Mux_s5_h I__7467 (
            .O(N__33387),
            .I(N__33381));
    Span4Mux_h I__7466 (
            .O(N__33384),
            .I(N__33378));
    Span12Mux_v I__7465 (
            .O(N__33381),
            .I(N__33375));
    Span4Mux_h I__7464 (
            .O(N__33378),
            .I(N__33372));
    Odrv12 I__7463 (
            .O(N__33375),
            .I(VCCIN_EN_c));
    Odrv4 I__7462 (
            .O(N__33372),
            .I(VCCIN_EN_c));
    InMux I__7461 (
            .O(N__33367),
            .I(\b2v_inst11.mult1_un89_sum_cry_7 ));
    InMux I__7460 (
            .O(N__33364),
            .I(N__33356));
    InMux I__7459 (
            .O(N__33363),
            .I(N__33349));
    InMux I__7458 (
            .O(N__33362),
            .I(N__33346));
    InMux I__7457 (
            .O(N__33361),
            .I(N__33343));
    InMux I__7456 (
            .O(N__33360),
            .I(N__33338));
    InMux I__7455 (
            .O(N__33359),
            .I(N__33338));
    LocalMux I__7454 (
            .O(N__33356),
            .I(N__33335));
    InMux I__7453 (
            .O(N__33355),
            .I(N__33332));
    CascadeMux I__7452 (
            .O(N__33354),
            .I(N__33329));
    CascadeMux I__7451 (
            .O(N__33353),
            .I(N__33326));
    InMux I__7450 (
            .O(N__33352),
            .I(N__33323));
    LocalMux I__7449 (
            .O(N__33349),
            .I(N__33317));
    LocalMux I__7448 (
            .O(N__33346),
            .I(N__33312));
    LocalMux I__7447 (
            .O(N__33343),
            .I(N__33312));
    LocalMux I__7446 (
            .O(N__33338),
            .I(N__33309));
    Span4Mux_s2_h I__7445 (
            .O(N__33335),
            .I(N__33304));
    LocalMux I__7444 (
            .O(N__33332),
            .I(N__33304));
    InMux I__7443 (
            .O(N__33329),
            .I(N__33301));
    InMux I__7442 (
            .O(N__33326),
            .I(N__33298));
    LocalMux I__7441 (
            .O(N__33323),
            .I(N__33295));
    InMux I__7440 (
            .O(N__33322),
            .I(N__33290));
    InMux I__7439 (
            .O(N__33321),
            .I(N__33290));
    InMux I__7438 (
            .O(N__33320),
            .I(N__33287));
    Span4Mux_h I__7437 (
            .O(N__33317),
            .I(N__33282));
    Span4Mux_h I__7436 (
            .O(N__33312),
            .I(N__33282));
    Span4Mux_v I__7435 (
            .O(N__33309),
            .I(N__33277));
    Span4Mux_h I__7434 (
            .O(N__33304),
            .I(N__33277));
    LocalMux I__7433 (
            .O(N__33301),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__7432 (
            .O(N__33298),
            .I(\b2v_inst11.dutycycle ));
    Odrv12 I__7431 (
            .O(N__33295),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__7430 (
            .O(N__33290),
            .I(\b2v_inst11.dutycycle ));
    LocalMux I__7429 (
            .O(N__33287),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__7428 (
            .O(N__33282),
            .I(\b2v_inst11.dutycycle ));
    Odrv4 I__7427 (
            .O(N__33277),
            .I(\b2v_inst11.dutycycle ));
    InMux I__7426 (
            .O(N__33262),
            .I(N__33258));
    CascadeMux I__7425 (
            .O(N__33261),
            .I(N__33255));
    LocalMux I__7424 (
            .O(N__33258),
            .I(N__33252));
    InMux I__7423 (
            .O(N__33255),
            .I(N__33249));
    Span4Mux_s2_h I__7422 (
            .O(N__33252),
            .I(N__33246));
    LocalMux I__7421 (
            .O(N__33249),
            .I(N__33243));
    Odrv4 I__7420 (
            .O(N__33246),
            .I(\b2v_inst11.mult1_un54_sum ));
    Odrv4 I__7419 (
            .O(N__33243),
            .I(\b2v_inst11.mult1_un54_sum ));
    InMux I__7418 (
            .O(N__33238),
            .I(N__33235));
    LocalMux I__7417 (
            .O(N__33235),
            .I(N__33232));
    Odrv12 I__7416 (
            .O(N__33232),
            .I(\b2v_inst11.mult1_un61_sum_i_8 ));
    InMux I__7415 (
            .O(N__33229),
            .I(N__33225));
    InMux I__7414 (
            .O(N__33228),
            .I(N__33222));
    LocalMux I__7413 (
            .O(N__33225),
            .I(N__33219));
    LocalMux I__7412 (
            .O(N__33222),
            .I(N__33216));
    Span4Mux_s2_h I__7411 (
            .O(N__33219),
            .I(N__33213));
    Span4Mux_s2_h I__7410 (
            .O(N__33216),
            .I(N__33210));
    Odrv4 I__7409 (
            .O(N__33213),
            .I(\b2v_inst11.mult1_un61_sum ));
    Odrv4 I__7408 (
            .O(N__33210),
            .I(\b2v_inst11.mult1_un61_sum ));
    InMux I__7407 (
            .O(N__33205),
            .I(N__33202));
    LocalMux I__7406 (
            .O(N__33202),
            .I(\b2v_inst11.mult1_un54_sum_i ));
    InMux I__7405 (
            .O(N__33199),
            .I(\b2v_inst11.mult1_un61_sum_cry_2 ));
    InMux I__7404 (
            .O(N__33196),
            .I(N__33193));
    LocalMux I__7403 (
            .O(N__33193),
            .I(\b2v_inst11.mult1_un89_sum_i_8 ));
    CascadeMux I__7402 (
            .O(N__33190),
            .I(N__33187));
    InMux I__7401 (
            .O(N__33187),
            .I(N__33184));
    LocalMux I__7400 (
            .O(N__33184),
            .I(N__33181));
    Span4Mux_v I__7399 (
            .O(N__33181),
            .I(N__33178));
    Odrv4 I__7398 (
            .O(N__33178),
            .I(\b2v_inst11.un85_clk_100khz_1 ));
    InMux I__7397 (
            .O(N__33175),
            .I(N__33172));
    LocalMux I__7396 (
            .O(N__33172),
            .I(\b2v_inst11.mult1_un82_sum_i_8 ));
    InMux I__7395 (
            .O(N__33169),
            .I(N__33165));
    InMux I__7394 (
            .O(N__33168),
            .I(N__33162));
    LocalMux I__7393 (
            .O(N__33165),
            .I(N__33159));
    LocalMux I__7392 (
            .O(N__33162),
            .I(N__33156));
    Span4Mux_s2_h I__7391 (
            .O(N__33159),
            .I(N__33153));
    Odrv4 I__7390 (
            .O(N__33156),
            .I(\b2v_inst11.mult1_un89_sum ));
    Odrv4 I__7389 (
            .O(N__33153),
            .I(\b2v_inst11.mult1_un89_sum ));
    InMux I__7388 (
            .O(N__33148),
            .I(N__33145));
    LocalMux I__7387 (
            .O(N__33145),
            .I(\b2v_inst11.mult1_un82_sum_i ));
    InMux I__7386 (
            .O(N__33142),
            .I(\b2v_inst11.mult1_un89_sum_cry_2 ));
    InMux I__7385 (
            .O(N__33139),
            .I(\b2v_inst11.mult1_un89_sum_cry_3 ));
    InMux I__7384 (
            .O(N__33136),
            .I(\b2v_inst11.mult1_un89_sum_cry_4 ));
    InMux I__7383 (
            .O(N__33133),
            .I(\b2v_inst11.mult1_un89_sum_cry_5 ));
    InMux I__7382 (
            .O(N__33130),
            .I(\b2v_inst11.mult1_un89_sum_cry_6 ));
    InMux I__7381 (
            .O(N__33127),
            .I(N__33124));
    LocalMux I__7380 (
            .O(N__33124),
            .I(N__33121));
    Span4Mux_h I__7379 (
            .O(N__33121),
            .I(N__33116));
    InMux I__7378 (
            .O(N__33120),
            .I(N__33113));
    InMux I__7377 (
            .O(N__33119),
            .I(N__33110));
    Odrv4 I__7376 (
            .O(N__33116),
            .I(\b2v_inst11.countZ0Z_12 ));
    LocalMux I__7375 (
            .O(N__33113),
            .I(\b2v_inst11.countZ0Z_12 ));
    LocalMux I__7374 (
            .O(N__33110),
            .I(\b2v_inst11.countZ0Z_12 ));
    CascadeMux I__7373 (
            .O(N__33103),
            .I(N__33100));
    InMux I__7372 (
            .O(N__33100),
            .I(N__33097));
    LocalMux I__7371 (
            .O(N__33097),
            .I(\b2v_inst11.N_5541_i ));
    InMux I__7370 (
            .O(N__33094),
            .I(N__33091));
    LocalMux I__7369 (
            .O(N__33091),
            .I(N__33088));
    Span4Mux_s3_h I__7368 (
            .O(N__33088),
            .I(N__33083));
    InMux I__7367 (
            .O(N__33087),
            .I(N__33080));
    InMux I__7366 (
            .O(N__33086),
            .I(N__33077));
    Odrv4 I__7365 (
            .O(N__33083),
            .I(\b2v_inst11.countZ0Z_13 ));
    LocalMux I__7364 (
            .O(N__33080),
            .I(\b2v_inst11.countZ0Z_13 ));
    LocalMux I__7363 (
            .O(N__33077),
            .I(\b2v_inst11.countZ0Z_13 ));
    CascadeMux I__7362 (
            .O(N__33070),
            .I(N__33067));
    InMux I__7361 (
            .O(N__33067),
            .I(N__33064));
    LocalMux I__7360 (
            .O(N__33064),
            .I(\b2v_inst11.N_5542_i ));
    InMux I__7359 (
            .O(N__33061),
            .I(N__33058));
    LocalMux I__7358 (
            .O(N__33058),
            .I(N__33055));
    Span4Mux_h I__7357 (
            .O(N__33055),
            .I(N__33052));
    Span4Mux_v I__7356 (
            .O(N__33052),
            .I(N__33047));
    InMux I__7355 (
            .O(N__33051),
            .I(N__33044));
    InMux I__7354 (
            .O(N__33050),
            .I(N__33041));
    Odrv4 I__7353 (
            .O(N__33047),
            .I(\b2v_inst11.countZ0Z_14 ));
    LocalMux I__7352 (
            .O(N__33044),
            .I(\b2v_inst11.countZ0Z_14 ));
    LocalMux I__7351 (
            .O(N__33041),
            .I(\b2v_inst11.countZ0Z_14 ));
    CascadeMux I__7350 (
            .O(N__33034),
            .I(N__33031));
    InMux I__7349 (
            .O(N__33031),
            .I(N__33028));
    LocalMux I__7348 (
            .O(N__33028),
            .I(\b2v_inst11.N_5543_i ));
    InMux I__7347 (
            .O(N__33025),
            .I(N__33022));
    LocalMux I__7346 (
            .O(N__33022),
            .I(N__33019));
    Span12Mux_s5_h I__7345 (
            .O(N__33019),
            .I(N__33014));
    InMux I__7344 (
            .O(N__33018),
            .I(N__33011));
    InMux I__7343 (
            .O(N__33017),
            .I(N__33008));
    Odrv12 I__7342 (
            .O(N__33014),
            .I(\b2v_inst11.countZ0Z_15 ));
    LocalMux I__7341 (
            .O(N__33011),
            .I(\b2v_inst11.countZ0Z_15 ));
    LocalMux I__7340 (
            .O(N__33008),
            .I(\b2v_inst11.countZ0Z_15 ));
    CascadeMux I__7339 (
            .O(N__33001),
            .I(N__32998));
    InMux I__7338 (
            .O(N__32998),
            .I(N__32995));
    LocalMux I__7337 (
            .O(N__32995),
            .I(\b2v_inst11.N_5544_i ));
    InMux I__7336 (
            .O(N__32992),
            .I(bfn_11_10_0_));
    CascadeMux I__7335 (
            .O(N__32989),
            .I(N__32984));
    InMux I__7334 (
            .O(N__32988),
            .I(N__32978));
    InMux I__7333 (
            .O(N__32987),
            .I(N__32978));
    InMux I__7332 (
            .O(N__32984),
            .I(N__32975));
    InMux I__7331 (
            .O(N__32983),
            .I(N__32972));
    LocalMux I__7330 (
            .O(N__32978),
            .I(N__32969));
    LocalMux I__7329 (
            .O(N__32975),
            .I(N__32966));
    LocalMux I__7328 (
            .O(N__32972),
            .I(N__32961));
    Span4Mux_s2_v I__7327 (
            .O(N__32969),
            .I(N__32961));
    Span12Mux_s6_v I__7326 (
            .O(N__32966),
            .I(N__32958));
    Span4Mux_v I__7325 (
            .O(N__32961),
            .I(N__32955));
    Odrv12 I__7324 (
            .O(N__32958),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__7323 (
            .O(N__32955),
            .I(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    InMux I__7322 (
            .O(N__32950),
            .I(N__32947));
    LocalMux I__7321 (
            .O(N__32947),
            .I(N__32944));
    Span4Mux_v I__7320 (
            .O(N__32944),
            .I(N__32941));
    Span4Mux_v I__7319 (
            .O(N__32941),
            .I(N__32936));
    InMux I__7318 (
            .O(N__32940),
            .I(N__32933));
    InMux I__7317 (
            .O(N__32939),
            .I(N__32930));
    Odrv4 I__7316 (
            .O(N__32936),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__7315 (
            .O(N__32933),
            .I(\b2v_inst11.countZ0Z_4 ));
    LocalMux I__7314 (
            .O(N__32930),
            .I(\b2v_inst11.countZ0Z_4 ));
    CascadeMux I__7313 (
            .O(N__32923),
            .I(N__32920));
    InMux I__7312 (
            .O(N__32920),
            .I(N__32917));
    LocalMux I__7311 (
            .O(N__32917),
            .I(\b2v_inst11.mult1_un138_sum_i_8 ));
    InMux I__7310 (
            .O(N__32914),
            .I(N__32911));
    LocalMux I__7309 (
            .O(N__32911),
            .I(\b2v_inst11.N_5533_i ));
    InMux I__7308 (
            .O(N__32908),
            .I(N__32905));
    LocalMux I__7307 (
            .O(N__32905),
            .I(N__32902));
    Span4Mux_v I__7306 (
            .O(N__32902),
            .I(N__32898));
    InMux I__7305 (
            .O(N__32901),
            .I(N__32895));
    Span4Mux_h I__7304 (
            .O(N__32898),
            .I(N__32889));
    LocalMux I__7303 (
            .O(N__32895),
            .I(N__32889));
    InMux I__7302 (
            .O(N__32894),
            .I(N__32886));
    Odrv4 I__7301 (
            .O(N__32889),
            .I(\b2v_inst11.countZ0Z_5 ));
    LocalMux I__7300 (
            .O(N__32886),
            .I(\b2v_inst11.countZ0Z_5 ));
    CascadeMux I__7299 (
            .O(N__32881),
            .I(N__32878));
    InMux I__7298 (
            .O(N__32878),
            .I(N__32875));
    LocalMux I__7297 (
            .O(N__32875),
            .I(N__32872));
    Span4Mux_v I__7296 (
            .O(N__32872),
            .I(N__32869));
    Odrv4 I__7295 (
            .O(N__32869),
            .I(\b2v_inst11.mult1_un131_sum_i_8 ));
    InMux I__7294 (
            .O(N__32866),
            .I(N__32863));
    LocalMux I__7293 (
            .O(N__32863),
            .I(\b2v_inst11.N_5534_i ));
    CascadeMux I__7292 (
            .O(N__32860),
            .I(N__32857));
    InMux I__7291 (
            .O(N__32857),
            .I(N__32854));
    LocalMux I__7290 (
            .O(N__32854),
            .I(\b2v_inst11.mult1_un124_sum_i_8 ));
    InMux I__7289 (
            .O(N__32851),
            .I(N__32848));
    LocalMux I__7288 (
            .O(N__32848),
            .I(N__32844));
    InMux I__7287 (
            .O(N__32847),
            .I(N__32841));
    Span12Mux_v I__7286 (
            .O(N__32844),
            .I(N__32837));
    LocalMux I__7285 (
            .O(N__32841),
            .I(N__32834));
    InMux I__7284 (
            .O(N__32840),
            .I(N__32831));
    Odrv12 I__7283 (
            .O(N__32837),
            .I(\b2v_inst11.countZ0Z_6 ));
    Odrv4 I__7282 (
            .O(N__32834),
            .I(\b2v_inst11.countZ0Z_6 ));
    LocalMux I__7281 (
            .O(N__32831),
            .I(\b2v_inst11.countZ0Z_6 ));
    InMux I__7280 (
            .O(N__32824),
            .I(N__32821));
    LocalMux I__7279 (
            .O(N__32821),
            .I(\b2v_inst11.N_5535_i ));
    InMux I__7278 (
            .O(N__32818),
            .I(N__32815));
    LocalMux I__7277 (
            .O(N__32815),
            .I(N__32812));
    Span4Mux_v I__7276 (
            .O(N__32812),
            .I(N__32808));
    InMux I__7275 (
            .O(N__32811),
            .I(N__32805));
    Span4Mux_v I__7274 (
            .O(N__32808),
            .I(N__32801));
    LocalMux I__7273 (
            .O(N__32805),
            .I(N__32798));
    InMux I__7272 (
            .O(N__32804),
            .I(N__32795));
    Span4Mux_h I__7271 (
            .O(N__32801),
            .I(N__32788));
    Span4Mux_s3_v I__7270 (
            .O(N__32798),
            .I(N__32788));
    LocalMux I__7269 (
            .O(N__32795),
            .I(N__32788));
    Odrv4 I__7268 (
            .O(N__32788),
            .I(\b2v_inst11.countZ0Z_7 ));
    CascadeMux I__7267 (
            .O(N__32785),
            .I(N__32782));
    InMux I__7266 (
            .O(N__32782),
            .I(N__32779));
    LocalMux I__7265 (
            .O(N__32779),
            .I(\b2v_inst11.mult1_un117_sum_i_8 ));
    InMux I__7264 (
            .O(N__32776),
            .I(N__32773));
    LocalMux I__7263 (
            .O(N__32773),
            .I(\b2v_inst11.N_5536_i ));
    InMux I__7262 (
            .O(N__32770),
            .I(N__32767));
    LocalMux I__7261 (
            .O(N__32767),
            .I(N__32763));
    InMux I__7260 (
            .O(N__32766),
            .I(N__32760));
    Span12Mux_s4_h I__7259 (
            .O(N__32763),
            .I(N__32756));
    LocalMux I__7258 (
            .O(N__32760),
            .I(N__32753));
    InMux I__7257 (
            .O(N__32759),
            .I(N__32750));
    Odrv12 I__7256 (
            .O(N__32756),
            .I(\b2v_inst11.countZ0Z_8 ));
    Odrv4 I__7255 (
            .O(N__32753),
            .I(\b2v_inst11.countZ0Z_8 ));
    LocalMux I__7254 (
            .O(N__32750),
            .I(\b2v_inst11.countZ0Z_8 ));
    InMux I__7253 (
            .O(N__32743),
            .I(N__32740));
    LocalMux I__7252 (
            .O(N__32740),
            .I(N__32737));
    Odrv4 I__7251 (
            .O(N__32737),
            .I(\b2v_inst11.mult1_un110_sum_i_8 ));
    CascadeMux I__7250 (
            .O(N__32734),
            .I(N__32731));
    InMux I__7249 (
            .O(N__32731),
            .I(N__32728));
    LocalMux I__7248 (
            .O(N__32728),
            .I(\b2v_inst11.N_5537_i ));
    InMux I__7247 (
            .O(N__32725),
            .I(N__32722));
    LocalMux I__7246 (
            .O(N__32722),
            .I(N__32719));
    Span4Mux_v I__7245 (
            .O(N__32719),
            .I(N__32715));
    InMux I__7244 (
            .O(N__32718),
            .I(N__32712));
    Span4Mux_h I__7243 (
            .O(N__32715),
            .I(N__32706));
    LocalMux I__7242 (
            .O(N__32712),
            .I(N__32706));
    InMux I__7241 (
            .O(N__32711),
            .I(N__32703));
    Span4Mux_v I__7240 (
            .O(N__32706),
            .I(N__32700));
    LocalMux I__7239 (
            .O(N__32703),
            .I(\b2v_inst11.countZ0Z_9 ));
    Odrv4 I__7238 (
            .O(N__32700),
            .I(\b2v_inst11.countZ0Z_9 ));
    CascadeMux I__7237 (
            .O(N__32695),
            .I(N__32692));
    InMux I__7236 (
            .O(N__32692),
            .I(N__32689));
    LocalMux I__7235 (
            .O(N__32689),
            .I(N__32686));
    Span4Mux_s3_h I__7234 (
            .O(N__32686),
            .I(N__32683));
    Odrv4 I__7233 (
            .O(N__32683),
            .I(\b2v_inst11.mult1_un103_sum_i_8 ));
    InMux I__7232 (
            .O(N__32680),
            .I(N__32677));
    LocalMux I__7231 (
            .O(N__32677),
            .I(\b2v_inst11.N_5538_i ));
    InMux I__7230 (
            .O(N__32674),
            .I(N__32670));
    CascadeMux I__7229 (
            .O(N__32673),
            .I(N__32667));
    LocalMux I__7228 (
            .O(N__32670),
            .I(N__32664));
    InMux I__7227 (
            .O(N__32667),
            .I(N__32661));
    Span4Mux_v I__7226 (
            .O(N__32664),
            .I(N__32658));
    LocalMux I__7225 (
            .O(N__32661),
            .I(N__32654));
    Span4Mux_h I__7224 (
            .O(N__32658),
            .I(N__32651));
    InMux I__7223 (
            .O(N__32657),
            .I(N__32648));
    Span4Mux_h I__7222 (
            .O(N__32654),
            .I(N__32645));
    Odrv4 I__7221 (
            .O(N__32651),
            .I(\b2v_inst11.countZ0Z_10 ));
    LocalMux I__7220 (
            .O(N__32648),
            .I(\b2v_inst11.countZ0Z_10 ));
    Odrv4 I__7219 (
            .O(N__32645),
            .I(\b2v_inst11.countZ0Z_10 ));
    CascadeMux I__7218 (
            .O(N__32638),
            .I(N__32635));
    InMux I__7217 (
            .O(N__32635),
            .I(N__32632));
    LocalMux I__7216 (
            .O(N__32632),
            .I(\b2v_inst11.N_5539_i ));
    InMux I__7215 (
            .O(N__32629),
            .I(N__32626));
    LocalMux I__7214 (
            .O(N__32626),
            .I(N__32622));
    InMux I__7213 (
            .O(N__32625),
            .I(N__32619));
    Span4Mux_v I__7212 (
            .O(N__32622),
            .I(N__32616));
    LocalMux I__7211 (
            .O(N__32619),
            .I(N__32612));
    Span4Mux_h I__7210 (
            .O(N__32616),
            .I(N__32609));
    InMux I__7209 (
            .O(N__32615),
            .I(N__32606));
    Span4Mux_h I__7208 (
            .O(N__32612),
            .I(N__32603));
    Odrv4 I__7207 (
            .O(N__32609),
            .I(\b2v_inst11.countZ0Z_11 ));
    LocalMux I__7206 (
            .O(N__32606),
            .I(\b2v_inst11.countZ0Z_11 ));
    Odrv4 I__7205 (
            .O(N__32603),
            .I(\b2v_inst11.countZ0Z_11 ));
    CascadeMux I__7204 (
            .O(N__32596),
            .I(N__32593));
    InMux I__7203 (
            .O(N__32593),
            .I(N__32590));
    LocalMux I__7202 (
            .O(N__32590),
            .I(\b2v_inst11.N_5540_i ));
    InMux I__7201 (
            .O(N__32587),
            .I(N__32583));
    CascadeMux I__7200 (
            .O(N__32586),
            .I(N__32579));
    LocalMux I__7199 (
            .O(N__32583),
            .I(N__32575));
    InMux I__7198 (
            .O(N__32582),
            .I(N__32570));
    InMux I__7197 (
            .O(N__32579),
            .I(N__32570));
    InMux I__7196 (
            .O(N__32578),
            .I(N__32567));
    Odrv12 I__7195 (
            .O(N__32575),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__7194 (
            .O(N__32570),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    LocalMux I__7193 (
            .O(N__32567),
            .I(\b2v_inst11.mult1_un117_sum_s_8 ));
    InMux I__7192 (
            .O(N__32560),
            .I(N__32557));
    LocalMux I__7191 (
            .O(N__32557),
            .I(N__32553));
    CascadeMux I__7190 (
            .O(N__32556),
            .I(N__32549));
    Span4Mux_h I__7189 (
            .O(N__32553),
            .I(N__32543));
    InMux I__7188 (
            .O(N__32552),
            .I(N__32540));
    InMux I__7187 (
            .O(N__32549),
            .I(N__32533));
    InMux I__7186 (
            .O(N__32548),
            .I(N__32533));
    InMux I__7185 (
            .O(N__32547),
            .I(N__32533));
    InMux I__7184 (
            .O(N__32546),
            .I(N__32530));
    Odrv4 I__7183 (
            .O(N__32543),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__7182 (
            .O(N__32540),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__7181 (
            .O(N__32533),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    LocalMux I__7180 (
            .O(N__32530),
            .I(\b2v_inst11.mult1_un124_sum_s_8 ));
    InMux I__7179 (
            .O(N__32521),
            .I(N__32516));
    CascadeMux I__7178 (
            .O(N__32520),
            .I(N__32513));
    CascadeMux I__7177 (
            .O(N__32519),
            .I(N__32510));
    LocalMux I__7176 (
            .O(N__32516),
            .I(N__32506));
    InMux I__7175 (
            .O(N__32513),
            .I(N__32503));
    InMux I__7174 (
            .O(N__32510),
            .I(N__32498));
    InMux I__7173 (
            .O(N__32509),
            .I(N__32498));
    Span4Mux_v I__7172 (
            .O(N__32506),
            .I(N__32494));
    LocalMux I__7171 (
            .O(N__32503),
            .I(N__32489));
    LocalMux I__7170 (
            .O(N__32498),
            .I(N__32489));
    InMux I__7169 (
            .O(N__32497),
            .I(N__32486));
    Odrv4 I__7168 (
            .O(N__32494),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    Odrv4 I__7167 (
            .O(N__32489),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    LocalMux I__7166 (
            .O(N__32486),
            .I(\b2v_inst11.mult1_un145_sum_s_8 ));
    InMux I__7165 (
            .O(N__32479),
            .I(N__32476));
    LocalMux I__7164 (
            .O(N__32476),
            .I(N__32472));
    CascadeMux I__7163 (
            .O(N__32475),
            .I(N__32469));
    Span4Mux_v I__7162 (
            .O(N__32472),
            .I(N__32463));
    InMux I__7161 (
            .O(N__32469),
            .I(N__32456));
    InMux I__7160 (
            .O(N__32468),
            .I(N__32456));
    InMux I__7159 (
            .O(N__32467),
            .I(N__32456));
    InMux I__7158 (
            .O(N__32466),
            .I(N__32453));
    Odrv4 I__7157 (
            .O(N__32463),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__7156 (
            .O(N__32456),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    LocalMux I__7155 (
            .O(N__32453),
            .I(\b2v_inst11.mult1_un138_sum_s_8 ));
    InMux I__7154 (
            .O(N__32446),
            .I(N__32443));
    LocalMux I__7153 (
            .O(N__32443),
            .I(N__32440));
    Span4Mux_v I__7152 (
            .O(N__32440),
            .I(N__32433));
    InMux I__7151 (
            .O(N__32439),
            .I(N__32430));
    InMux I__7150 (
            .O(N__32438),
            .I(N__32427));
    InMux I__7149 (
            .O(N__32437),
            .I(N__32422));
    InMux I__7148 (
            .O(N__32436),
            .I(N__32422));
    Span4Mux_h I__7147 (
            .O(N__32433),
            .I(N__32417));
    LocalMux I__7146 (
            .O(N__32430),
            .I(N__32417));
    LocalMux I__7145 (
            .O(N__32427),
            .I(\b2v_inst11.countZ0Z_0 ));
    LocalMux I__7144 (
            .O(N__32422),
            .I(\b2v_inst11.countZ0Z_0 ));
    Odrv4 I__7143 (
            .O(N__32417),
            .I(\b2v_inst11.countZ0Z_0 ));
    InMux I__7142 (
            .O(N__32410),
            .I(N__32407));
    LocalMux I__7141 (
            .O(N__32407),
            .I(\b2v_inst11.un1_count_cry_0_i ));
    InMux I__7140 (
            .O(N__32404),
            .I(N__32401));
    LocalMux I__7139 (
            .O(N__32401),
            .I(N__32397));
    CascadeMux I__7138 (
            .O(N__32400),
            .I(N__32394));
    Span4Mux_v I__7137 (
            .O(N__32397),
            .I(N__32390));
    InMux I__7136 (
            .O(N__32394),
            .I(N__32387));
    InMux I__7135 (
            .O(N__32393),
            .I(N__32384));
    Span4Mux_h I__7134 (
            .O(N__32390),
            .I(N__32379));
    LocalMux I__7133 (
            .O(N__32387),
            .I(N__32379));
    LocalMux I__7132 (
            .O(N__32384),
            .I(\b2v_inst11.countZ0Z_1 ));
    Odrv4 I__7131 (
            .O(N__32379),
            .I(\b2v_inst11.countZ0Z_1 ));
    InMux I__7130 (
            .O(N__32374),
            .I(N__32371));
    LocalMux I__7129 (
            .O(N__32371),
            .I(\b2v_inst11.N_5530_i ));
    InMux I__7128 (
            .O(N__32368),
            .I(N__32365));
    LocalMux I__7127 (
            .O(N__32365),
            .I(N__32362));
    Span4Mux_s1_h I__7126 (
            .O(N__32362),
            .I(N__32358));
    InMux I__7125 (
            .O(N__32361),
            .I(N__32354));
    Span4Mux_v I__7124 (
            .O(N__32358),
            .I(N__32351));
    InMux I__7123 (
            .O(N__32357),
            .I(N__32348));
    LocalMux I__7122 (
            .O(N__32354),
            .I(N__32345));
    Span4Mux_h I__7121 (
            .O(N__32351),
            .I(N__32340));
    LocalMux I__7120 (
            .O(N__32348),
            .I(N__32340));
    Span4Mux_h I__7119 (
            .O(N__32345),
            .I(N__32337));
    Odrv4 I__7118 (
            .O(N__32340),
            .I(\b2v_inst11.countZ0Z_2 ));
    Odrv4 I__7117 (
            .O(N__32337),
            .I(\b2v_inst11.countZ0Z_2 ));
    CascadeMux I__7116 (
            .O(N__32332),
            .I(N__32329));
    InMux I__7115 (
            .O(N__32329),
            .I(N__32326));
    LocalMux I__7114 (
            .O(N__32326),
            .I(\b2v_inst11.un85_clk_100khz_2 ));
    InMux I__7113 (
            .O(N__32323),
            .I(N__32320));
    LocalMux I__7112 (
            .O(N__32320),
            .I(\b2v_inst11.N_5531_i ));
    InMux I__7111 (
            .O(N__32317),
            .I(N__32314));
    LocalMux I__7110 (
            .O(N__32314),
            .I(N__32311));
    Span4Mux_v I__7109 (
            .O(N__32311),
            .I(N__32307));
    CascadeMux I__7108 (
            .O(N__32310),
            .I(N__32303));
    Span4Mux_v I__7107 (
            .O(N__32307),
            .I(N__32300));
    InMux I__7106 (
            .O(N__32306),
            .I(N__32297));
    InMux I__7105 (
            .O(N__32303),
            .I(N__32294));
    Odrv4 I__7104 (
            .O(N__32300),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__7103 (
            .O(N__32297),
            .I(\b2v_inst11.countZ0Z_3 ));
    LocalMux I__7102 (
            .O(N__32294),
            .I(\b2v_inst11.countZ0Z_3 ));
    CascadeMux I__7101 (
            .O(N__32287),
            .I(N__32284));
    InMux I__7100 (
            .O(N__32284),
            .I(N__32281));
    LocalMux I__7099 (
            .O(N__32281),
            .I(N__32278));
    Odrv4 I__7098 (
            .O(N__32278),
            .I(\b2v_inst11.mult1_un145_sum_i_8 ));
    InMux I__7097 (
            .O(N__32275),
            .I(N__32272));
    LocalMux I__7096 (
            .O(N__32272),
            .I(\b2v_inst11.N_5532_i ));
    InMux I__7095 (
            .O(N__32269),
            .I(N__32266));
    LocalMux I__7094 (
            .O(N__32266),
            .I(N__32263));
    Odrv12 I__7093 (
            .O(N__32263),
            .I(\b2v_inst5.un2_count_1_axb_5 ));
    InMux I__7092 (
            .O(N__32260),
            .I(N__32257));
    LocalMux I__7091 (
            .O(N__32257),
            .I(\b2v_inst5.count_1_6 ));
    InMux I__7090 (
            .O(N__32254),
            .I(N__32248));
    InMux I__7089 (
            .O(N__32253),
            .I(N__32248));
    LocalMux I__7088 (
            .O(N__32248),
            .I(N__32245));
    Odrv4 I__7087 (
            .O(N__32245),
            .I(\b2v_inst5.count_rst_8 ));
    InMux I__7086 (
            .O(N__32242),
            .I(N__32239));
    LocalMux I__7085 (
            .O(N__32239),
            .I(N__32236));
    Odrv12 I__7084 (
            .O(N__32236),
            .I(\b2v_inst5.countZ0Z_6 ));
    InMux I__7083 (
            .O(N__32233),
            .I(N__32228));
    InMux I__7082 (
            .O(N__32232),
            .I(N__32223));
    InMux I__7081 (
            .O(N__32231),
            .I(N__32223));
    LocalMux I__7080 (
            .O(N__32228),
            .I(N__32218));
    LocalMux I__7079 (
            .O(N__32223),
            .I(N__32218));
    Odrv4 I__7078 (
            .O(N__32218),
            .I(\b2v_inst5.count_rst_9 ));
    CascadeMux I__7077 (
            .O(N__32215),
            .I(\b2v_inst5.countZ0Z_6_cascade_ ));
    InMux I__7076 (
            .O(N__32212),
            .I(N__32206));
    InMux I__7075 (
            .O(N__32211),
            .I(N__32206));
    LocalMux I__7074 (
            .O(N__32206),
            .I(\b2v_inst5.count_1_5 ));
    InMux I__7073 (
            .O(N__32203),
            .I(N__32200));
    LocalMux I__7072 (
            .O(N__32200),
            .I(N__32197));
    Span4Mux_v I__7071 (
            .O(N__32197),
            .I(N__32194));
    Odrv4 I__7070 (
            .O(N__32194),
            .I(\b2v_inst5.un12_clk_100khz_3 ));
    InMux I__7069 (
            .O(N__32191),
            .I(N__32188));
    LocalMux I__7068 (
            .O(N__32188),
            .I(N__32185));
    Odrv4 I__7067 (
            .O(N__32185),
            .I(\b2v_inst5.un2_count_1_axb_7 ));
    InMux I__7066 (
            .O(N__32182),
            .I(N__32163));
    InMux I__7065 (
            .O(N__32181),
            .I(N__32163));
    InMux I__7064 (
            .O(N__32180),
            .I(N__32163));
    InMux I__7063 (
            .O(N__32179),
            .I(N__32160));
    InMux I__7062 (
            .O(N__32178),
            .I(N__32155));
    InMux I__7061 (
            .O(N__32177),
            .I(N__32155));
    InMux I__7060 (
            .O(N__32176),
            .I(N__32150));
    InMux I__7059 (
            .O(N__32175),
            .I(N__32150));
    SRMux I__7058 (
            .O(N__32174),
            .I(N__32147));
    SRMux I__7057 (
            .O(N__32173),
            .I(N__32144));
    SRMux I__7056 (
            .O(N__32172),
            .I(N__32136));
    SRMux I__7055 (
            .O(N__32171),
            .I(N__32132));
    SRMux I__7054 (
            .O(N__32170),
            .I(N__32129));
    LocalMux I__7053 (
            .O(N__32163),
            .I(N__32120));
    LocalMux I__7052 (
            .O(N__32160),
            .I(N__32120));
    LocalMux I__7051 (
            .O(N__32155),
            .I(N__32120));
    LocalMux I__7050 (
            .O(N__32150),
            .I(N__32120));
    LocalMux I__7049 (
            .O(N__32147),
            .I(N__32117));
    LocalMux I__7048 (
            .O(N__32144),
            .I(N__32114));
    InMux I__7047 (
            .O(N__32143),
            .I(N__32103));
    InMux I__7046 (
            .O(N__32142),
            .I(N__32103));
    InMux I__7045 (
            .O(N__32141),
            .I(N__32103));
    InMux I__7044 (
            .O(N__32140),
            .I(N__32103));
    InMux I__7043 (
            .O(N__32139),
            .I(N__32103));
    LocalMux I__7042 (
            .O(N__32136),
            .I(N__32100));
    SRMux I__7041 (
            .O(N__32135),
            .I(N__32097));
    LocalMux I__7040 (
            .O(N__32132),
            .I(N__32082));
    LocalMux I__7039 (
            .O(N__32129),
            .I(N__32077));
    Span4Mux_s3_v I__7038 (
            .O(N__32120),
            .I(N__32077));
    Span4Mux_s1_h I__7037 (
            .O(N__32117),
            .I(N__32070));
    Span4Mux_h I__7036 (
            .O(N__32114),
            .I(N__32070));
    LocalMux I__7035 (
            .O(N__32103),
            .I(N__32070));
    Span4Mux_v I__7034 (
            .O(N__32100),
            .I(N__32067));
    LocalMux I__7033 (
            .O(N__32097),
            .I(N__32064));
    InMux I__7032 (
            .O(N__32096),
            .I(N__32057));
    InMux I__7031 (
            .O(N__32095),
            .I(N__32057));
    InMux I__7030 (
            .O(N__32094),
            .I(N__32057));
    InMux I__7029 (
            .O(N__32093),
            .I(N__32046));
    SRMux I__7028 (
            .O(N__32092),
            .I(N__32046));
    InMux I__7027 (
            .O(N__32091),
            .I(N__32046));
    InMux I__7026 (
            .O(N__32090),
            .I(N__32046));
    InMux I__7025 (
            .O(N__32089),
            .I(N__32046));
    InMux I__7024 (
            .O(N__32088),
            .I(N__32037));
    InMux I__7023 (
            .O(N__32087),
            .I(N__32037));
    InMux I__7022 (
            .O(N__32086),
            .I(N__32037));
    InMux I__7021 (
            .O(N__32085),
            .I(N__32037));
    Span4Mux_v I__7020 (
            .O(N__32082),
            .I(N__32032));
    Span4Mux_v I__7019 (
            .O(N__32077),
            .I(N__32032));
    Span4Mux_v I__7018 (
            .O(N__32070),
            .I(N__32029));
    Span4Mux_v I__7017 (
            .O(N__32067),
            .I(N__32026));
    Span4Mux_v I__7016 (
            .O(N__32064),
            .I(N__32023));
    LocalMux I__7015 (
            .O(N__32057),
            .I(N__32020));
    LocalMux I__7014 (
            .O(N__32046),
            .I(N__32015));
    LocalMux I__7013 (
            .O(N__32037),
            .I(N__32015));
    Span4Mux_v I__7012 (
            .O(N__32032),
            .I(N__32010));
    Span4Mux_v I__7011 (
            .O(N__32029),
            .I(N__32010));
    Span4Mux_h I__7010 (
            .O(N__32026),
            .I(N__32007));
    Span4Mux_h I__7009 (
            .O(N__32023),
            .I(N__32002));
    Span4Mux_v I__7008 (
            .O(N__32020),
            .I(N__32002));
    Span12Mux_v I__7007 (
            .O(N__32015),
            .I(N__31999));
    Span4Mux_h I__7006 (
            .O(N__32010),
            .I(N__31996));
    Odrv4 I__7005 (
            .O(N__32007),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__7004 (
            .O(N__32002),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv12 I__7003 (
            .O(N__31999),
            .I(\b2v_inst5.count_0_sqmuxa ));
    Odrv4 I__7002 (
            .O(N__31996),
            .I(\b2v_inst5.count_0_sqmuxa ));
    InMux I__7001 (
            .O(N__31987),
            .I(N__31981));
    InMux I__7000 (
            .O(N__31986),
            .I(N__31981));
    LocalMux I__6999 (
            .O(N__31981),
            .I(\b2v_inst5.count_1_7 ));
    InMux I__6998 (
            .O(N__31978),
            .I(N__31969));
    InMux I__6997 (
            .O(N__31977),
            .I(N__31969));
    InMux I__6996 (
            .O(N__31976),
            .I(N__31969));
    LocalMux I__6995 (
            .O(N__31969),
            .I(N__31966));
    Odrv4 I__6994 (
            .O(N__31966),
            .I(\b2v_inst5.count_rst_7 ));
    CascadeMux I__6993 (
            .O(N__31963),
            .I(N__31960));
    InMux I__6992 (
            .O(N__31960),
            .I(N__31957));
    LocalMux I__6991 (
            .O(N__31957),
            .I(N__31953));
    InMux I__6990 (
            .O(N__31956),
            .I(N__31950));
    Span4Mux_v I__6989 (
            .O(N__31953),
            .I(N__31945));
    LocalMux I__6988 (
            .O(N__31950),
            .I(N__31945));
    Odrv4 I__6987 (
            .O(N__31945),
            .I(\b2v_inst5.countZ0Z_11 ));
    InMux I__6986 (
            .O(N__31942),
            .I(N__31934));
    CEMux I__6985 (
            .O(N__31941),
            .I(N__31934));
    InMux I__6984 (
            .O(N__31940),
            .I(N__31929));
    CEMux I__6983 (
            .O(N__31939),
            .I(N__31929));
    LocalMux I__6982 (
            .O(N__31934),
            .I(N__31924));
    LocalMux I__6981 (
            .O(N__31929),
            .I(N__31921));
    CEMux I__6980 (
            .O(N__31928),
            .I(N__31918));
    CEMux I__6979 (
            .O(N__31927),
            .I(N__31915));
    Span4Mux_v I__6978 (
            .O(N__31924),
            .I(N__31900));
    Span4Mux_h I__6977 (
            .O(N__31921),
            .I(N__31900));
    LocalMux I__6976 (
            .O(N__31918),
            .I(N__31900));
    LocalMux I__6975 (
            .O(N__31915),
            .I(N__31897));
    InMux I__6974 (
            .O(N__31914),
            .I(N__31888));
    InMux I__6973 (
            .O(N__31913),
            .I(N__31888));
    InMux I__6972 (
            .O(N__31912),
            .I(N__31888));
    InMux I__6971 (
            .O(N__31911),
            .I(N__31888));
    InMux I__6970 (
            .O(N__31910),
            .I(N__31875));
    CEMux I__6969 (
            .O(N__31909),
            .I(N__31875));
    InMux I__6968 (
            .O(N__31908),
            .I(N__31865));
    CEMux I__6967 (
            .O(N__31907),
            .I(N__31865));
    Span4Mux_s3_v I__6966 (
            .O(N__31900),
            .I(N__31858));
    Span4Mux_s1_h I__6965 (
            .O(N__31897),
            .I(N__31858));
    LocalMux I__6964 (
            .O(N__31888),
            .I(N__31858));
    InMux I__6963 (
            .O(N__31887),
            .I(N__31849));
    InMux I__6962 (
            .O(N__31886),
            .I(N__31849));
    InMux I__6961 (
            .O(N__31885),
            .I(N__31849));
    InMux I__6960 (
            .O(N__31884),
            .I(N__31849));
    CEMux I__6959 (
            .O(N__31883),
            .I(N__31840));
    InMux I__6958 (
            .O(N__31882),
            .I(N__31840));
    InMux I__6957 (
            .O(N__31881),
            .I(N__31840));
    InMux I__6956 (
            .O(N__31880),
            .I(N__31840));
    LocalMux I__6955 (
            .O(N__31875),
            .I(N__31837));
    InMux I__6954 (
            .O(N__31874),
            .I(N__31828));
    InMux I__6953 (
            .O(N__31873),
            .I(N__31828));
    InMux I__6952 (
            .O(N__31872),
            .I(N__31828));
    InMux I__6951 (
            .O(N__31871),
            .I(N__31823));
    InMux I__6950 (
            .O(N__31870),
            .I(N__31823));
    LocalMux I__6949 (
            .O(N__31865),
            .I(N__31820));
    Span4Mux_h I__6948 (
            .O(N__31858),
            .I(N__31813));
    LocalMux I__6947 (
            .O(N__31849),
            .I(N__31813));
    LocalMux I__6946 (
            .O(N__31840),
            .I(N__31813));
    Span4Mux_h I__6945 (
            .O(N__31837),
            .I(N__31810));
    InMux I__6944 (
            .O(N__31836),
            .I(N__31805));
    InMux I__6943 (
            .O(N__31835),
            .I(N__31805));
    LocalMux I__6942 (
            .O(N__31828),
            .I(N__31800));
    LocalMux I__6941 (
            .O(N__31823),
            .I(N__31800));
    Span4Mux_v I__6940 (
            .O(N__31820),
            .I(N__31795));
    Span4Mux_v I__6939 (
            .O(N__31813),
            .I(N__31795));
    Span4Mux_v I__6938 (
            .O(N__31810),
            .I(N__31792));
    LocalMux I__6937 (
            .O(N__31805),
            .I(N__31789));
    Sp12to4 I__6936 (
            .O(N__31800),
            .I(N__31786));
    Span4Mux_v I__6935 (
            .O(N__31795),
            .I(N__31783));
    Span4Mux_v I__6934 (
            .O(N__31792),
            .I(N__31780));
    Span4Mux_v I__6933 (
            .O(N__31789),
            .I(N__31777));
    Span12Mux_v I__6932 (
            .O(N__31786),
            .I(N__31774));
    Span4Mux_h I__6931 (
            .O(N__31783),
            .I(N__31771));
    Odrv4 I__6930 (
            .O(N__31780),
            .I(\b2v_inst5.curr_state_RNIFLPH1Z0Z_1 ));
    Odrv4 I__6929 (
            .O(N__31777),
            .I(\b2v_inst5.curr_state_RNIFLPH1Z0Z_1 ));
    Odrv12 I__6928 (
            .O(N__31774),
            .I(\b2v_inst5.curr_state_RNIFLPH1Z0Z_1 ));
    Odrv4 I__6927 (
            .O(N__31771),
            .I(\b2v_inst5.curr_state_RNIFLPH1Z0Z_1 ));
    CascadeMux I__6926 (
            .O(N__31762),
            .I(N__31759));
    InMux I__6925 (
            .O(N__31759),
            .I(N__31756));
    LocalMux I__6924 (
            .O(N__31756),
            .I(N__31753));
    Span4Mux_v I__6923 (
            .O(N__31753),
            .I(N__31750));
    Odrv4 I__6922 (
            .O(N__31750),
            .I(\b2v_inst5.un12_clk_100khz_2 ));
    CascadeMux I__6921 (
            .O(N__31747),
            .I(N__31743));
    CascadeMux I__6920 (
            .O(N__31746),
            .I(N__31740));
    InMux I__6919 (
            .O(N__31743),
            .I(N__31736));
    InMux I__6918 (
            .O(N__31740),
            .I(N__31731));
    InMux I__6917 (
            .O(N__31739),
            .I(N__31731));
    LocalMux I__6916 (
            .O(N__31736),
            .I(N__31727));
    LocalMux I__6915 (
            .O(N__31731),
            .I(N__31724));
    InMux I__6914 (
            .O(N__31730),
            .I(N__31721));
    Span4Mux_s2_v I__6913 (
            .O(N__31727),
            .I(N__31716));
    Span4Mux_s2_v I__6912 (
            .O(N__31724),
            .I(N__31716));
    LocalMux I__6911 (
            .O(N__31721),
            .I(N__31713));
    Span4Mux_v I__6910 (
            .O(N__31716),
            .I(N__31710));
    Span4Mux_v I__6909 (
            .O(N__31713),
            .I(N__31707));
    Span4Mux_v I__6908 (
            .O(N__31710),
            .I(N__31703));
    Sp12to4 I__6907 (
            .O(N__31707),
            .I(N__31700));
    InMux I__6906 (
            .O(N__31706),
            .I(N__31697));
    Odrv4 I__6905 (
            .O(N__31703),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    Odrv12 I__6904 (
            .O(N__31700),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    LocalMux I__6903 (
            .O(N__31697),
            .I(\b2v_inst11.mult1_un152_sum_s_8 ));
    InMux I__6902 (
            .O(N__31690),
            .I(N__31686));
    CascadeMux I__6901 (
            .O(N__31689),
            .I(N__31682));
    LocalMux I__6900 (
            .O(N__31686),
            .I(N__31678));
    InMux I__6899 (
            .O(N__31685),
            .I(N__31673));
    InMux I__6898 (
            .O(N__31682),
            .I(N__31673));
    InMux I__6897 (
            .O(N__31681),
            .I(N__31670));
    Odrv4 I__6896 (
            .O(N__31678),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__6895 (
            .O(N__31673),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    LocalMux I__6894 (
            .O(N__31670),
            .I(\b2v_inst11.mult1_un110_sum_s_8 ));
    CascadeMux I__6893 (
            .O(N__31663),
            .I(\b2v_inst5.count_rst_5_cascade_ ));
    InMux I__6892 (
            .O(N__31660),
            .I(N__31656));
    InMux I__6891 (
            .O(N__31659),
            .I(N__31653));
    LocalMux I__6890 (
            .O(N__31656),
            .I(\b2v_inst5.un2_count_1_axb_9 ));
    LocalMux I__6889 (
            .O(N__31653),
            .I(\b2v_inst5.un2_count_1_axb_9 ));
    CascadeMux I__6888 (
            .O(N__31648),
            .I(N__31644));
    InMux I__6887 (
            .O(N__31647),
            .I(N__31639));
    InMux I__6886 (
            .O(N__31644),
            .I(N__31639));
    LocalMux I__6885 (
            .O(N__31639),
            .I(\b2v_inst5.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__6884 (
            .O(N__31636),
            .I(\b2v_inst5.un2_count_1_axb_9_cascade_ ));
    InMux I__6883 (
            .O(N__31633),
            .I(N__31627));
    InMux I__6882 (
            .O(N__31632),
            .I(N__31627));
    LocalMux I__6881 (
            .O(N__31627),
            .I(\b2v_inst5.count_1_9 ));
    CascadeMux I__6880 (
            .O(N__31624),
            .I(N__31621));
    InMux I__6879 (
            .O(N__31621),
            .I(N__31618));
    LocalMux I__6878 (
            .O(N__31618),
            .I(\b2v_inst5.count_rst_5 ));
    InMux I__6877 (
            .O(N__31615),
            .I(N__31612));
    LocalMux I__6876 (
            .O(N__31612),
            .I(N__31609));
    Span4Mux_h I__6875 (
            .O(N__31609),
            .I(N__31606));
    Odrv4 I__6874 (
            .O(N__31606),
            .I(\b2v_inst5.un12_clk_100khz_6 ));
    CascadeMux I__6873 (
            .O(N__31603),
            .I(\b2v_inst5.count_rst_4_cascade_ ));
    CascadeMux I__6872 (
            .O(N__31600),
            .I(N__31596));
    InMux I__6871 (
            .O(N__31599),
            .I(N__31592));
    InMux I__6870 (
            .O(N__31596),
            .I(N__31587));
    InMux I__6869 (
            .O(N__31595),
            .I(N__31587));
    LocalMux I__6868 (
            .O(N__31592),
            .I(\b2v_inst5.countZ0Z_10 ));
    LocalMux I__6867 (
            .O(N__31587),
            .I(\b2v_inst5.countZ0Z_10 ));
    InMux I__6866 (
            .O(N__31582),
            .I(N__31576));
    InMux I__6865 (
            .O(N__31581),
            .I(N__31576));
    LocalMux I__6864 (
            .O(N__31576),
            .I(\b2v_inst5.un2_count_1_cry_9_THRU_CO ));
    CascadeMux I__6863 (
            .O(N__31573),
            .I(\b2v_inst5.countZ0Z_10_cascade_ ));
    InMux I__6862 (
            .O(N__31570),
            .I(N__31567));
    LocalMux I__6861 (
            .O(N__31567),
            .I(\b2v_inst5.count_1_10 ));
    CascadeMux I__6860 (
            .O(N__31564),
            .I(N__31561));
    InMux I__6859 (
            .O(N__31561),
            .I(N__31557));
    InMux I__6858 (
            .O(N__31560),
            .I(N__31552));
    LocalMux I__6857 (
            .O(N__31557),
            .I(N__31549));
    InMux I__6856 (
            .O(N__31556),
            .I(N__31543));
    InMux I__6855 (
            .O(N__31555),
            .I(N__31543));
    LocalMux I__6854 (
            .O(N__31552),
            .I(N__31540));
    Span4Mux_s3_h I__6853 (
            .O(N__31549),
            .I(N__31537));
    InMux I__6852 (
            .O(N__31548),
            .I(N__31534));
    LocalMux I__6851 (
            .O(N__31543),
            .I(\b2v_inst5.un2_count_1_cry_0 ));
    Odrv12 I__6850 (
            .O(N__31540),
            .I(\b2v_inst5.un2_count_1_cry_0 ));
    Odrv4 I__6849 (
            .O(N__31537),
            .I(\b2v_inst5.un2_count_1_cry_0 ));
    LocalMux I__6848 (
            .O(N__31534),
            .I(\b2v_inst5.un2_count_1_cry_0 ));
    InMux I__6847 (
            .O(N__31525),
            .I(N__31514));
    InMux I__6846 (
            .O(N__31524),
            .I(N__31511));
    InMux I__6845 (
            .O(N__31523),
            .I(N__31502));
    InMux I__6844 (
            .O(N__31522),
            .I(N__31502));
    InMux I__6843 (
            .O(N__31521),
            .I(N__31502));
    InMux I__6842 (
            .O(N__31520),
            .I(N__31502));
    InMux I__6841 (
            .O(N__31519),
            .I(N__31495));
    InMux I__6840 (
            .O(N__31518),
            .I(N__31495));
    InMux I__6839 (
            .O(N__31517),
            .I(N__31495));
    LocalMux I__6838 (
            .O(N__31514),
            .I(N__31488));
    LocalMux I__6837 (
            .O(N__31511),
            .I(N__31481));
    LocalMux I__6836 (
            .O(N__31502),
            .I(N__31481));
    LocalMux I__6835 (
            .O(N__31495),
            .I(N__31481));
    InMux I__6834 (
            .O(N__31494),
            .I(N__31478));
    InMux I__6833 (
            .O(N__31493),
            .I(N__31471));
    InMux I__6832 (
            .O(N__31492),
            .I(N__31471));
    InMux I__6831 (
            .O(N__31491),
            .I(N__31471));
    Span4Mux_s3_h I__6830 (
            .O(N__31488),
            .I(N__31466));
    Span4Mux_s3_h I__6829 (
            .O(N__31481),
            .I(N__31466));
    LocalMux I__6828 (
            .O(N__31478),
            .I(\b2v_inst5.N_1_i ));
    LocalMux I__6827 (
            .O(N__31471),
            .I(\b2v_inst5.N_1_i ));
    Odrv4 I__6826 (
            .O(N__31466),
            .I(\b2v_inst5.N_1_i ));
    InMux I__6825 (
            .O(N__31459),
            .I(N__31456));
    LocalMux I__6824 (
            .O(N__31456),
            .I(N__31453));
    Odrv4 I__6823 (
            .O(N__31453),
            .I(\b2v_inst5.count_1_0 ));
    InMux I__6822 (
            .O(N__31450),
            .I(bfn_11_4_0_));
    InMux I__6821 (
            .O(N__31447),
            .I(\b2v_inst5.un2_count_1_cry_9 ));
    InMux I__6820 (
            .O(N__31444),
            .I(N__31440));
    InMux I__6819 (
            .O(N__31443),
            .I(N__31437));
    LocalMux I__6818 (
            .O(N__31440),
            .I(N__31432));
    LocalMux I__6817 (
            .O(N__31437),
            .I(N__31432));
    Odrv12 I__6816 (
            .O(N__31432),
            .I(\b2v_inst5.count_rst_3 ));
    InMux I__6815 (
            .O(N__31429),
            .I(\b2v_inst5.un2_count_1_cry_10 ));
    InMux I__6814 (
            .O(N__31426),
            .I(N__31422));
    InMux I__6813 (
            .O(N__31425),
            .I(N__31419));
    LocalMux I__6812 (
            .O(N__31422),
            .I(N__31416));
    LocalMux I__6811 (
            .O(N__31419),
            .I(\b2v_inst5.countZ0Z_12 ));
    Odrv4 I__6810 (
            .O(N__31416),
            .I(\b2v_inst5.countZ0Z_12 ));
    InMux I__6809 (
            .O(N__31411),
            .I(N__31407));
    InMux I__6808 (
            .O(N__31410),
            .I(N__31404));
    LocalMux I__6807 (
            .O(N__31407),
            .I(N__31401));
    LocalMux I__6806 (
            .O(N__31404),
            .I(N__31398));
    Odrv12 I__6805 (
            .O(N__31401),
            .I(\b2v_inst5.count_rst_2 ));
    Odrv4 I__6804 (
            .O(N__31398),
            .I(\b2v_inst5.count_rst_2 ));
    InMux I__6803 (
            .O(N__31393),
            .I(\b2v_inst5.un2_count_1_cry_11 ));
    InMux I__6802 (
            .O(N__31390),
            .I(N__31387));
    LocalMux I__6801 (
            .O(N__31387),
            .I(N__31383));
    InMux I__6800 (
            .O(N__31386),
            .I(N__31380));
    Span4Mux_s2_h I__6799 (
            .O(N__31383),
            .I(N__31377));
    LocalMux I__6798 (
            .O(N__31380),
            .I(\b2v_inst5.un2_count_1_axb_13 ));
    Odrv4 I__6797 (
            .O(N__31377),
            .I(\b2v_inst5.un2_count_1_axb_13 ));
    CascadeMux I__6796 (
            .O(N__31372),
            .I(N__31368));
    InMux I__6795 (
            .O(N__31371),
            .I(N__31365));
    InMux I__6794 (
            .O(N__31368),
            .I(N__31362));
    LocalMux I__6793 (
            .O(N__31365),
            .I(N__31357));
    LocalMux I__6792 (
            .O(N__31362),
            .I(N__31357));
    Span4Mux_v I__6791 (
            .O(N__31357),
            .I(N__31354));
    Span4Mux_h I__6790 (
            .O(N__31354),
            .I(N__31351));
    Odrv4 I__6789 (
            .O(N__31351),
            .I(\b2v_inst5.un2_count_1_cry_12_THRU_CO ));
    InMux I__6788 (
            .O(N__31348),
            .I(\b2v_inst5.un2_count_1_cry_12 ));
    CascadeMux I__6787 (
            .O(N__31345),
            .I(N__31342));
    InMux I__6786 (
            .O(N__31342),
            .I(N__31338));
    InMux I__6785 (
            .O(N__31341),
            .I(N__31335));
    LocalMux I__6784 (
            .O(N__31338),
            .I(N__31332));
    LocalMux I__6783 (
            .O(N__31335),
            .I(N__31329));
    Odrv4 I__6782 (
            .O(N__31332),
            .I(\b2v_inst5.countZ0Z_14 ));
    Odrv4 I__6781 (
            .O(N__31329),
            .I(\b2v_inst5.countZ0Z_14 ));
    InMux I__6780 (
            .O(N__31324),
            .I(N__31320));
    InMux I__6779 (
            .O(N__31323),
            .I(N__31317));
    LocalMux I__6778 (
            .O(N__31320),
            .I(N__31312));
    LocalMux I__6777 (
            .O(N__31317),
            .I(N__31312));
    Span4Mux_h I__6776 (
            .O(N__31312),
            .I(N__31309));
    Odrv4 I__6775 (
            .O(N__31309),
            .I(\b2v_inst5.count_rst_0 ));
    InMux I__6774 (
            .O(N__31306),
            .I(\b2v_inst5.un2_count_1_cry_13 ));
    InMux I__6773 (
            .O(N__31303),
            .I(N__31300));
    LocalMux I__6772 (
            .O(N__31300),
            .I(N__31296));
    InMux I__6771 (
            .O(N__31299),
            .I(N__31293));
    Odrv12 I__6770 (
            .O(N__31296),
            .I(\b2v_inst5.countZ0Z_15 ));
    LocalMux I__6769 (
            .O(N__31293),
            .I(\b2v_inst5.countZ0Z_15 ));
    InMux I__6768 (
            .O(N__31288),
            .I(\b2v_inst5.un2_count_1_cry_14 ));
    InMux I__6767 (
            .O(N__31285),
            .I(N__31282));
    LocalMux I__6766 (
            .O(N__31282),
            .I(N__31279));
    Span4Mux_h I__6765 (
            .O(N__31279),
            .I(N__31275));
    InMux I__6764 (
            .O(N__31278),
            .I(N__31272));
    Odrv4 I__6763 (
            .O(N__31275),
            .I(\b2v_inst5.count_rst ));
    LocalMux I__6762 (
            .O(N__31272),
            .I(\b2v_inst5.count_rst ));
    InMux I__6761 (
            .O(N__31267),
            .I(N__31264));
    LocalMux I__6760 (
            .O(N__31264),
            .I(N__31261));
    Span4Mux_h I__6759 (
            .O(N__31261),
            .I(N__31258));
    Odrv4 I__6758 (
            .O(N__31258),
            .I(\b2v_inst5.count_1_15 ));
    InMux I__6757 (
            .O(N__31255),
            .I(N__31252));
    LocalMux I__6756 (
            .O(N__31252),
            .I(N__31247));
    InMux I__6755 (
            .O(N__31251),
            .I(N__31244));
    InMux I__6754 (
            .O(N__31250),
            .I(N__31241));
    Span4Mux_s2_h I__6753 (
            .O(N__31247),
            .I(N__31238));
    LocalMux I__6752 (
            .O(N__31244),
            .I(\b2v_inst5.countZ0Z_1 ));
    LocalMux I__6751 (
            .O(N__31241),
            .I(\b2v_inst5.countZ0Z_1 ));
    Odrv4 I__6750 (
            .O(N__31238),
            .I(\b2v_inst5.countZ0Z_1 ));
    InMux I__6749 (
            .O(N__31231),
            .I(N__31228));
    LocalMux I__6748 (
            .O(N__31228),
            .I(N__31225));
    Span4Mux_s3_v I__6747 (
            .O(N__31225),
            .I(N__31222));
    Odrv4 I__6746 (
            .O(N__31222),
            .I(\b2v_inst5.un2_count_1_axb_2 ));
    CascadeMux I__6745 (
            .O(N__31219),
            .I(N__31216));
    InMux I__6744 (
            .O(N__31216),
            .I(N__31207));
    InMux I__6743 (
            .O(N__31215),
            .I(N__31207));
    InMux I__6742 (
            .O(N__31214),
            .I(N__31207));
    LocalMux I__6741 (
            .O(N__31207),
            .I(N__31204));
    Span4Mux_h I__6740 (
            .O(N__31204),
            .I(N__31201));
    Odrv4 I__6739 (
            .O(N__31201),
            .I(\b2v_inst5.count_rst_12 ));
    InMux I__6738 (
            .O(N__31198),
            .I(\b2v_inst5.un2_count_1_cry_1 ));
    InMux I__6737 (
            .O(N__31195),
            .I(N__31192));
    LocalMux I__6736 (
            .O(N__31192),
            .I(N__31188));
    InMux I__6735 (
            .O(N__31191),
            .I(N__31185));
    Span4Mux_s2_h I__6734 (
            .O(N__31188),
            .I(N__31182));
    LocalMux I__6733 (
            .O(N__31185),
            .I(\b2v_inst5.countZ0Z_3 ));
    Odrv4 I__6732 (
            .O(N__31182),
            .I(\b2v_inst5.countZ0Z_3 ));
    CascadeMux I__6731 (
            .O(N__31177),
            .I(N__31173));
    InMux I__6730 (
            .O(N__31176),
            .I(N__31168));
    InMux I__6729 (
            .O(N__31173),
            .I(N__31168));
    LocalMux I__6728 (
            .O(N__31168),
            .I(N__31165));
    Span4Mux_h I__6727 (
            .O(N__31165),
            .I(N__31162));
    Odrv4 I__6726 (
            .O(N__31162),
            .I(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ));
    InMux I__6725 (
            .O(N__31159),
            .I(\b2v_inst5.un2_count_1_cry_2 ));
    InMux I__6724 (
            .O(N__31156),
            .I(N__31153));
    LocalMux I__6723 (
            .O(N__31153),
            .I(N__31149));
    CascadeMux I__6722 (
            .O(N__31152),
            .I(N__31146));
    Span4Mux_h I__6721 (
            .O(N__31149),
            .I(N__31143));
    InMux I__6720 (
            .O(N__31146),
            .I(N__31140));
    Span4Mux_v I__6719 (
            .O(N__31143),
            .I(N__31137));
    LocalMux I__6718 (
            .O(N__31140),
            .I(\b2v_inst5.un2_count_1_axb_4 ));
    Odrv4 I__6717 (
            .O(N__31137),
            .I(\b2v_inst5.un2_count_1_axb_4 ));
    InMux I__6716 (
            .O(N__31132),
            .I(N__31126));
    InMux I__6715 (
            .O(N__31131),
            .I(N__31126));
    LocalMux I__6714 (
            .O(N__31126),
            .I(N__31123));
    Span4Mux_v I__6713 (
            .O(N__31123),
            .I(N__31120));
    Span4Mux_h I__6712 (
            .O(N__31120),
            .I(N__31117));
    Odrv4 I__6711 (
            .O(N__31117),
            .I(\b2v_inst5.un2_count_1_cry_3_THRU_CO ));
    InMux I__6710 (
            .O(N__31114),
            .I(\b2v_inst5.un2_count_1_cry_3 ));
    InMux I__6709 (
            .O(N__31111),
            .I(\b2v_inst5.un2_count_1_cry_4 ));
    InMux I__6708 (
            .O(N__31108),
            .I(\b2v_inst5.un2_count_1_cry_5 ));
    InMux I__6707 (
            .O(N__31105),
            .I(\b2v_inst5.un2_count_1_cry_6 ));
    CascadeMux I__6706 (
            .O(N__31102),
            .I(N__31098));
    InMux I__6705 (
            .O(N__31101),
            .I(N__31095));
    InMux I__6704 (
            .O(N__31098),
            .I(N__31092));
    LocalMux I__6703 (
            .O(N__31095),
            .I(N__31089));
    LocalMux I__6702 (
            .O(N__31092),
            .I(N__31086));
    Span4Mux_s3_v I__6701 (
            .O(N__31089),
            .I(N__31082));
    Span4Mux_v I__6700 (
            .O(N__31086),
            .I(N__31079));
    InMux I__6699 (
            .O(N__31085),
            .I(N__31076));
    Span4Mux_h I__6698 (
            .O(N__31082),
            .I(N__31073));
    Odrv4 I__6697 (
            .O(N__31079),
            .I(\b2v_inst5.countZ0Z_8 ));
    LocalMux I__6696 (
            .O(N__31076),
            .I(\b2v_inst5.countZ0Z_8 ));
    Odrv4 I__6695 (
            .O(N__31073),
            .I(\b2v_inst5.countZ0Z_8 ));
    CascadeMux I__6694 (
            .O(N__31066),
            .I(N__31063));
    InMux I__6693 (
            .O(N__31063),
            .I(N__31060));
    LocalMux I__6692 (
            .O(N__31060),
            .I(N__31056));
    InMux I__6691 (
            .O(N__31059),
            .I(N__31053));
    Span4Mux_v I__6690 (
            .O(N__31056),
            .I(N__31048));
    LocalMux I__6689 (
            .O(N__31053),
            .I(N__31048));
    Span4Mux_h I__6688 (
            .O(N__31048),
            .I(N__31045));
    Odrv4 I__6687 (
            .O(N__31045),
            .I(\b2v_inst5.un2_count_1_cry_7_THRU_CO ));
    InMux I__6686 (
            .O(N__31042),
            .I(\b2v_inst5.un2_count_1_cry_7 ));
    InMux I__6685 (
            .O(N__31039),
            .I(N__31033));
    InMux I__6684 (
            .O(N__31038),
            .I(N__31033));
    LocalMux I__6683 (
            .O(N__31033),
            .I(N__31030));
    Span4Mux_s2_h I__6682 (
            .O(N__31030),
            .I(N__31027));
    Odrv4 I__6681 (
            .O(N__31027),
            .I(\b2v_inst36.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__6680 (
            .O(N__31024),
            .I(\b2v_inst36.countZ0Z_5_cascade_ ));
    InMux I__6679 (
            .O(N__31021),
            .I(N__31018));
    LocalMux I__6678 (
            .O(N__31018),
            .I(\b2v_inst36.count_2_5 ));
    InMux I__6677 (
            .O(N__31015),
            .I(N__31010));
    InMux I__6676 (
            .O(N__31014),
            .I(N__31005));
    InMux I__6675 (
            .O(N__31013),
            .I(N__31005));
    LocalMux I__6674 (
            .O(N__31010),
            .I(N__30999));
    LocalMux I__6673 (
            .O(N__31005),
            .I(N__30999));
    InMux I__6672 (
            .O(N__31004),
            .I(N__30996));
    Span4Mux_s3_h I__6671 (
            .O(N__30999),
            .I(N__30993));
    LocalMux I__6670 (
            .O(N__30996),
            .I(\b2v_inst36.countZ0Z_7 ));
    Odrv4 I__6669 (
            .O(N__30993),
            .I(\b2v_inst36.countZ0Z_7 ));
    CascadeMux I__6668 (
            .O(N__30988),
            .I(N__30982));
    InMux I__6667 (
            .O(N__30987),
            .I(N__30970));
    InMux I__6666 (
            .O(N__30986),
            .I(N__30961));
    InMux I__6665 (
            .O(N__30985),
            .I(N__30961));
    InMux I__6664 (
            .O(N__30982),
            .I(N__30961));
    InMux I__6663 (
            .O(N__30981),
            .I(N__30961));
    CascadeMux I__6662 (
            .O(N__30980),
            .I(N__30953));
    InMux I__6661 (
            .O(N__30979),
            .I(N__30945));
    InMux I__6660 (
            .O(N__30978),
            .I(N__30945));
    InMux I__6659 (
            .O(N__30977),
            .I(N__30938));
    InMux I__6658 (
            .O(N__30976),
            .I(N__30938));
    InMux I__6657 (
            .O(N__30975),
            .I(N__30938));
    InMux I__6656 (
            .O(N__30974),
            .I(N__30933));
    InMux I__6655 (
            .O(N__30973),
            .I(N__30933));
    LocalMux I__6654 (
            .O(N__30970),
            .I(N__30928));
    LocalMux I__6653 (
            .O(N__30961),
            .I(N__30928));
    CascadeMux I__6652 (
            .O(N__30960),
            .I(N__30924));
    InMux I__6651 (
            .O(N__30959),
            .I(N__30917));
    InMux I__6650 (
            .O(N__30958),
            .I(N__30917));
    InMux I__6649 (
            .O(N__30957),
            .I(N__30917));
    CascadeMux I__6648 (
            .O(N__30956),
            .I(N__30913));
    InMux I__6647 (
            .O(N__30953),
            .I(N__30909));
    InMux I__6646 (
            .O(N__30952),
            .I(N__30902));
    InMux I__6645 (
            .O(N__30951),
            .I(N__30902));
    InMux I__6644 (
            .O(N__30950),
            .I(N__30902));
    LocalMux I__6643 (
            .O(N__30945),
            .I(N__30899));
    LocalMux I__6642 (
            .O(N__30938),
            .I(N__30892));
    LocalMux I__6641 (
            .O(N__30933),
            .I(N__30892));
    Span4Mux_s3_h I__6640 (
            .O(N__30928),
            .I(N__30892));
    InMux I__6639 (
            .O(N__30927),
            .I(N__30887));
    InMux I__6638 (
            .O(N__30924),
            .I(N__30887));
    LocalMux I__6637 (
            .O(N__30917),
            .I(N__30884));
    InMux I__6636 (
            .O(N__30916),
            .I(N__30877));
    InMux I__6635 (
            .O(N__30913),
            .I(N__30877));
    InMux I__6634 (
            .O(N__30912),
            .I(N__30877));
    LocalMux I__6633 (
            .O(N__30909),
            .I(\b2v_inst36.N_2942_i ));
    LocalMux I__6632 (
            .O(N__30902),
            .I(\b2v_inst36.N_2942_i ));
    Odrv4 I__6631 (
            .O(N__30899),
            .I(\b2v_inst36.N_2942_i ));
    Odrv4 I__6630 (
            .O(N__30892),
            .I(\b2v_inst36.N_2942_i ));
    LocalMux I__6629 (
            .O(N__30887),
            .I(\b2v_inst36.N_2942_i ));
    Odrv4 I__6628 (
            .O(N__30884),
            .I(\b2v_inst36.N_2942_i ));
    LocalMux I__6627 (
            .O(N__30877),
            .I(\b2v_inst36.N_2942_i ));
    CascadeMux I__6626 (
            .O(N__30862),
            .I(N__30849));
    CascadeMux I__6625 (
            .O(N__30861),
            .I(N__30846));
    InMux I__6624 (
            .O(N__30860),
            .I(N__30835));
    InMux I__6623 (
            .O(N__30859),
            .I(N__30835));
    InMux I__6622 (
            .O(N__30858),
            .I(N__30835));
    InMux I__6621 (
            .O(N__30857),
            .I(N__30828));
    InMux I__6620 (
            .O(N__30856),
            .I(N__30828));
    InMux I__6619 (
            .O(N__30855),
            .I(N__30828));
    InMux I__6618 (
            .O(N__30854),
            .I(N__30821));
    InMux I__6617 (
            .O(N__30853),
            .I(N__30821));
    InMux I__6616 (
            .O(N__30852),
            .I(N__30821));
    InMux I__6615 (
            .O(N__30849),
            .I(N__30816));
    InMux I__6614 (
            .O(N__30846),
            .I(N__30816));
    InMux I__6613 (
            .O(N__30845),
            .I(N__30804));
    InMux I__6612 (
            .O(N__30844),
            .I(N__30804));
    InMux I__6611 (
            .O(N__30843),
            .I(N__30804));
    InMux I__6610 (
            .O(N__30842),
            .I(N__30801));
    LocalMux I__6609 (
            .O(N__30835),
            .I(N__30796));
    LocalMux I__6608 (
            .O(N__30828),
            .I(N__30796));
    LocalMux I__6607 (
            .O(N__30821),
            .I(N__30791));
    LocalMux I__6606 (
            .O(N__30816),
            .I(N__30791));
    InMux I__6605 (
            .O(N__30815),
            .I(N__30780));
    InMux I__6604 (
            .O(N__30814),
            .I(N__30780));
    InMux I__6603 (
            .O(N__30813),
            .I(N__30780));
    InMux I__6602 (
            .O(N__30812),
            .I(N__30780));
    InMux I__6601 (
            .O(N__30811),
            .I(N__30780));
    LocalMux I__6600 (
            .O(N__30804),
            .I(N__30777));
    LocalMux I__6599 (
            .O(N__30801),
            .I(\b2v_inst36.N_1_i ));
    Odrv4 I__6598 (
            .O(N__30796),
            .I(\b2v_inst36.N_1_i ));
    Odrv12 I__6597 (
            .O(N__30791),
            .I(\b2v_inst36.N_1_i ));
    LocalMux I__6596 (
            .O(N__30780),
            .I(\b2v_inst36.N_1_i ));
    Odrv4 I__6595 (
            .O(N__30777),
            .I(\b2v_inst36.N_1_i ));
    InMux I__6594 (
            .O(N__30766),
            .I(N__30762));
    InMux I__6593 (
            .O(N__30765),
            .I(N__30759));
    LocalMux I__6592 (
            .O(N__30762),
            .I(N__30756));
    LocalMux I__6591 (
            .O(N__30759),
            .I(N__30753));
    Span4Mux_s1_h I__6590 (
            .O(N__30756),
            .I(N__30750));
    Odrv4 I__6589 (
            .O(N__30753),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    Odrv4 I__6588 (
            .O(N__30750),
            .I(\b2v_inst36.un2_count_1_cry_6_THRU_CO ));
    InMux I__6587 (
            .O(N__30745),
            .I(N__30742));
    LocalMux I__6586 (
            .O(N__30742),
            .I(N__30739));
    Span4Mux_h I__6585 (
            .O(N__30739),
            .I(N__30736));
    Odrv4 I__6584 (
            .O(N__30736),
            .I(\b2v_inst36.count_2_7 ));
    CEMux I__6583 (
            .O(N__30733),
            .I(N__30727));
    CEMux I__6582 (
            .O(N__30732),
            .I(N__30721));
    CEMux I__6581 (
            .O(N__30731),
            .I(N__30718));
    CEMux I__6580 (
            .O(N__30730),
            .I(N__30715));
    LocalMux I__6579 (
            .O(N__30727),
            .I(N__30712));
    InMux I__6578 (
            .O(N__30726),
            .I(N__30702));
    InMux I__6577 (
            .O(N__30725),
            .I(N__30702));
    InMux I__6576 (
            .O(N__30724),
            .I(N__30690));
    LocalMux I__6575 (
            .O(N__30721),
            .I(N__30687));
    LocalMux I__6574 (
            .O(N__30718),
            .I(N__30684));
    LocalMux I__6573 (
            .O(N__30715),
            .I(N__30681));
    IoSpan4Mux I__6572 (
            .O(N__30712),
            .I(N__30677));
    InMux I__6571 (
            .O(N__30711),
            .I(N__30672));
    CEMux I__6570 (
            .O(N__30710),
            .I(N__30672));
    InMux I__6569 (
            .O(N__30709),
            .I(N__30665));
    InMux I__6568 (
            .O(N__30708),
            .I(N__30665));
    InMux I__6567 (
            .O(N__30707),
            .I(N__30665));
    LocalMux I__6566 (
            .O(N__30702),
            .I(N__30662));
    InMux I__6565 (
            .O(N__30701),
            .I(N__30655));
    CEMux I__6564 (
            .O(N__30700),
            .I(N__30655));
    CEMux I__6563 (
            .O(N__30699),
            .I(N__30644));
    InMux I__6562 (
            .O(N__30698),
            .I(N__30644));
    InMux I__6561 (
            .O(N__30697),
            .I(N__30644));
    InMux I__6560 (
            .O(N__30696),
            .I(N__30644));
    InMux I__6559 (
            .O(N__30695),
            .I(N__30644));
    InMux I__6558 (
            .O(N__30694),
            .I(N__30639));
    InMux I__6557 (
            .O(N__30693),
            .I(N__30639));
    LocalMux I__6556 (
            .O(N__30690),
            .I(N__30634));
    Span4Mux_s2_v I__6555 (
            .O(N__30687),
            .I(N__30634));
    Span4Mux_s2_v I__6554 (
            .O(N__30684),
            .I(N__30629));
    Span4Mux_s2_v I__6553 (
            .O(N__30681),
            .I(N__30629));
    InMux I__6552 (
            .O(N__30680),
            .I(N__30626));
    Span4Mux_s0_v I__6551 (
            .O(N__30677),
            .I(N__30617));
    LocalMux I__6550 (
            .O(N__30672),
            .I(N__30617));
    LocalMux I__6549 (
            .O(N__30665),
            .I(N__30617));
    Span4Mux_s3_h I__6548 (
            .O(N__30662),
            .I(N__30617));
    InMux I__6547 (
            .O(N__30661),
            .I(N__30612));
    InMux I__6546 (
            .O(N__30660),
            .I(N__30612));
    LocalMux I__6545 (
            .O(N__30655),
            .I(N__30605));
    LocalMux I__6544 (
            .O(N__30644),
            .I(N__30605));
    LocalMux I__6543 (
            .O(N__30639),
            .I(N__30605));
    Odrv4 I__6542 (
            .O(N__30634),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__6541 (
            .O(N__30629),
            .I(\b2v_inst36.count_en ));
    LocalMux I__6540 (
            .O(N__30626),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__6539 (
            .O(N__30617),
            .I(\b2v_inst36.count_en ));
    LocalMux I__6538 (
            .O(N__30612),
            .I(\b2v_inst36.count_en ));
    Odrv4 I__6537 (
            .O(N__30605),
            .I(\b2v_inst36.count_en ));
    SRMux I__6536 (
            .O(N__30592),
            .I(N__30584));
    SRMux I__6535 (
            .O(N__30591),
            .I(N__30581));
    SRMux I__6534 (
            .O(N__30590),
            .I(N__30577));
    SRMux I__6533 (
            .O(N__30589),
            .I(N__30574));
    SRMux I__6532 (
            .O(N__30588),
            .I(N__30571));
    SRMux I__6531 (
            .O(N__30587),
            .I(N__30568));
    LocalMux I__6530 (
            .O(N__30584),
            .I(N__30565));
    LocalMux I__6529 (
            .O(N__30581),
            .I(N__30562));
    SRMux I__6528 (
            .O(N__30580),
            .I(N__30559));
    LocalMux I__6527 (
            .O(N__30577),
            .I(N__30556));
    LocalMux I__6526 (
            .O(N__30574),
            .I(N__30553));
    LocalMux I__6525 (
            .O(N__30571),
            .I(N__30550));
    LocalMux I__6524 (
            .O(N__30568),
            .I(N__30547));
    Span4Mux_s2_v I__6523 (
            .O(N__30565),
            .I(N__30540));
    Span4Mux_s2_v I__6522 (
            .O(N__30562),
            .I(N__30540));
    LocalMux I__6521 (
            .O(N__30559),
            .I(N__30540));
    Span4Mux_s3_v I__6520 (
            .O(N__30556),
            .I(N__30537));
    Span4Mux_s2_v I__6519 (
            .O(N__30553),
            .I(N__30532));
    Span4Mux_h I__6518 (
            .O(N__30550),
            .I(N__30527));
    Span4Mux_h I__6517 (
            .O(N__30547),
            .I(N__30527));
    Span4Mux_h I__6516 (
            .O(N__30540),
            .I(N__30524));
    Span4Mux_v I__6515 (
            .O(N__30537),
            .I(N__30521));
    InMux I__6514 (
            .O(N__30536),
            .I(N__30516));
    InMux I__6513 (
            .O(N__30535),
            .I(N__30516));
    Odrv4 I__6512 (
            .O(N__30532),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__6511 (
            .O(N__30527),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__6510 (
            .O(N__30524),
            .I(\b2v_inst36.count_0_sqmuxa ));
    Odrv4 I__6509 (
            .O(N__30521),
            .I(\b2v_inst36.count_0_sqmuxa ));
    LocalMux I__6508 (
            .O(N__30516),
            .I(\b2v_inst36.count_0_sqmuxa ));
    InMux I__6507 (
            .O(N__30505),
            .I(N__30502));
    LocalMux I__6506 (
            .O(N__30502),
            .I(\b2v_inst6.count_0_14 ));
    CascadeMux I__6505 (
            .O(N__30499),
            .I(\b2v_inst6.countZ0Z_14_cascade_ ));
    InMux I__6504 (
            .O(N__30496),
            .I(N__30493));
    LocalMux I__6503 (
            .O(N__30493),
            .I(\b2v_inst6.count_0_6 ));
    CascadeMux I__6502 (
            .O(N__30490),
            .I(N__30485));
    CascadeMux I__6501 (
            .O(N__30489),
            .I(N__30482));
    CascadeMux I__6500 (
            .O(N__30488),
            .I(N__30479));
    InMux I__6499 (
            .O(N__30485),
            .I(N__30476));
    InMux I__6498 (
            .O(N__30482),
            .I(N__30471));
    InMux I__6497 (
            .O(N__30479),
            .I(N__30471));
    LocalMux I__6496 (
            .O(N__30476),
            .I(\b2v_inst11.mult1_un152_sum_i_0_8 ));
    LocalMux I__6495 (
            .O(N__30471),
            .I(\b2v_inst11.mult1_un152_sum_i_0_8 ));
    InMux I__6494 (
            .O(N__30466),
            .I(N__30463));
    LocalMux I__6493 (
            .O(N__30463),
            .I(N__30460));
    Span4Mux_s2_v I__6492 (
            .O(N__30460),
            .I(N__30457));
    Odrv4 I__6491 (
            .O(N__30457),
            .I(\b2v_inst5.N_51 ));
    InMux I__6490 (
            .O(N__30454),
            .I(N__30451));
    LocalMux I__6489 (
            .O(N__30451),
            .I(N__30448));
    Span4Mux_h I__6488 (
            .O(N__30448),
            .I(N__30445));
    Odrv4 I__6487 (
            .O(N__30445),
            .I(\b2v_inst5.curr_state_0_1 ));
    IoInMux I__6486 (
            .O(N__30442),
            .I(N__30439));
    LocalMux I__6485 (
            .O(N__30439),
            .I(N__30433));
    InMux I__6484 (
            .O(N__30438),
            .I(N__30430));
    InMux I__6483 (
            .O(N__30437),
            .I(N__30427));
    InMux I__6482 (
            .O(N__30436),
            .I(N__30424));
    Span12Mux_s0_v I__6481 (
            .O(N__30433),
            .I(N__30421));
    LocalMux I__6480 (
            .O(N__30430),
            .I(N__30416));
    LocalMux I__6479 (
            .O(N__30427),
            .I(N__30416));
    LocalMux I__6478 (
            .O(N__30424),
            .I(N__30413));
    Odrv12 I__6477 (
            .O(N__30421),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6476 (
            .O(N__30416),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6475 (
            .O(N__30413),
            .I(CONSTANT_ONE_NET));
    InMux I__6474 (
            .O(N__30406),
            .I(N__30403));
    LocalMux I__6473 (
            .O(N__30403),
            .I(N__30400));
    Span4Mux_s1_v I__6472 (
            .O(N__30400),
            .I(N__30395));
    InMux I__6471 (
            .O(N__30399),
            .I(N__30392));
    InMux I__6470 (
            .O(N__30398),
            .I(N__30389));
    Odrv4 I__6469 (
            .O(N__30395),
            .I(\b2v_inst36.countZ0Z_2 ));
    LocalMux I__6468 (
            .O(N__30392),
            .I(\b2v_inst36.countZ0Z_2 ));
    LocalMux I__6467 (
            .O(N__30389),
            .I(\b2v_inst36.countZ0Z_2 ));
    InMux I__6466 (
            .O(N__30382),
            .I(N__30379));
    LocalMux I__6465 (
            .O(N__30379),
            .I(N__30376));
    Span4Mux_h I__6464 (
            .O(N__30376),
            .I(N__30373));
    Odrv4 I__6463 (
            .O(N__30373),
            .I(\b2v_inst36.un12_clk_100khz_11 ));
    CascadeMux I__6462 (
            .O(N__30370),
            .I(\b2v_inst36.count_rst_11_cascade_ ));
    InMux I__6461 (
            .O(N__30367),
            .I(N__30360));
    InMux I__6460 (
            .O(N__30366),
            .I(N__30360));
    InMux I__6459 (
            .O(N__30365),
            .I(N__30357));
    LocalMux I__6458 (
            .O(N__30360),
            .I(N__30352));
    LocalMux I__6457 (
            .O(N__30357),
            .I(N__30352));
    Odrv4 I__6456 (
            .O(N__30352),
            .I(\b2v_inst36.countZ0Z_3 ));
    InMux I__6455 (
            .O(N__30349),
            .I(N__30343));
    InMux I__6454 (
            .O(N__30348),
            .I(N__30343));
    LocalMux I__6453 (
            .O(N__30343),
            .I(N__30340));
    Odrv4 I__6452 (
            .O(N__30340),
            .I(\b2v_inst36.un2_count_1_cry_2_THRU_CO ));
    CascadeMux I__6451 (
            .O(N__30337),
            .I(\b2v_inst36.countZ0Z_3_cascade_ ));
    InMux I__6450 (
            .O(N__30334),
            .I(N__30331));
    LocalMux I__6449 (
            .O(N__30331),
            .I(\b2v_inst36.count_2_3 ));
    CascadeMux I__6448 (
            .O(N__30328),
            .I(\b2v_inst36.count_rst_9_cascade_ ));
    CascadeMux I__6447 (
            .O(N__30325),
            .I(N__30322));
    InMux I__6446 (
            .O(N__30322),
            .I(N__30317));
    InMux I__6445 (
            .O(N__30321),
            .I(N__30314));
    InMux I__6444 (
            .O(N__30320),
            .I(N__30311));
    LocalMux I__6443 (
            .O(N__30317),
            .I(N__30308));
    LocalMux I__6442 (
            .O(N__30314),
            .I(N__30305));
    LocalMux I__6441 (
            .O(N__30311),
            .I(\b2v_inst36.countZ0Z_5 ));
    Odrv4 I__6440 (
            .O(N__30308),
            .I(\b2v_inst36.countZ0Z_5 ));
    Odrv4 I__6439 (
            .O(N__30305),
            .I(\b2v_inst36.countZ0Z_5 ));
    InMux I__6438 (
            .O(N__30298),
            .I(N__30292));
    CascadeMux I__6437 (
            .O(N__30297),
            .I(N__30288));
    CascadeMux I__6436 (
            .O(N__30296),
            .I(N__30284));
    InMux I__6435 (
            .O(N__30295),
            .I(N__30280));
    LocalMux I__6434 (
            .O(N__30292),
            .I(N__30275));
    InMux I__6433 (
            .O(N__30291),
            .I(N__30272));
    InMux I__6432 (
            .O(N__30288),
            .I(N__30269));
    InMux I__6431 (
            .O(N__30287),
            .I(N__30266));
    InMux I__6430 (
            .O(N__30284),
            .I(N__30261));
    InMux I__6429 (
            .O(N__30283),
            .I(N__30261));
    LocalMux I__6428 (
            .O(N__30280),
            .I(N__30258));
    InMux I__6427 (
            .O(N__30279),
            .I(N__30255));
    CascadeMux I__6426 (
            .O(N__30278),
            .I(N__30252));
    Span4Mux_h I__6425 (
            .O(N__30275),
            .I(N__30249));
    LocalMux I__6424 (
            .O(N__30272),
            .I(N__30246));
    LocalMux I__6423 (
            .O(N__30269),
            .I(N__30243));
    LocalMux I__6422 (
            .O(N__30266),
            .I(N__30238));
    LocalMux I__6421 (
            .O(N__30261),
            .I(N__30235));
    Span4Mux_s2_h I__6420 (
            .O(N__30258),
            .I(N__30230));
    LocalMux I__6419 (
            .O(N__30255),
            .I(N__30230));
    InMux I__6418 (
            .O(N__30252),
            .I(N__30227));
    Span4Mux_v I__6417 (
            .O(N__30249),
            .I(N__30224));
    Span4Mux_v I__6416 (
            .O(N__30246),
            .I(N__30219));
    Span4Mux_v I__6415 (
            .O(N__30243),
            .I(N__30219));
    InMux I__6414 (
            .O(N__30242),
            .I(N__30216));
    InMux I__6413 (
            .O(N__30241),
            .I(N__30213));
    Span4Mux_v I__6412 (
            .O(N__30238),
            .I(N__30206));
    Span4Mux_h I__6411 (
            .O(N__30235),
            .I(N__30206));
    Span4Mux_h I__6410 (
            .O(N__30230),
            .I(N__30206));
    LocalMux I__6409 (
            .O(N__30227),
            .I(N__30203));
    Odrv4 I__6408 (
            .O(N__30224),
            .I(dutycycle_RNIU8G3G_0_2));
    Odrv4 I__6407 (
            .O(N__30219),
            .I(dutycycle_RNIU8G3G_0_2));
    LocalMux I__6406 (
            .O(N__30216),
            .I(dutycycle_RNIU8G3G_0_2));
    LocalMux I__6405 (
            .O(N__30213),
            .I(dutycycle_RNIU8G3G_0_2));
    Odrv4 I__6404 (
            .O(N__30206),
            .I(dutycycle_RNIU8G3G_0_2));
    Odrv4 I__6403 (
            .O(N__30203),
            .I(dutycycle_RNIU8G3G_0_2));
    InMux I__6402 (
            .O(N__30190),
            .I(N__30187));
    LocalMux I__6401 (
            .O(N__30187),
            .I(\b2v_inst11.mult1_un152_sum_i ));
    InMux I__6400 (
            .O(N__30184),
            .I(\b2v_inst11.mult1_un159_sum_cry_1 ));
    InMux I__6399 (
            .O(N__30181),
            .I(N__30178));
    LocalMux I__6398 (
            .O(N__30178),
            .I(N__30175));
    Span12Mux_s6_h I__6397 (
            .O(N__30175),
            .I(N__30172));
    Odrv12 I__6396 (
            .O(N__30172),
            .I(\b2v_inst11.mult1_un152_sum_cry_3_s ));
    InMux I__6395 (
            .O(N__30169),
            .I(\b2v_inst11.mult1_un159_sum_cry_2 ));
    InMux I__6394 (
            .O(N__30166),
            .I(N__30163));
    LocalMux I__6393 (
            .O(N__30163),
            .I(N__30160));
    Span4Mux_s2_v I__6392 (
            .O(N__30160),
            .I(N__30157));
    Span4Mux_v I__6391 (
            .O(N__30157),
            .I(N__30154));
    Span4Mux_v I__6390 (
            .O(N__30154),
            .I(N__30151));
    Odrv4 I__6389 (
            .O(N__30151),
            .I(\b2v_inst11.mult1_un152_sum_cry_4_s ));
    InMux I__6388 (
            .O(N__30148),
            .I(\b2v_inst11.mult1_un159_sum_cry_3 ));
    InMux I__6387 (
            .O(N__30145),
            .I(N__30142));
    LocalMux I__6386 (
            .O(N__30142),
            .I(N__30139));
    Span4Mux_s2_v I__6385 (
            .O(N__30139),
            .I(N__30136));
    Span4Mux_v I__6384 (
            .O(N__30136),
            .I(N__30133));
    Span4Mux_v I__6383 (
            .O(N__30133),
            .I(N__30130));
    Odrv4 I__6382 (
            .O(N__30130),
            .I(\b2v_inst11.mult1_un152_sum_cry_5_s ));
    InMux I__6381 (
            .O(N__30127),
            .I(\b2v_inst11.mult1_un159_sum_cry_4 ));
    InMux I__6380 (
            .O(N__30124),
            .I(N__30121));
    LocalMux I__6379 (
            .O(N__30121),
            .I(N__30118));
    Span4Mux_s2_v I__6378 (
            .O(N__30118),
            .I(N__30115));
    Span4Mux_v I__6377 (
            .O(N__30115),
            .I(N__30112));
    Span4Mux_v I__6376 (
            .O(N__30112),
            .I(N__30109));
    Odrv4 I__6375 (
            .O(N__30109),
            .I(\b2v_inst11.mult1_un152_sum_cry_6_s ));
    InMux I__6374 (
            .O(N__30106),
            .I(\b2v_inst11.mult1_un159_sum_cry_5 ));
    InMux I__6373 (
            .O(N__30103),
            .I(N__30100));
    LocalMux I__6372 (
            .O(N__30100),
            .I(N__30097));
    Span12Mux_s10_v I__6371 (
            .O(N__30097),
            .I(N__30094));
    Odrv12 I__6370 (
            .O(N__30094),
            .I(\b2v_inst11.mult1_un159_sum_axb_7 ));
    InMux I__6369 (
            .O(N__30091),
            .I(\b2v_inst11.mult1_un159_sum_cry_6 ));
    InMux I__6368 (
            .O(N__30088),
            .I(N__30083));
    InMux I__6367 (
            .O(N__30087),
            .I(N__30080));
    InMux I__6366 (
            .O(N__30086),
            .I(N__30077));
    LocalMux I__6365 (
            .O(N__30083),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    LocalMux I__6364 (
            .O(N__30080),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    LocalMux I__6363 (
            .O(N__30077),
            .I(\b2v_inst11.mult1_un47_sum_s_6 ));
    CascadeMux I__6362 (
            .O(N__30070),
            .I(N__30067));
    InMux I__6361 (
            .O(N__30067),
            .I(N__30064));
    LocalMux I__6360 (
            .O(N__30064),
            .I(\b2v_inst11.mult1_un47_sum_l_fx_6 ));
    InMux I__6359 (
            .O(N__30061),
            .I(\b2v_inst11.mult1_un54_sum_cry_6 ));
    CascadeMux I__6358 (
            .O(N__30058),
            .I(N__30055));
    InMux I__6357 (
            .O(N__30055),
            .I(N__30051));
    CascadeMux I__6356 (
            .O(N__30054),
            .I(N__30048));
    LocalMux I__6355 (
            .O(N__30051),
            .I(N__30045));
    InMux I__6354 (
            .O(N__30048),
            .I(N__30042));
    Odrv4 I__6353 (
            .O(N__30045),
            .I(\b2v_inst11.mult1_un40_sum_i_5 ));
    LocalMux I__6352 (
            .O(N__30042),
            .I(\b2v_inst11.mult1_un40_sum_i_5 ));
    InMux I__6351 (
            .O(N__30037),
            .I(\b2v_inst11.mult1_un54_sum_cry_7 ));
    InMux I__6350 (
            .O(N__30034),
            .I(N__30031));
    LocalMux I__6349 (
            .O(N__30031),
            .I(\b2v_inst11.mult1_un47_sum_l_fx_3 ));
    CascadeMux I__6348 (
            .O(N__30028),
            .I(N__30025));
    InMux I__6347 (
            .O(N__30025),
            .I(N__30021));
    InMux I__6346 (
            .O(N__30024),
            .I(N__30018));
    LocalMux I__6345 (
            .O(N__30021),
            .I(N__30015));
    LocalMux I__6344 (
            .O(N__30018),
            .I(\b2v_inst11.mult1_un47_sum ));
    Odrv12 I__6343 (
            .O(N__30015),
            .I(\b2v_inst11.mult1_un47_sum ));
    CascadeMux I__6342 (
            .O(N__30010),
            .I(N__30007));
    InMux I__6341 (
            .O(N__30007),
            .I(N__30000));
    InMux I__6340 (
            .O(N__30006),
            .I(N__30000));
    InMux I__6339 (
            .O(N__30005),
            .I(N__29997));
    LocalMux I__6338 (
            .O(N__30000),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    LocalMux I__6337 (
            .O(N__29997),
            .I(\b2v_inst11.mult1_un47_sum_cry_3_s ));
    InMux I__6336 (
            .O(N__29992),
            .I(\b2v_inst11.mult1_un47_sum_cry_2 ));
    CascadeMux I__6335 (
            .O(N__29989),
            .I(N__29986));
    InMux I__6334 (
            .O(N__29986),
            .I(N__29983));
    LocalMux I__6333 (
            .O(N__29983),
            .I(N__29980));
    Odrv4 I__6332 (
            .O(N__29980),
            .I(\b2v_inst11.mult1_un47_sum_s_4_sf ));
    CascadeMux I__6331 (
            .O(N__29977),
            .I(N__29974));
    InMux I__6330 (
            .O(N__29974),
            .I(N__29971));
    LocalMux I__6329 (
            .O(N__29971),
            .I(\b2v_inst11.mult1_un47_sum_cry_4_s ));
    InMux I__6328 (
            .O(N__29968),
            .I(\b2v_inst11.mult1_un47_sum_cry_3 ));
    CascadeMux I__6327 (
            .O(N__29965),
            .I(N__29962));
    InMux I__6326 (
            .O(N__29962),
            .I(N__29959));
    LocalMux I__6325 (
            .O(N__29959),
            .I(N__29956));
    Odrv4 I__6324 (
            .O(N__29956),
            .I(\b2v_inst11.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__6323 (
            .O(N__29953),
            .I(N__29950));
    InMux I__6322 (
            .O(N__29950),
            .I(N__29947));
    LocalMux I__6321 (
            .O(N__29947),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_s ));
    InMux I__6320 (
            .O(N__29944),
            .I(\b2v_inst11.mult1_un47_sum_cry_4 ));
    InMux I__6319 (
            .O(N__29941),
            .I(\b2v_inst11.mult1_un47_sum_cry_5 ));
    InMux I__6318 (
            .O(N__29938),
            .I(N__29934));
    InMux I__6317 (
            .O(N__29937),
            .I(N__29931));
    LocalMux I__6316 (
            .O(N__29934),
            .I(N__29928));
    LocalMux I__6315 (
            .O(N__29931),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ));
    Odrv4 I__6314 (
            .O(N__29928),
            .I(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ));
    CascadeMux I__6313 (
            .O(N__29923),
            .I(N__29917));
    InMux I__6312 (
            .O(N__29922),
            .I(N__29914));
    InMux I__6311 (
            .O(N__29921),
            .I(N__29911));
    InMux I__6310 (
            .O(N__29920),
            .I(N__29906));
    InMux I__6309 (
            .O(N__29917),
            .I(N__29906));
    LocalMux I__6308 (
            .O(N__29914),
            .I(N__29901));
    LocalMux I__6307 (
            .O(N__29911),
            .I(N__29901));
    LocalMux I__6306 (
            .O(N__29906),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ));
    Odrv12 I__6305 (
            .O(N__29901),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ));
    CascadeMux I__6304 (
            .O(N__29896),
            .I(N__29893));
    InMux I__6303 (
            .O(N__29893),
            .I(N__29890));
    LocalMux I__6302 (
            .O(N__29890),
            .I(\b2v_inst11.un1_dutycycle_53_i_29 ));
    CascadeMux I__6301 (
            .O(N__29887),
            .I(N__29884));
    InMux I__6300 (
            .O(N__29884),
            .I(N__29880));
    CascadeMux I__6299 (
            .O(N__29883),
            .I(N__29871));
    LocalMux I__6298 (
            .O(N__29880),
            .I(N__29868));
    InMux I__6297 (
            .O(N__29879),
            .I(N__29863));
    InMux I__6296 (
            .O(N__29878),
            .I(N__29863));
    InMux I__6295 (
            .O(N__29877),
            .I(N__29856));
    InMux I__6294 (
            .O(N__29876),
            .I(N__29856));
    InMux I__6293 (
            .O(N__29875),
            .I(N__29856));
    InMux I__6292 (
            .O(N__29874),
            .I(N__29851));
    InMux I__6291 (
            .O(N__29871),
            .I(N__29851));
    Span4Mux_s3_h I__6290 (
            .O(N__29868),
            .I(N__29846));
    LocalMux I__6289 (
            .O(N__29863),
            .I(N__29846));
    LocalMux I__6288 (
            .O(N__29856),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    LocalMux I__6287 (
            .O(N__29851),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    Odrv4 I__6286 (
            .O(N__29846),
            .I(\b2v_inst11.curr_stateZ0Z_0 ));
    InMux I__6285 (
            .O(N__29839),
            .I(N__29833));
    InMux I__6284 (
            .O(N__29838),
            .I(N__29829));
    InMux I__6283 (
            .O(N__29837),
            .I(N__29824));
    InMux I__6282 (
            .O(N__29836),
            .I(N__29824));
    LocalMux I__6281 (
            .O(N__29833),
            .I(N__29821));
    InMux I__6280 (
            .O(N__29832),
            .I(N__29818));
    LocalMux I__6279 (
            .O(N__29829),
            .I(N__29813));
    LocalMux I__6278 (
            .O(N__29824),
            .I(N__29813));
    Odrv4 I__6277 (
            .O(N__29821),
            .I(\b2v_inst11.count_RNIZ0Z_13 ));
    LocalMux I__6276 (
            .O(N__29818),
            .I(\b2v_inst11.count_RNIZ0Z_13 ));
    Odrv4 I__6275 (
            .O(N__29813),
            .I(\b2v_inst11.count_RNIZ0Z_13 ));
    InMux I__6274 (
            .O(N__29806),
            .I(N__29803));
    LocalMux I__6273 (
            .O(N__29803),
            .I(N__29800));
    Span4Mux_s3_v I__6272 (
            .O(N__29800),
            .I(N__29797));
    Odrv4 I__6271 (
            .O(N__29797),
            .I(\b2v_inst11.curr_state_4_0 ));
    CascadeMux I__6270 (
            .O(N__29794),
            .I(N__29790));
    InMux I__6269 (
            .O(N__29793),
            .I(N__29787));
    InMux I__6268 (
            .O(N__29790),
            .I(N__29784));
    LocalMux I__6267 (
            .O(N__29787),
            .I(\b2v_inst11.CO2_THRU_CO ));
    LocalMux I__6266 (
            .O(N__29784),
            .I(\b2v_inst11.CO2_THRU_CO ));
    CascadeMux I__6265 (
            .O(N__29779),
            .I(N__29775));
    InMux I__6264 (
            .O(N__29778),
            .I(N__29771));
    InMux I__6263 (
            .O(N__29775),
            .I(N__29766));
    InMux I__6262 (
            .O(N__29774),
            .I(N__29766));
    LocalMux I__6261 (
            .O(N__29771),
            .I(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ));
    LocalMux I__6260 (
            .O(N__29766),
            .I(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ));
    CascadeMux I__6259 (
            .O(N__29761),
            .I(N__29758));
    InMux I__6258 (
            .O(N__29758),
            .I(N__29755));
    LocalMux I__6257 (
            .O(N__29755),
            .I(N__29752));
    Odrv4 I__6256 (
            .O(N__29752),
            .I(\b2v_inst11.mult1_un47_sum_i ));
    InMux I__6255 (
            .O(N__29749),
            .I(\b2v_inst11.mult1_un54_sum_cry_2 ));
    InMux I__6254 (
            .O(N__29746),
            .I(\b2v_inst11.mult1_un54_sum_cry_3 ));
    InMux I__6253 (
            .O(N__29743),
            .I(\b2v_inst11.mult1_un54_sum_cry_4 ));
    InMux I__6252 (
            .O(N__29740),
            .I(\b2v_inst11.mult1_un54_sum_cry_5 ));
    CascadeMux I__6251 (
            .O(N__29737),
            .I(N__29733));
    InMux I__6250 (
            .O(N__29736),
            .I(N__29727));
    InMux I__6249 (
            .O(N__29733),
            .I(N__29722));
    InMux I__6248 (
            .O(N__29732),
            .I(N__29719));
    InMux I__6247 (
            .O(N__29731),
            .I(N__29716));
    InMux I__6246 (
            .O(N__29730),
            .I(N__29713));
    LocalMux I__6245 (
            .O(N__29727),
            .I(N__29710));
    InMux I__6244 (
            .O(N__29726),
            .I(N__29707));
    CascadeMux I__6243 (
            .O(N__29725),
            .I(N__29702));
    LocalMux I__6242 (
            .O(N__29722),
            .I(N__29699));
    LocalMux I__6241 (
            .O(N__29719),
            .I(N__29696));
    LocalMux I__6240 (
            .O(N__29716),
            .I(N__29691));
    LocalMux I__6239 (
            .O(N__29713),
            .I(N__29691));
    Span4Mux_h I__6238 (
            .O(N__29710),
            .I(N__29688));
    LocalMux I__6237 (
            .O(N__29707),
            .I(N__29685));
    InMux I__6236 (
            .O(N__29706),
            .I(N__29680));
    InMux I__6235 (
            .O(N__29705),
            .I(N__29680));
    InMux I__6234 (
            .O(N__29702),
            .I(N__29677));
    Span4Mux_h I__6233 (
            .O(N__29699),
            .I(N__29670));
    Span4Mux_v I__6232 (
            .O(N__29696),
            .I(N__29670));
    Span4Mux_v I__6231 (
            .O(N__29691),
            .I(N__29670));
    Odrv4 I__6230 (
            .O(N__29688),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__6229 (
            .O(N__29685),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__6228 (
            .O(N__29680),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    LocalMux I__6227 (
            .O(N__29677),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    Odrv4 I__6226 (
            .O(N__29670),
            .I(\b2v_inst11.dutycycleZ0Z_12 ));
    CascadeMux I__6225 (
            .O(N__29659),
            .I(N__29656));
    InMux I__6224 (
            .O(N__29656),
            .I(N__29653));
    LocalMux I__6223 (
            .O(N__29653),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_13 ));
    InMux I__6222 (
            .O(N__29650),
            .I(\b2v_inst11.un1_dutycycle_53_cry_13 ));
    CascadeMux I__6221 (
            .O(N__29647),
            .I(N__29644));
    InMux I__6220 (
            .O(N__29644),
            .I(N__29641));
    LocalMux I__6219 (
            .O(N__29641),
            .I(N__29638));
    Span4Mux_h I__6218 (
            .O(N__29638),
            .I(N__29635));
    Span4Mux_v I__6217 (
            .O(N__29635),
            .I(N__29632));
    Odrv4 I__6216 (
            .O(N__29632),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_15 ));
    InMux I__6215 (
            .O(N__29629),
            .I(\b2v_inst11.un1_dutycycle_53_cry_14 ));
    InMux I__6214 (
            .O(N__29626),
            .I(N__29623));
    LocalMux I__6213 (
            .O(N__29623),
            .I(N__29620));
    Span4Mux_v I__6212 (
            .O(N__29620),
            .I(N__29617));
    Odrv4 I__6211 (
            .O(N__29617),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_14 ));
    InMux I__6210 (
            .O(N__29614),
            .I(N__29609));
    InMux I__6209 (
            .O(N__29613),
            .I(N__29604));
    InMux I__6208 (
            .O(N__29612),
            .I(N__29601));
    LocalMux I__6207 (
            .O(N__29609),
            .I(N__29598));
    InMux I__6206 (
            .O(N__29608),
            .I(N__29595));
    CascadeMux I__6205 (
            .O(N__29607),
            .I(N__29591));
    LocalMux I__6204 (
            .O(N__29604),
            .I(N__29586));
    LocalMux I__6203 (
            .O(N__29601),
            .I(N__29583));
    Span4Mux_h I__6202 (
            .O(N__29598),
            .I(N__29580));
    LocalMux I__6201 (
            .O(N__29595),
            .I(N__29577));
    InMux I__6200 (
            .O(N__29594),
            .I(N__29574));
    InMux I__6199 (
            .O(N__29591),
            .I(N__29571));
    InMux I__6198 (
            .O(N__29590),
            .I(N__29568));
    InMux I__6197 (
            .O(N__29589),
            .I(N__29565));
    Span4Mux_h I__6196 (
            .O(N__29586),
            .I(N__29560));
    Span4Mux_h I__6195 (
            .O(N__29583),
            .I(N__29560));
    Odrv4 I__6194 (
            .O(N__29580),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    Odrv12 I__6193 (
            .O(N__29577),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__6192 (
            .O(N__29574),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__6191 (
            .O(N__29571),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__6190 (
            .O(N__29568),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    LocalMux I__6189 (
            .O(N__29565),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    Odrv4 I__6188 (
            .O(N__29560),
            .I(\b2v_inst11.dutycycleZ0Z_11 ));
    InMux I__6187 (
            .O(N__29545),
            .I(bfn_9_11_0_));
    InMux I__6186 (
            .O(N__29542),
            .I(\b2v_inst11.CO2 ));
    CascadeMux I__6185 (
            .O(N__29539),
            .I(N__29527));
    InMux I__6184 (
            .O(N__29538),
            .I(N__29519));
    InMux I__6183 (
            .O(N__29537),
            .I(N__29519));
    CascadeMux I__6182 (
            .O(N__29536),
            .I(N__29513));
    CascadeMux I__6181 (
            .O(N__29535),
            .I(N__29510));
    InMux I__6180 (
            .O(N__29534),
            .I(N__29506));
    InMux I__6179 (
            .O(N__29533),
            .I(N__29503));
    CascadeMux I__6178 (
            .O(N__29532),
            .I(N__29500));
    InMux I__6177 (
            .O(N__29531),
            .I(N__29495));
    CascadeMux I__6176 (
            .O(N__29530),
            .I(N__29492));
    InMux I__6175 (
            .O(N__29527),
            .I(N__29483));
    InMux I__6174 (
            .O(N__29526),
            .I(N__29483));
    InMux I__6173 (
            .O(N__29525),
            .I(N__29483));
    InMux I__6172 (
            .O(N__29524),
            .I(N__29479));
    LocalMux I__6171 (
            .O(N__29519),
            .I(N__29476));
    InMux I__6170 (
            .O(N__29518),
            .I(N__29465));
    InMux I__6169 (
            .O(N__29517),
            .I(N__29465));
    InMux I__6168 (
            .O(N__29516),
            .I(N__29465));
    InMux I__6167 (
            .O(N__29513),
            .I(N__29465));
    InMux I__6166 (
            .O(N__29510),
            .I(N__29465));
    InMux I__6165 (
            .O(N__29509),
            .I(N__29462));
    LocalMux I__6164 (
            .O(N__29506),
            .I(N__29459));
    LocalMux I__6163 (
            .O(N__29503),
            .I(N__29456));
    InMux I__6162 (
            .O(N__29500),
            .I(N__29449));
    InMux I__6161 (
            .O(N__29499),
            .I(N__29449));
    InMux I__6160 (
            .O(N__29498),
            .I(N__29449));
    LocalMux I__6159 (
            .O(N__29495),
            .I(N__29446));
    InMux I__6158 (
            .O(N__29492),
            .I(N__29439));
    InMux I__6157 (
            .O(N__29491),
            .I(N__29439));
    InMux I__6156 (
            .O(N__29490),
            .I(N__29439));
    LocalMux I__6155 (
            .O(N__29483),
            .I(N__29436));
    InMux I__6154 (
            .O(N__29482),
            .I(N__29433));
    LocalMux I__6153 (
            .O(N__29479),
            .I(N__29426));
    Span4Mux_v I__6152 (
            .O(N__29476),
            .I(N__29426));
    LocalMux I__6151 (
            .O(N__29465),
            .I(N__29426));
    LocalMux I__6150 (
            .O(N__29462),
            .I(N__29417));
    Span4Mux_h I__6149 (
            .O(N__29459),
            .I(N__29417));
    Span4Mux_h I__6148 (
            .O(N__29456),
            .I(N__29417));
    LocalMux I__6147 (
            .O(N__29449),
            .I(N__29417));
    Span4Mux_h I__6146 (
            .O(N__29446),
            .I(N__29410));
    LocalMux I__6145 (
            .O(N__29439),
            .I(N__29410));
    Span4Mux_h I__6144 (
            .O(N__29436),
            .I(N__29410));
    LocalMux I__6143 (
            .O(N__29433),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__6142 (
            .O(N__29426),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__6141 (
            .O(N__29417),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    Odrv4 I__6140 (
            .O(N__29410),
            .I(\b2v_inst11.dutycycleZ0Z_7 ));
    CascadeMux I__6139 (
            .O(N__29401),
            .I(N__29394));
    CascadeMux I__6138 (
            .O(N__29400),
            .I(N__29385));
    InMux I__6137 (
            .O(N__29399),
            .I(N__29382));
    InMux I__6136 (
            .O(N__29398),
            .I(N__29379));
    CascadeMux I__6135 (
            .O(N__29397),
            .I(N__29376));
    InMux I__6134 (
            .O(N__29394),
            .I(N__29371));
    InMux I__6133 (
            .O(N__29393),
            .I(N__29371));
    InMux I__6132 (
            .O(N__29392),
            .I(N__29368));
    InMux I__6131 (
            .O(N__29391),
            .I(N__29365));
    InMux I__6130 (
            .O(N__29390),
            .I(N__29362));
    CascadeMux I__6129 (
            .O(N__29389),
            .I(N__29359));
    InMux I__6128 (
            .O(N__29388),
            .I(N__29356));
    InMux I__6127 (
            .O(N__29385),
            .I(N__29353));
    LocalMux I__6126 (
            .O(N__29382),
            .I(N__29348));
    LocalMux I__6125 (
            .O(N__29379),
            .I(N__29348));
    InMux I__6124 (
            .O(N__29376),
            .I(N__29345));
    LocalMux I__6123 (
            .O(N__29371),
            .I(N__29341));
    LocalMux I__6122 (
            .O(N__29368),
            .I(N__29334));
    LocalMux I__6121 (
            .O(N__29365),
            .I(N__29334));
    LocalMux I__6120 (
            .O(N__29362),
            .I(N__29334));
    InMux I__6119 (
            .O(N__29359),
            .I(N__29331));
    LocalMux I__6118 (
            .O(N__29356),
            .I(N__29326));
    LocalMux I__6117 (
            .O(N__29353),
            .I(N__29323));
    Span4Mux_h I__6116 (
            .O(N__29348),
            .I(N__29320));
    LocalMux I__6115 (
            .O(N__29345),
            .I(N__29317));
    InMux I__6114 (
            .O(N__29344),
            .I(N__29314));
    Span4Mux_s3_h I__6113 (
            .O(N__29341),
            .I(N__29307));
    Span4Mux_v I__6112 (
            .O(N__29334),
            .I(N__29307));
    LocalMux I__6111 (
            .O(N__29331),
            .I(N__29307));
    InMux I__6110 (
            .O(N__29330),
            .I(N__29304));
    InMux I__6109 (
            .O(N__29329),
            .I(N__29301));
    Span4Mux_h I__6108 (
            .O(N__29326),
            .I(N__29298));
    Span12Mux_s4_h I__6107 (
            .O(N__29323),
            .I(N__29295));
    Span4Mux_v I__6106 (
            .O(N__29320),
            .I(N__29292));
    Span4Mux_h I__6105 (
            .O(N__29317),
            .I(N__29285));
    LocalMux I__6104 (
            .O(N__29314),
            .I(N__29285));
    Span4Mux_h I__6103 (
            .O(N__29307),
            .I(N__29285));
    LocalMux I__6102 (
            .O(N__29304),
            .I(dutycycle_RNISSAOS1_0_5));
    LocalMux I__6101 (
            .O(N__29301),
            .I(dutycycle_RNISSAOS1_0_5));
    Odrv4 I__6100 (
            .O(N__29298),
            .I(dutycycle_RNISSAOS1_0_5));
    Odrv12 I__6099 (
            .O(N__29295),
            .I(dutycycle_RNISSAOS1_0_5));
    Odrv4 I__6098 (
            .O(N__29292),
            .I(dutycycle_RNISSAOS1_0_5));
    Odrv4 I__6097 (
            .O(N__29285),
            .I(dutycycle_RNISSAOS1_0_5));
    CascadeMux I__6096 (
            .O(N__29272),
            .I(N__29269));
    InMux I__6095 (
            .O(N__29269),
            .I(N__29266));
    LocalMux I__6094 (
            .O(N__29266),
            .I(N__29263));
    Odrv4 I__6093 (
            .O(N__29263),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_1 ));
    InMux I__6092 (
            .O(N__29260),
            .I(N__29257));
    LocalMux I__6091 (
            .O(N__29257),
            .I(N__29254));
    Odrv4 I__6090 (
            .O(N__29254),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_9 ));
    InMux I__6089 (
            .O(N__29251),
            .I(N__29247));
    InMux I__6088 (
            .O(N__29250),
            .I(N__29244));
    LocalMux I__6087 (
            .O(N__29247),
            .I(\b2v_inst11.mult1_un103_sum ));
    LocalMux I__6086 (
            .O(N__29244),
            .I(\b2v_inst11.mult1_un103_sum ));
    InMux I__6085 (
            .O(N__29239),
            .I(\b2v_inst11.un1_dutycycle_53_cry_5 ));
    InMux I__6084 (
            .O(N__29236),
            .I(N__29233));
    LocalMux I__6083 (
            .O(N__29233),
            .I(N__29230));
    Span4Mux_h I__6082 (
            .O(N__29230),
            .I(N__29227));
    Odrv4 I__6081 (
            .O(N__29227),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_9 ));
    CascadeMux I__6080 (
            .O(N__29224),
            .I(N__29220));
    InMux I__6079 (
            .O(N__29223),
            .I(N__29212));
    InMux I__6078 (
            .O(N__29220),
            .I(N__29209));
    InMux I__6077 (
            .O(N__29219),
            .I(N__29204));
    InMux I__6076 (
            .O(N__29218),
            .I(N__29204));
    CascadeMux I__6075 (
            .O(N__29217),
            .I(N__29201));
    InMux I__6074 (
            .O(N__29216),
            .I(N__29195));
    CascadeMux I__6073 (
            .O(N__29215),
            .I(N__29192));
    LocalMux I__6072 (
            .O(N__29212),
            .I(N__29186));
    LocalMux I__6071 (
            .O(N__29209),
            .I(N__29181));
    LocalMux I__6070 (
            .O(N__29204),
            .I(N__29181));
    InMux I__6069 (
            .O(N__29201),
            .I(N__29178));
    InMux I__6068 (
            .O(N__29200),
            .I(N__29173));
    InMux I__6067 (
            .O(N__29199),
            .I(N__29173));
    InMux I__6066 (
            .O(N__29198),
            .I(N__29170));
    LocalMux I__6065 (
            .O(N__29195),
            .I(N__29167));
    InMux I__6064 (
            .O(N__29192),
            .I(N__29164));
    InMux I__6063 (
            .O(N__29191),
            .I(N__29157));
    InMux I__6062 (
            .O(N__29190),
            .I(N__29157));
    InMux I__6061 (
            .O(N__29189),
            .I(N__29157));
    Span4Mux_v I__6060 (
            .O(N__29186),
            .I(N__29152));
    Span4Mux_h I__6059 (
            .O(N__29181),
            .I(N__29152));
    LocalMux I__6058 (
            .O(N__29178),
            .I(N__29143));
    LocalMux I__6057 (
            .O(N__29173),
            .I(N__29143));
    LocalMux I__6056 (
            .O(N__29170),
            .I(N__29143));
    Span4Mux_h I__6055 (
            .O(N__29167),
            .I(N__29143));
    LocalMux I__6054 (
            .O(N__29164),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    LocalMux I__6053 (
            .O(N__29157),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__6052 (
            .O(N__29152),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    Odrv4 I__6051 (
            .O(N__29143),
            .I(\b2v_inst11.dutycycleZ0Z_4 ));
    InMux I__6050 (
            .O(N__29134),
            .I(\b2v_inst11.un1_dutycycle_53_cry_6 ));
    InMux I__6049 (
            .O(N__29131),
            .I(N__29125));
    InMux I__6048 (
            .O(N__29130),
            .I(N__29120));
    InMux I__6047 (
            .O(N__29129),
            .I(N__29120));
    InMux I__6046 (
            .O(N__29128),
            .I(N__29117));
    LocalMux I__6045 (
            .O(N__29125),
            .I(N__29112));
    LocalMux I__6044 (
            .O(N__29120),
            .I(N__29109));
    LocalMux I__6043 (
            .O(N__29117),
            .I(N__29106));
    InMux I__6042 (
            .O(N__29116),
            .I(N__29103));
    InMux I__6041 (
            .O(N__29115),
            .I(N__29098));
    Span4Mux_h I__6040 (
            .O(N__29112),
            .I(N__29095));
    Span4Mux_v I__6039 (
            .O(N__29109),
            .I(N__29088));
    Span4Mux_h I__6038 (
            .O(N__29106),
            .I(N__29088));
    LocalMux I__6037 (
            .O(N__29103),
            .I(N__29088));
    InMux I__6036 (
            .O(N__29102),
            .I(N__29083));
    InMux I__6035 (
            .O(N__29101),
            .I(N__29083));
    LocalMux I__6034 (
            .O(N__29098),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__6033 (
            .O(N__29095),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    Odrv4 I__6032 (
            .O(N__29088),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    LocalMux I__6031 (
            .O(N__29083),
            .I(\b2v_inst11.dutycycleZ0Z_6 ));
    CascadeMux I__6030 (
            .O(N__29074),
            .I(N__29071));
    InMux I__6029 (
            .O(N__29071),
            .I(N__29068));
    LocalMux I__6028 (
            .O(N__29068),
            .I(N__29065));
    Span4Mux_h I__6027 (
            .O(N__29065),
            .I(N__29062));
    Odrv4 I__6026 (
            .O(N__29062),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_11 ));
    InMux I__6025 (
            .O(N__29059),
            .I(bfn_9_10_0_));
    InMux I__6024 (
            .O(N__29056),
            .I(N__29053));
    LocalMux I__6023 (
            .O(N__29053),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_12 ));
    InMux I__6022 (
            .O(N__29050),
            .I(N__29041));
    InMux I__6021 (
            .O(N__29049),
            .I(N__29041));
    CascadeMux I__6020 (
            .O(N__29048),
            .I(N__29038));
    InMux I__6019 (
            .O(N__29047),
            .I(N__29034));
    CascadeMux I__6018 (
            .O(N__29046),
            .I(N__29030));
    LocalMux I__6017 (
            .O(N__29041),
            .I(N__29024));
    InMux I__6016 (
            .O(N__29038),
            .I(N__29021));
    InMux I__6015 (
            .O(N__29037),
            .I(N__29018));
    LocalMux I__6014 (
            .O(N__29034),
            .I(N__29015));
    InMux I__6013 (
            .O(N__29033),
            .I(N__29012));
    InMux I__6012 (
            .O(N__29030),
            .I(N__29009));
    CascadeMux I__6011 (
            .O(N__29029),
            .I(N__29006));
    CascadeMux I__6010 (
            .O(N__29028),
            .I(N__29002));
    CascadeMux I__6009 (
            .O(N__29027),
            .I(N__28997));
    Span4Mux_v I__6008 (
            .O(N__29024),
            .I(N__28994));
    LocalMux I__6007 (
            .O(N__29021),
            .I(N__28989));
    LocalMux I__6006 (
            .O(N__29018),
            .I(N__28989));
    Span4Mux_h I__6005 (
            .O(N__29015),
            .I(N__28986));
    LocalMux I__6004 (
            .O(N__29012),
            .I(N__28983));
    LocalMux I__6003 (
            .O(N__29009),
            .I(N__28980));
    InMux I__6002 (
            .O(N__29006),
            .I(N__28977));
    InMux I__6001 (
            .O(N__29005),
            .I(N__28974));
    InMux I__6000 (
            .O(N__29002),
            .I(N__28965));
    InMux I__5999 (
            .O(N__29001),
            .I(N__28965));
    InMux I__5998 (
            .O(N__29000),
            .I(N__28965));
    InMux I__5997 (
            .O(N__28997),
            .I(N__28965));
    Span4Mux_h I__5996 (
            .O(N__28994),
            .I(N__28960));
    Span4Mux_h I__5995 (
            .O(N__28989),
            .I(N__28960));
    Odrv4 I__5994 (
            .O(N__28986),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__5993 (
            .O(N__28983),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv12 I__5992 (
            .O(N__28980),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__5991 (
            .O(N__28977),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__5990 (
            .O(N__28974),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    LocalMux I__5989 (
            .O(N__28965),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    Odrv4 I__5988 (
            .O(N__28960),
            .I(\b2v_inst11.dutycycleZ0Z_9 ));
    InMux I__5987 (
            .O(N__28945),
            .I(\b2v_inst11.un1_dutycycle_53_cry_8 ));
    CascadeMux I__5986 (
            .O(N__28942),
            .I(N__28939));
    InMux I__5985 (
            .O(N__28939),
            .I(N__28936));
    LocalMux I__5984 (
            .O(N__28936),
            .I(N__28933));
    Span4Mux_v I__5983 (
            .O(N__28933),
            .I(N__28930));
    Odrv4 I__5982 (
            .O(N__28930),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_13 ));
    InMux I__5981 (
            .O(N__28927),
            .I(\b2v_inst11.un1_dutycycle_53_cry_9 ));
    CascadeMux I__5980 (
            .O(N__28924),
            .I(N__28921));
    InMux I__5979 (
            .O(N__28921),
            .I(N__28918));
    LocalMux I__5978 (
            .O(N__28918),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_14 ));
    InMux I__5977 (
            .O(N__28915),
            .I(\b2v_inst11.un1_dutycycle_53_cry_10 ));
    CascadeMux I__5976 (
            .O(N__28912),
            .I(N__28909));
    InMux I__5975 (
            .O(N__28909),
            .I(N__28906));
    LocalMux I__5974 (
            .O(N__28906),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_11 ));
    InMux I__5973 (
            .O(N__28903),
            .I(\b2v_inst11.un1_dutycycle_53_cry_11 ));
    InMux I__5972 (
            .O(N__28900),
            .I(N__28892));
    InMux I__5971 (
            .O(N__28899),
            .I(N__28889));
    InMux I__5970 (
            .O(N__28898),
            .I(N__28886));
    InMux I__5969 (
            .O(N__28897),
            .I(N__28883));
    InMux I__5968 (
            .O(N__28896),
            .I(N__28878));
    InMux I__5967 (
            .O(N__28895),
            .I(N__28875));
    LocalMux I__5966 (
            .O(N__28892),
            .I(N__28872));
    LocalMux I__5965 (
            .O(N__28889),
            .I(N__28865));
    LocalMux I__5964 (
            .O(N__28886),
            .I(N__28865));
    LocalMux I__5963 (
            .O(N__28883),
            .I(N__28865));
    InMux I__5962 (
            .O(N__28882),
            .I(N__28860));
    InMux I__5961 (
            .O(N__28881),
            .I(N__28860));
    LocalMux I__5960 (
            .O(N__28878),
            .I(N__28855));
    LocalMux I__5959 (
            .O(N__28875),
            .I(N__28855));
    Odrv12 I__5958 (
            .O(N__28872),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__5957 (
            .O(N__28865),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    LocalMux I__5956 (
            .O(N__28860),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    Odrv4 I__5955 (
            .O(N__28855),
            .I(\b2v_inst11.dutycycleZ0Z_8 ));
    CascadeMux I__5954 (
            .O(N__28846),
            .I(N__28843));
    InMux I__5953 (
            .O(N__28843),
            .I(N__28840));
    LocalMux I__5952 (
            .O(N__28840),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ));
    InMux I__5951 (
            .O(N__28837),
            .I(\b2v_inst11.un1_dutycycle_53_cry_12 ));
    InMux I__5950 (
            .O(N__28834),
            .I(\b2v_inst11.mult1_un103_sum_cry_7 ));
    CascadeMux I__5949 (
            .O(N__28831),
            .I(N__28826));
    InMux I__5948 (
            .O(N__28830),
            .I(N__28822));
    InMux I__5947 (
            .O(N__28829),
            .I(N__28817));
    InMux I__5946 (
            .O(N__28826),
            .I(N__28817));
    InMux I__5945 (
            .O(N__28825),
            .I(N__28814));
    LocalMux I__5944 (
            .O(N__28822),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    LocalMux I__5943 (
            .O(N__28817),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    LocalMux I__5942 (
            .O(N__28814),
            .I(\b2v_inst11.mult1_un103_sum_s_8 ));
    CascadeMux I__5941 (
            .O(N__28807),
            .I(\b2v_inst11.mult1_un103_sum_s_8_cascade_ ));
    CascadeMux I__5940 (
            .O(N__28804),
            .I(N__28800));
    CascadeMux I__5939 (
            .O(N__28803),
            .I(N__28796));
    InMux I__5938 (
            .O(N__28800),
            .I(N__28789));
    InMux I__5937 (
            .O(N__28799),
            .I(N__28789));
    InMux I__5936 (
            .O(N__28796),
            .I(N__28789));
    LocalMux I__5935 (
            .O(N__28789),
            .I(\b2v_inst11.mult1_un103_sum_i_0_8 ));
    InMux I__5934 (
            .O(N__28786),
            .I(N__28781));
    InMux I__5933 (
            .O(N__28785),
            .I(N__28776));
    InMux I__5932 (
            .O(N__28784),
            .I(N__28776));
    LocalMux I__5931 (
            .O(N__28781),
            .I(N__28769));
    LocalMux I__5930 (
            .O(N__28776),
            .I(N__28766));
    InMux I__5929 (
            .O(N__28775),
            .I(N__28759));
    InMux I__5928 (
            .O(N__28774),
            .I(N__28759));
    InMux I__5927 (
            .O(N__28773),
            .I(N__28759));
    InMux I__5926 (
            .O(N__28772),
            .I(N__28751));
    Span4Mux_v I__5925 (
            .O(N__28769),
            .I(N__28744));
    Span4Mux_v I__5924 (
            .O(N__28766),
            .I(N__28744));
    LocalMux I__5923 (
            .O(N__28759),
            .I(N__28744));
    CascadeMux I__5922 (
            .O(N__28758),
            .I(N__28741));
    CascadeMux I__5921 (
            .O(N__28757),
            .I(N__28738));
    InMux I__5920 (
            .O(N__28756),
            .I(N__28735));
    InMux I__5919 (
            .O(N__28755),
            .I(N__28730));
    InMux I__5918 (
            .O(N__28754),
            .I(N__28730));
    LocalMux I__5917 (
            .O(N__28751),
            .I(N__28725));
    Span4Mux_h I__5916 (
            .O(N__28744),
            .I(N__28725));
    InMux I__5915 (
            .O(N__28741),
            .I(N__28722));
    InMux I__5914 (
            .O(N__28738),
            .I(N__28719));
    LocalMux I__5913 (
            .O(N__28735),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__5912 (
            .O(N__28730),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    Odrv4 I__5911 (
            .O(N__28725),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__5910 (
            .O(N__28722),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    LocalMux I__5909 (
            .O(N__28719),
            .I(\b2v_inst11.dutycycleZ0Z_3 ));
    InMux I__5908 (
            .O(N__28708),
            .I(N__28704));
    InMux I__5907 (
            .O(N__28707),
            .I(N__28701));
    LocalMux I__5906 (
            .O(N__28704),
            .I(N__28696));
    LocalMux I__5905 (
            .O(N__28701),
            .I(N__28696));
    Odrv4 I__5904 (
            .O(N__28696),
            .I(\b2v_inst11.un1_dutycycle_53_axb_0 ));
    InMux I__5903 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__5902 (
            .O(N__28690),
            .I(N__28687));
    Span4Mux_h I__5901 (
            .O(N__28687),
            .I(N__28684));
    Odrv4 I__5900 (
            .O(N__28684),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_1 ));
    InMux I__5899 (
            .O(N__28681),
            .I(N__28678));
    LocalMux I__5898 (
            .O(N__28678),
            .I(N__28674));
    InMux I__5897 (
            .O(N__28677),
            .I(N__28671));
    Span4Mux_h I__5896 (
            .O(N__28674),
            .I(N__28666));
    LocalMux I__5895 (
            .O(N__28671),
            .I(N__28666));
    Span4Mux_v I__5894 (
            .O(N__28666),
            .I(N__28663));
    Odrv4 I__5893 (
            .O(N__28663),
            .I(\b2v_inst11.mult1_un138_sum ));
    InMux I__5892 (
            .O(N__28660),
            .I(\b2v_inst11.un1_dutycycle_53_cry_0 ));
    InMux I__5891 (
            .O(N__28657),
            .I(N__28653));
    InMux I__5890 (
            .O(N__28656),
            .I(N__28650));
    LocalMux I__5889 (
            .O(N__28653),
            .I(N__28647));
    LocalMux I__5888 (
            .O(N__28650),
            .I(N__28642));
    Span4Mux_h I__5887 (
            .O(N__28647),
            .I(N__28642));
    Odrv4 I__5886 (
            .O(N__28642),
            .I(\b2v_inst11.mult1_un131_sum ));
    InMux I__5885 (
            .O(N__28639),
            .I(\b2v_inst11.un1_dutycycle_53_cry_1 ));
    InMux I__5884 (
            .O(N__28636),
            .I(N__28633));
    LocalMux I__5883 (
            .O(N__28633),
            .I(N__28630));
    Odrv4 I__5882 (
            .O(N__28630),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_2 ));
    InMux I__5881 (
            .O(N__28627),
            .I(N__28623));
    InMux I__5880 (
            .O(N__28626),
            .I(N__28620));
    LocalMux I__5879 (
            .O(N__28623),
            .I(N__28615));
    LocalMux I__5878 (
            .O(N__28620),
            .I(N__28615));
    Span4Mux_h I__5877 (
            .O(N__28615),
            .I(N__28612));
    Odrv4 I__5876 (
            .O(N__28612),
            .I(\b2v_inst11.mult1_un124_sum ));
    InMux I__5875 (
            .O(N__28609),
            .I(\b2v_inst11.un1_dutycycle_53_cry_2 ));
    CascadeMux I__5874 (
            .O(N__28606),
            .I(N__28602));
    InMux I__5873 (
            .O(N__28605),
            .I(N__28599));
    InMux I__5872 (
            .O(N__28602),
            .I(N__28596));
    LocalMux I__5871 (
            .O(N__28599),
            .I(N__28593));
    LocalMux I__5870 (
            .O(N__28596),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_3 ));
    Odrv4 I__5869 (
            .O(N__28593),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_3 ));
    CascadeMux I__5868 (
            .O(N__28588),
            .I(N__28585));
    InMux I__5867 (
            .O(N__28585),
            .I(N__28582));
    LocalMux I__5866 (
            .O(N__28582),
            .I(N__28579));
    Odrv4 I__5865 (
            .O(N__28579),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_3 ));
    InMux I__5864 (
            .O(N__28576),
            .I(N__28572));
    InMux I__5863 (
            .O(N__28575),
            .I(N__28569));
    LocalMux I__5862 (
            .O(N__28572),
            .I(N__28564));
    LocalMux I__5861 (
            .O(N__28569),
            .I(N__28564));
    Odrv4 I__5860 (
            .O(N__28564),
            .I(\b2v_inst11.mult1_un117_sum ));
    InMux I__5859 (
            .O(N__28561),
            .I(\b2v_inst11.un1_dutycycle_53_cry_3 ));
    CascadeMux I__5858 (
            .O(N__28558),
            .I(N__28555));
    InMux I__5857 (
            .O(N__28555),
            .I(N__28552));
    LocalMux I__5856 (
            .O(N__28552),
            .I(N__28549));
    Span4Mux_s3_h I__5855 (
            .O(N__28549),
            .I(N__28546));
    Odrv4 I__5854 (
            .O(N__28546),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_8 ));
    InMux I__5853 (
            .O(N__28543),
            .I(N__28539));
    InMux I__5852 (
            .O(N__28542),
            .I(N__28536));
    LocalMux I__5851 (
            .O(N__28539),
            .I(N__28533));
    LocalMux I__5850 (
            .O(N__28536),
            .I(\b2v_inst11.mult1_un110_sum ));
    Odrv4 I__5849 (
            .O(N__28533),
            .I(\b2v_inst11.mult1_un110_sum ));
    InMux I__5848 (
            .O(N__28528),
            .I(\b2v_inst11.un1_dutycycle_53_cry_4 ));
    CascadeMux I__5847 (
            .O(N__28525),
            .I(N__28522));
    InMux I__5846 (
            .O(N__28522),
            .I(N__28519));
    LocalMux I__5845 (
            .O(N__28519),
            .I(\b2v_inst11.mult1_un117_sum_axb_8 ));
    InMux I__5844 (
            .O(N__28516),
            .I(\b2v_inst11.mult1_un110_sum_cry_6 ));
    InMux I__5843 (
            .O(N__28513),
            .I(\b2v_inst11.mult1_un110_sum_cry_7 ));
    CascadeMux I__5842 (
            .O(N__28510),
            .I(\b2v_inst11.mult1_un110_sum_s_8_cascade_ ));
    CascadeMux I__5841 (
            .O(N__28507),
            .I(N__28503));
    CascadeMux I__5840 (
            .O(N__28506),
            .I(N__28499));
    InMux I__5839 (
            .O(N__28503),
            .I(N__28492));
    InMux I__5838 (
            .O(N__28502),
            .I(N__28492));
    InMux I__5837 (
            .O(N__28499),
            .I(N__28492));
    LocalMux I__5836 (
            .O(N__28492),
            .I(\b2v_inst11.mult1_un110_sum_i_0_8 ));
    CascadeMux I__5835 (
            .O(N__28489),
            .I(N__28486));
    InMux I__5834 (
            .O(N__28486),
            .I(N__28483));
    LocalMux I__5833 (
            .O(N__28483),
            .I(\b2v_inst11.mult1_un103_sum_cry_3_s ));
    InMux I__5832 (
            .O(N__28480),
            .I(\b2v_inst11.mult1_un103_sum_cry_2 ));
    InMux I__5831 (
            .O(N__28477),
            .I(N__28474));
    LocalMux I__5830 (
            .O(N__28474),
            .I(\b2v_inst11.mult1_un103_sum_cry_4_s ));
    InMux I__5829 (
            .O(N__28471),
            .I(\b2v_inst11.mult1_un103_sum_cry_3 ));
    CascadeMux I__5828 (
            .O(N__28468),
            .I(N__28465));
    InMux I__5827 (
            .O(N__28465),
            .I(N__28462));
    LocalMux I__5826 (
            .O(N__28462),
            .I(\b2v_inst11.mult1_un103_sum_cry_5_s ));
    InMux I__5825 (
            .O(N__28459),
            .I(\b2v_inst11.mult1_un103_sum_cry_4 ));
    InMux I__5824 (
            .O(N__28456),
            .I(N__28453));
    LocalMux I__5823 (
            .O(N__28453),
            .I(\b2v_inst11.mult1_un103_sum_cry_6_s ));
    InMux I__5822 (
            .O(N__28450),
            .I(\b2v_inst11.mult1_un103_sum_cry_5 ));
    CascadeMux I__5821 (
            .O(N__28447),
            .I(N__28443));
    CascadeMux I__5820 (
            .O(N__28446),
            .I(N__28439));
    InMux I__5819 (
            .O(N__28443),
            .I(N__28432));
    InMux I__5818 (
            .O(N__28442),
            .I(N__28432));
    InMux I__5817 (
            .O(N__28439),
            .I(N__28432));
    LocalMux I__5816 (
            .O(N__28432),
            .I(\b2v_inst11.mult1_un96_sum_i_0_8 ));
    CascadeMux I__5815 (
            .O(N__28429),
            .I(N__28426));
    InMux I__5814 (
            .O(N__28426),
            .I(N__28423));
    LocalMux I__5813 (
            .O(N__28423),
            .I(\b2v_inst11.mult1_un110_sum_axb_8 ));
    InMux I__5812 (
            .O(N__28420),
            .I(\b2v_inst11.mult1_un103_sum_cry_6 ));
    CascadeMux I__5811 (
            .O(N__28417),
            .I(N__28414));
    InMux I__5810 (
            .O(N__28414),
            .I(N__28411));
    LocalMux I__5809 (
            .O(N__28411),
            .I(\b2v_inst11.mult1_un138_sum_cry_6_s ));
    InMux I__5808 (
            .O(N__28408),
            .I(N__28405));
    LocalMux I__5807 (
            .O(N__28405),
            .I(N__28402));
    Odrv4 I__5806 (
            .O(N__28402),
            .I(\b2v_inst11.mult1_un152_sum_axb_8 ));
    InMux I__5805 (
            .O(N__28399),
            .I(\b2v_inst11.mult1_un145_sum_cry_6 ));
    InMux I__5804 (
            .O(N__28396),
            .I(N__28393));
    LocalMux I__5803 (
            .O(N__28393),
            .I(\b2v_inst11.mult1_un145_sum_axb_8 ));
    InMux I__5802 (
            .O(N__28390),
            .I(\b2v_inst11.mult1_un145_sum_cry_7 ));
    CascadeMux I__5801 (
            .O(N__28387),
            .I(N__28382));
    CascadeMux I__5800 (
            .O(N__28386),
            .I(N__28379));
    InMux I__5799 (
            .O(N__28385),
            .I(N__28374));
    InMux I__5798 (
            .O(N__28382),
            .I(N__28374));
    InMux I__5797 (
            .O(N__28379),
            .I(N__28371));
    LocalMux I__5796 (
            .O(N__28374),
            .I(\b2v_inst11.mult1_un138_sum_i_0_8 ));
    LocalMux I__5795 (
            .O(N__28371),
            .I(\b2v_inst11.mult1_un138_sum_i_0_8 ));
    InMux I__5794 (
            .O(N__28366),
            .I(N__28363));
    LocalMux I__5793 (
            .O(N__28363),
            .I(\b2v_inst11.mult1_un103_sum_i ));
    CascadeMux I__5792 (
            .O(N__28360),
            .I(N__28357));
    InMux I__5791 (
            .O(N__28357),
            .I(N__28354));
    LocalMux I__5790 (
            .O(N__28354),
            .I(\b2v_inst11.mult1_un110_sum_cry_3_s ));
    InMux I__5789 (
            .O(N__28351),
            .I(\b2v_inst11.mult1_un110_sum_cry_2 ));
    InMux I__5788 (
            .O(N__28348),
            .I(N__28345));
    LocalMux I__5787 (
            .O(N__28345),
            .I(\b2v_inst11.mult1_un110_sum_cry_4_s ));
    InMux I__5786 (
            .O(N__28342),
            .I(\b2v_inst11.mult1_un110_sum_cry_3 ));
    CascadeMux I__5785 (
            .O(N__28339),
            .I(N__28336));
    InMux I__5784 (
            .O(N__28336),
            .I(N__28333));
    LocalMux I__5783 (
            .O(N__28333),
            .I(\b2v_inst11.mult1_un110_sum_cry_5_s ));
    InMux I__5782 (
            .O(N__28330),
            .I(\b2v_inst11.mult1_un110_sum_cry_4 ));
    InMux I__5781 (
            .O(N__28327),
            .I(N__28324));
    LocalMux I__5780 (
            .O(N__28324),
            .I(\b2v_inst11.mult1_un110_sum_cry_6_s ));
    InMux I__5779 (
            .O(N__28321),
            .I(\b2v_inst11.mult1_un110_sum_cry_5 ));
    CascadeMux I__5778 (
            .O(N__28318),
            .I(\b2v_inst5.un2_count_1_axb_13_cascade_ ));
    InMux I__5777 (
            .O(N__28315),
            .I(N__28312));
    LocalMux I__5776 (
            .O(N__28312),
            .I(\b2v_inst5.count_rst_1 ));
    CascadeMux I__5775 (
            .O(N__28309),
            .I(N__28306));
    InMux I__5774 (
            .O(N__28306),
            .I(N__28302));
    InMux I__5773 (
            .O(N__28305),
            .I(N__28299));
    LocalMux I__5772 (
            .O(N__28302),
            .I(\b2v_inst5.count_1_13 ));
    LocalMux I__5771 (
            .O(N__28299),
            .I(\b2v_inst5.count_1_13 ));
    InMux I__5770 (
            .O(N__28294),
            .I(N__28291));
    LocalMux I__5769 (
            .O(N__28291),
            .I(N__28288));
    Span4Mux_v I__5768 (
            .O(N__28288),
            .I(N__28285));
    Odrv4 I__5767 (
            .O(N__28285),
            .I(\b2v_inst5.un12_clk_100khz_5 ));
    InMux I__5766 (
            .O(N__28282),
            .I(N__28279));
    LocalMux I__5765 (
            .O(N__28279),
            .I(N__28276));
    Span4Mux_h I__5764 (
            .O(N__28276),
            .I(N__28273));
    Odrv4 I__5763 (
            .O(N__28273),
            .I(\b2v_inst5.count_rst_6 ));
    InMux I__5762 (
            .O(N__28270),
            .I(N__28267));
    LocalMux I__5761 (
            .O(N__28267),
            .I(N__28264));
    Odrv4 I__5760 (
            .O(N__28264),
            .I(\b2v_inst5.un12_clk_100khz_8 ));
    InMux I__5759 (
            .O(N__28261),
            .I(N__28258));
    LocalMux I__5758 (
            .O(N__28258),
            .I(N__28255));
    Span4Mux_v I__5757 (
            .O(N__28255),
            .I(N__28252));
    Odrv4 I__5756 (
            .O(N__28252),
            .I(\b2v_inst11.mult1_un138_sum_i ));
    InMux I__5755 (
            .O(N__28249),
            .I(N__28246));
    LocalMux I__5754 (
            .O(N__28246),
            .I(N__28243));
    Odrv12 I__5753 (
            .O(N__28243),
            .I(\b2v_inst11.mult1_un145_sum_cry_3_s ));
    InMux I__5752 (
            .O(N__28240),
            .I(\b2v_inst11.mult1_un145_sum_cry_2 ));
    InMux I__5751 (
            .O(N__28237),
            .I(N__28234));
    LocalMux I__5750 (
            .O(N__28234),
            .I(\b2v_inst11.mult1_un138_sum_cry_3_s ));
    InMux I__5749 (
            .O(N__28231),
            .I(N__28228));
    LocalMux I__5748 (
            .O(N__28228),
            .I(N__28225));
    Odrv12 I__5747 (
            .O(N__28225),
            .I(\b2v_inst11.mult1_un145_sum_cry_4_s ));
    InMux I__5746 (
            .O(N__28222),
            .I(\b2v_inst11.mult1_un145_sum_cry_3 ));
    CascadeMux I__5745 (
            .O(N__28219),
            .I(N__28216));
    InMux I__5744 (
            .O(N__28216),
            .I(N__28213));
    LocalMux I__5743 (
            .O(N__28213),
            .I(\b2v_inst11.mult1_un138_sum_cry_4_s ));
    InMux I__5742 (
            .O(N__28210),
            .I(N__28207));
    LocalMux I__5741 (
            .O(N__28207),
            .I(N__28204));
    Odrv4 I__5740 (
            .O(N__28204),
            .I(\b2v_inst11.mult1_un145_sum_cry_5_s ));
    InMux I__5739 (
            .O(N__28201),
            .I(\b2v_inst11.mult1_un145_sum_cry_4 ));
    InMux I__5738 (
            .O(N__28198),
            .I(N__28195));
    LocalMux I__5737 (
            .O(N__28195),
            .I(\b2v_inst11.mult1_un138_sum_cry_5_s ));
    InMux I__5736 (
            .O(N__28192),
            .I(N__28189));
    LocalMux I__5735 (
            .O(N__28189),
            .I(N__28186));
    Odrv4 I__5734 (
            .O(N__28186),
            .I(\b2v_inst11.mult1_un145_sum_cry_6_s ));
    InMux I__5733 (
            .O(N__28183),
            .I(\b2v_inst11.mult1_un145_sum_cry_5 ));
    CascadeMux I__5732 (
            .O(N__28180),
            .I(\b2v_inst5.count_RNIZ0Z_1_cascade_ ));
    InMux I__5731 (
            .O(N__28177),
            .I(N__28174));
    LocalMux I__5730 (
            .O(N__28174),
            .I(\b2v_inst5.count_1_3 ));
    InMux I__5729 (
            .O(N__28171),
            .I(N__28168));
    LocalMux I__5728 (
            .O(N__28168),
            .I(\b2v_inst5.count_RNIZ0Z_1 ));
    InMux I__5727 (
            .O(N__28165),
            .I(N__28162));
    LocalMux I__5726 (
            .O(N__28162),
            .I(\b2v_inst5.count_1_1 ));
    CascadeMux I__5725 (
            .O(N__28159),
            .I(\b2v_inst5.count_rst_14_cascade_ ));
    CascadeMux I__5724 (
            .O(N__28156),
            .I(\b2v_inst5.count_rst_1_cascade_ ));
    CascadeMux I__5723 (
            .O(N__28153),
            .I(\b2v_inst36.count_rst_4_cascade_ ));
    InMux I__5722 (
            .O(N__28150),
            .I(N__28146));
    CascadeMux I__5721 (
            .O(N__28149),
            .I(N__28143));
    LocalMux I__5720 (
            .O(N__28146),
            .I(N__28139));
    InMux I__5719 (
            .O(N__28143),
            .I(N__28136));
    InMux I__5718 (
            .O(N__28142),
            .I(N__28133));
    Odrv4 I__5717 (
            .O(N__28139),
            .I(\b2v_inst36.countZ0Z_10 ));
    LocalMux I__5716 (
            .O(N__28136),
            .I(\b2v_inst36.countZ0Z_10 ));
    LocalMux I__5715 (
            .O(N__28133),
            .I(\b2v_inst36.countZ0Z_10 ));
    InMux I__5714 (
            .O(N__28126),
            .I(N__28120));
    InMux I__5713 (
            .O(N__28125),
            .I(N__28120));
    LocalMux I__5712 (
            .O(N__28120),
            .I(\b2v_inst36.un2_count_1_cry_9_THRU_CO ));
    CascadeMux I__5711 (
            .O(N__28117),
            .I(\b2v_inst36.countZ0Z_10_cascade_ ));
    InMux I__5710 (
            .O(N__28114),
            .I(N__28111));
    LocalMux I__5709 (
            .O(N__28111),
            .I(\b2v_inst36.count_2_10 ));
    InMux I__5708 (
            .O(N__28108),
            .I(N__28104));
    InMux I__5707 (
            .O(N__28107),
            .I(N__28101));
    LocalMux I__5706 (
            .O(N__28104),
            .I(\b2v_inst36.countZ0Z_13 ));
    LocalMux I__5705 (
            .O(N__28101),
            .I(\b2v_inst36.countZ0Z_13 ));
    InMux I__5704 (
            .O(N__28096),
            .I(N__28090));
    InMux I__5703 (
            .O(N__28095),
            .I(N__28090));
    LocalMux I__5702 (
            .O(N__28090),
            .I(\b2v_inst36.count_rst_1 ));
    InMux I__5701 (
            .O(N__28087),
            .I(N__28084));
    LocalMux I__5700 (
            .O(N__28084),
            .I(\b2v_inst36.count_2_13 ));
    InMux I__5699 (
            .O(N__28081),
            .I(N__28078));
    LocalMux I__5698 (
            .O(N__28078),
            .I(N__28075));
    Odrv12 I__5697 (
            .O(N__28075),
            .I(\b2v_inst36.count_2_15 ));
    InMux I__5696 (
            .O(N__28072),
            .I(N__28068));
    InMux I__5695 (
            .O(N__28071),
            .I(N__28065));
    LocalMux I__5694 (
            .O(N__28068),
            .I(\b2v_inst36.count_rst ));
    LocalMux I__5693 (
            .O(N__28065),
            .I(\b2v_inst36.count_rst ));
    InMux I__5692 (
            .O(N__28060),
            .I(N__28056));
    InMux I__5691 (
            .O(N__28059),
            .I(N__28053));
    LocalMux I__5690 (
            .O(N__28056),
            .I(\b2v_inst36.countZ0Z_15 ));
    LocalMux I__5689 (
            .O(N__28053),
            .I(\b2v_inst36.countZ0Z_15 ));
    InMux I__5688 (
            .O(N__28048),
            .I(N__28045));
    LocalMux I__5687 (
            .O(N__28045),
            .I(N__28042));
    Span4Mux_v I__5686 (
            .O(N__28042),
            .I(N__28039));
    Odrv4 I__5685 (
            .O(N__28039),
            .I(\b2v_inst5.un12_clk_100khz_4 ));
    InMux I__5684 (
            .O(N__28036),
            .I(N__28030));
    InMux I__5683 (
            .O(N__28035),
            .I(N__28030));
    LocalMux I__5682 (
            .O(N__28030),
            .I(\b2v_inst5.count_1_2 ));
    InMux I__5681 (
            .O(N__28027),
            .I(N__28022));
    InMux I__5680 (
            .O(N__28026),
            .I(N__28019));
    InMux I__5679 (
            .O(N__28025),
            .I(N__28016));
    LocalMux I__5678 (
            .O(N__28022),
            .I(\b2v_inst36.countZ0Z_11 ));
    LocalMux I__5677 (
            .O(N__28019),
            .I(\b2v_inst36.countZ0Z_11 ));
    LocalMux I__5676 (
            .O(N__28016),
            .I(\b2v_inst36.countZ0Z_11 ));
    InMux I__5675 (
            .O(N__28009),
            .I(N__28003));
    InMux I__5674 (
            .O(N__28008),
            .I(N__28003));
    LocalMux I__5673 (
            .O(N__28003),
            .I(\b2v_inst36.un2_count_1_cry_10_THRU_CO ));
    InMux I__5672 (
            .O(N__28000),
            .I(\b2v_inst36.un2_count_1_cry_10 ));
    InMux I__5671 (
            .O(N__27997),
            .I(N__27993));
    CascadeMux I__5670 (
            .O(N__27996),
            .I(N__27990));
    LocalMux I__5669 (
            .O(N__27993),
            .I(N__27987));
    InMux I__5668 (
            .O(N__27990),
            .I(N__27984));
    Span4Mux_h I__5667 (
            .O(N__27987),
            .I(N__27981));
    LocalMux I__5666 (
            .O(N__27984),
            .I(\b2v_inst36.countZ0Z_12 ));
    Odrv4 I__5665 (
            .O(N__27981),
            .I(\b2v_inst36.countZ0Z_12 ));
    InMux I__5664 (
            .O(N__27976),
            .I(N__27972));
    InMux I__5663 (
            .O(N__27975),
            .I(N__27969));
    LocalMux I__5662 (
            .O(N__27972),
            .I(N__27964));
    LocalMux I__5661 (
            .O(N__27969),
            .I(N__27964));
    Span4Mux_s1_v I__5660 (
            .O(N__27964),
            .I(N__27961));
    Odrv4 I__5659 (
            .O(N__27961),
            .I(\b2v_inst36.count_rst_2 ));
    InMux I__5658 (
            .O(N__27958),
            .I(\b2v_inst36.un2_count_1_cry_11 ));
    InMux I__5657 (
            .O(N__27955),
            .I(\b2v_inst36.un2_count_1_cry_12 ));
    CascadeMux I__5656 (
            .O(N__27952),
            .I(N__27949));
    InMux I__5655 (
            .O(N__27949),
            .I(N__27945));
    InMux I__5654 (
            .O(N__27948),
            .I(N__27942));
    LocalMux I__5653 (
            .O(N__27945),
            .I(N__27937));
    LocalMux I__5652 (
            .O(N__27942),
            .I(N__27937));
    Odrv4 I__5651 (
            .O(N__27937),
            .I(\b2v_inst36.countZ0Z_14 ));
    InMux I__5650 (
            .O(N__27934),
            .I(N__27930));
    InMux I__5649 (
            .O(N__27933),
            .I(N__27927));
    LocalMux I__5648 (
            .O(N__27930),
            .I(N__27924));
    LocalMux I__5647 (
            .O(N__27927),
            .I(N__27921));
    Odrv4 I__5646 (
            .O(N__27924),
            .I(\b2v_inst36.count_rst_0 ));
    Odrv4 I__5645 (
            .O(N__27921),
            .I(\b2v_inst36.count_rst_0 ));
    InMux I__5644 (
            .O(N__27916),
            .I(\b2v_inst36.un2_count_1_cry_13 ));
    InMux I__5643 (
            .O(N__27913),
            .I(\b2v_inst36.un2_count_1_cry_14 ));
    InMux I__5642 (
            .O(N__27910),
            .I(N__27907));
    LocalMux I__5641 (
            .O(N__27907),
            .I(\b2v_inst36.count_rst_6 ));
    InMux I__5640 (
            .O(N__27904),
            .I(N__27899));
    InMux I__5639 (
            .O(N__27903),
            .I(N__27896));
    InMux I__5638 (
            .O(N__27902),
            .I(N__27893));
    LocalMux I__5637 (
            .O(N__27899),
            .I(N__27890));
    LocalMux I__5636 (
            .O(N__27896),
            .I(N__27887));
    LocalMux I__5635 (
            .O(N__27893),
            .I(N__27884));
    Odrv4 I__5634 (
            .O(N__27890),
            .I(\b2v_inst36.countZ0Z_8 ));
    Odrv12 I__5633 (
            .O(N__27887),
            .I(\b2v_inst36.countZ0Z_8 ));
    Odrv4 I__5632 (
            .O(N__27884),
            .I(\b2v_inst36.countZ0Z_8 ));
    InMux I__5631 (
            .O(N__27877),
            .I(N__27873));
    InMux I__5630 (
            .O(N__27876),
            .I(N__27870));
    LocalMux I__5629 (
            .O(N__27873),
            .I(N__27865));
    LocalMux I__5628 (
            .O(N__27870),
            .I(N__27865));
    Span4Mux_h I__5627 (
            .O(N__27865),
            .I(N__27862));
    Odrv4 I__5626 (
            .O(N__27862),
            .I(\b2v_inst36.un2_count_1_cry_7_THRU_CO ));
    CascadeMux I__5625 (
            .O(N__27859),
            .I(\b2v_inst36.countZ0Z_8_cascade_ ));
    InMux I__5624 (
            .O(N__27856),
            .I(N__27853));
    LocalMux I__5623 (
            .O(N__27853),
            .I(\b2v_inst36.count_2_8 ));
    InMux I__5622 (
            .O(N__27850),
            .I(N__27844));
    InMux I__5621 (
            .O(N__27849),
            .I(N__27844));
    LocalMux I__5620 (
            .O(N__27844),
            .I(\b2v_inst36.un2_count_1_cry_1_THRU_CO ));
    InMux I__5619 (
            .O(N__27841),
            .I(\b2v_inst36.un2_count_1_cry_1 ));
    InMux I__5618 (
            .O(N__27838),
            .I(\b2v_inst36.un2_count_1_cry_2 ));
    InMux I__5617 (
            .O(N__27835),
            .I(N__27831));
    InMux I__5616 (
            .O(N__27834),
            .I(N__27828));
    LocalMux I__5615 (
            .O(N__27831),
            .I(N__27825));
    LocalMux I__5614 (
            .O(N__27828),
            .I(\b2v_inst36.countZ0Z_4 ));
    Odrv12 I__5613 (
            .O(N__27825),
            .I(\b2v_inst36.countZ0Z_4 ));
    InMux I__5612 (
            .O(N__27820),
            .I(N__27814));
    InMux I__5611 (
            .O(N__27819),
            .I(N__27814));
    LocalMux I__5610 (
            .O(N__27814),
            .I(N__27811));
    Odrv4 I__5609 (
            .O(N__27811),
            .I(\b2v_inst36.count_rst_10 ));
    InMux I__5608 (
            .O(N__27808),
            .I(\b2v_inst36.un2_count_1_cry_3 ));
    InMux I__5607 (
            .O(N__27805),
            .I(\b2v_inst36.un2_count_1_cry_4 ));
    InMux I__5606 (
            .O(N__27802),
            .I(N__27798));
    InMux I__5605 (
            .O(N__27801),
            .I(N__27795));
    LocalMux I__5604 (
            .O(N__27798),
            .I(N__27790));
    LocalMux I__5603 (
            .O(N__27795),
            .I(N__27790));
    Odrv4 I__5602 (
            .O(N__27790),
            .I(\b2v_inst36.countZ0Z_6 ));
    InMux I__5601 (
            .O(N__27787),
            .I(N__27781));
    InMux I__5600 (
            .O(N__27786),
            .I(N__27781));
    LocalMux I__5599 (
            .O(N__27781),
            .I(N__27778));
    Odrv12 I__5598 (
            .O(N__27778),
            .I(\b2v_inst36.count_rst_8 ));
    InMux I__5597 (
            .O(N__27775),
            .I(\b2v_inst36.un2_count_1_cry_5 ));
    InMux I__5596 (
            .O(N__27772),
            .I(\b2v_inst36.un2_count_1_cry_6 ));
    InMux I__5595 (
            .O(N__27769),
            .I(\b2v_inst36.un2_count_1_cry_7 ));
    InMux I__5594 (
            .O(N__27766),
            .I(N__27763));
    LocalMux I__5593 (
            .O(N__27763),
            .I(N__27759));
    InMux I__5592 (
            .O(N__27762),
            .I(N__27756));
    Span4Mux_h I__5591 (
            .O(N__27759),
            .I(N__27753));
    LocalMux I__5590 (
            .O(N__27756),
            .I(\b2v_inst36.countZ0Z_9 ));
    Odrv4 I__5589 (
            .O(N__27753),
            .I(\b2v_inst36.countZ0Z_9 ));
    InMux I__5588 (
            .O(N__27748),
            .I(N__27744));
    InMux I__5587 (
            .O(N__27747),
            .I(N__27741));
    LocalMux I__5586 (
            .O(N__27744),
            .I(N__27736));
    LocalMux I__5585 (
            .O(N__27741),
            .I(N__27736));
    Span4Mux_s1_v I__5584 (
            .O(N__27736),
            .I(N__27733));
    Odrv4 I__5583 (
            .O(N__27733),
            .I(\b2v_inst36.count_rst_5 ));
    InMux I__5582 (
            .O(N__27730),
            .I(bfn_9_2_0_));
    InMux I__5581 (
            .O(N__27727),
            .I(\b2v_inst36.un2_count_1_cry_9 ));
    InMux I__5580 (
            .O(N__27724),
            .I(N__27715));
    InMux I__5579 (
            .O(N__27723),
            .I(N__27711));
    InMux I__5578 (
            .O(N__27722),
            .I(N__27707));
    InMux I__5577 (
            .O(N__27721),
            .I(N__27702));
    InMux I__5576 (
            .O(N__27720),
            .I(N__27702));
    InMux I__5575 (
            .O(N__27719),
            .I(N__27695));
    InMux I__5574 (
            .O(N__27718),
            .I(N__27695));
    LocalMux I__5573 (
            .O(N__27715),
            .I(N__27692));
    CascadeMux I__5572 (
            .O(N__27714),
            .I(N__27689));
    LocalMux I__5571 (
            .O(N__27711),
            .I(N__27684));
    InMux I__5570 (
            .O(N__27710),
            .I(N__27681));
    LocalMux I__5569 (
            .O(N__27707),
            .I(N__27676));
    LocalMux I__5568 (
            .O(N__27702),
            .I(N__27676));
    CascadeMux I__5567 (
            .O(N__27701),
            .I(N__27673));
    CascadeMux I__5566 (
            .O(N__27700),
            .I(N__27665));
    LocalMux I__5565 (
            .O(N__27695),
            .I(N__27660));
    Span4Mux_h I__5564 (
            .O(N__27692),
            .I(N__27654));
    InMux I__5563 (
            .O(N__27689),
            .I(N__27651));
    InMux I__5562 (
            .O(N__27688),
            .I(N__27646));
    InMux I__5561 (
            .O(N__27687),
            .I(N__27646));
    Span4Mux_h I__5560 (
            .O(N__27684),
            .I(N__27639));
    LocalMux I__5559 (
            .O(N__27681),
            .I(N__27639));
    Span4Mux_h I__5558 (
            .O(N__27676),
            .I(N__27639));
    InMux I__5557 (
            .O(N__27673),
            .I(N__27634));
    InMux I__5556 (
            .O(N__27672),
            .I(N__27634));
    InMux I__5555 (
            .O(N__27671),
            .I(N__27629));
    InMux I__5554 (
            .O(N__27670),
            .I(N__27629));
    InMux I__5553 (
            .O(N__27669),
            .I(N__27624));
    InMux I__5552 (
            .O(N__27668),
            .I(N__27624));
    InMux I__5551 (
            .O(N__27665),
            .I(N__27617));
    InMux I__5550 (
            .O(N__27664),
            .I(N__27617));
    InMux I__5549 (
            .O(N__27663),
            .I(N__27617));
    Span4Mux_h I__5548 (
            .O(N__27660),
            .I(N__27614));
    InMux I__5547 (
            .O(N__27659),
            .I(N__27607));
    InMux I__5546 (
            .O(N__27658),
            .I(N__27607));
    InMux I__5545 (
            .O(N__27657),
            .I(N__27607));
    Span4Mux_v I__5544 (
            .O(N__27654),
            .I(N__27604));
    LocalMux I__5543 (
            .O(N__27651),
            .I(N__27596));
    LocalMux I__5542 (
            .O(N__27646),
            .I(N__27596));
    Span4Mux_v I__5541 (
            .O(N__27639),
            .I(N__27596));
    LocalMux I__5540 (
            .O(N__27634),
            .I(N__27586));
    LocalMux I__5539 (
            .O(N__27629),
            .I(N__27586));
    LocalMux I__5538 (
            .O(N__27624),
            .I(N__27586));
    LocalMux I__5537 (
            .O(N__27617),
            .I(N__27586));
    Span4Mux_v I__5536 (
            .O(N__27614),
            .I(N__27581));
    LocalMux I__5535 (
            .O(N__27607),
            .I(N__27581));
    Span4Mux_v I__5534 (
            .O(N__27604),
            .I(N__27578));
    IoInMux I__5533 (
            .O(N__27603),
            .I(N__27575));
    Span4Mux_v I__5532 (
            .O(N__27596),
            .I(N__27572));
    InMux I__5531 (
            .O(N__27595),
            .I(N__27569));
    Span4Mux_v I__5530 (
            .O(N__27586),
            .I(N__27564));
    Span4Mux_h I__5529 (
            .O(N__27581),
            .I(N__27564));
    Odrv4 I__5528 (
            .O(N__27578),
            .I(G_146));
    LocalMux I__5527 (
            .O(N__27575),
            .I(G_146));
    Odrv4 I__5526 (
            .O(N__27572),
            .I(G_146));
    LocalMux I__5525 (
            .O(N__27569),
            .I(G_146));
    Odrv4 I__5524 (
            .O(N__27564),
            .I(G_146));
    InMux I__5523 (
            .O(N__27553),
            .I(N__27549));
    InMux I__5522 (
            .O(N__27552),
            .I(N__27546));
    LocalMux I__5521 (
            .O(N__27549),
            .I(N__27543));
    LocalMux I__5520 (
            .O(N__27546),
            .I(N__27538));
    Span4Mux_h I__5519 (
            .O(N__27543),
            .I(N__27538));
    Odrv4 I__5518 (
            .O(N__27538),
            .I(N_15_i_0_a4_1));
    InMux I__5517 (
            .O(N__27535),
            .I(N__27531));
    InMux I__5516 (
            .O(N__27534),
            .I(N__27528));
    LocalMux I__5515 (
            .O(N__27531),
            .I(N__27525));
    LocalMux I__5514 (
            .O(N__27528),
            .I(N__27522));
    Span4Mux_h I__5513 (
            .O(N__27525),
            .I(N__27519));
    Span4Mux_h I__5512 (
            .O(N__27522),
            .I(N__27516));
    Odrv4 I__5511 (
            .O(N__27519),
            .I(N_73_mux_i_i_a7_0_0));
    Odrv4 I__5510 (
            .O(N__27516),
            .I(N_73_mux_i_i_a7_0_0));
    InMux I__5509 (
            .O(N__27511),
            .I(N__27505));
    InMux I__5508 (
            .O(N__27510),
            .I(N__27505));
    LocalMux I__5507 (
            .O(N__27505),
            .I(N__27502));
    Odrv4 I__5506 (
            .O(N__27502),
            .I(\b2v_inst11.count_1_8 ));
    InMux I__5505 (
            .O(N__27499),
            .I(N__27496));
    LocalMux I__5504 (
            .O(N__27496),
            .I(\b2v_inst11.count_0_8 ));
    InMux I__5503 (
            .O(N__27493),
            .I(N__27490));
    LocalMux I__5502 (
            .O(N__27490),
            .I(N__27487));
    Odrv4 I__5501 (
            .O(N__27487),
            .I(\b2v_inst11.g0_2_1 ));
    InMux I__5500 (
            .O(N__27484),
            .I(N__27480));
    InMux I__5499 (
            .O(N__27483),
            .I(N__27477));
    LocalMux I__5498 (
            .O(N__27480),
            .I(\b2v_inst11.pwm_outZ0 ));
    LocalMux I__5497 (
            .O(N__27477),
            .I(\b2v_inst11.pwm_outZ0 ));
    SRMux I__5496 (
            .O(N__27472),
            .I(N__27469));
    LocalMux I__5495 (
            .O(N__27469),
            .I(N__27466));
    Odrv12 I__5494 (
            .O(N__27466),
            .I(\b2v_inst11.pwm_out_1_sqmuxa ));
    CascadeMux I__5493 (
            .O(N__27463),
            .I(\b2v_inst11.curr_state_3_0_cascade_ ));
    CascadeMux I__5492 (
            .O(N__27460),
            .I(\b2v_inst11.curr_stateZ0Z_0_cascade_ ));
    InMux I__5491 (
            .O(N__27457),
            .I(N__27441));
    InMux I__5490 (
            .O(N__27456),
            .I(N__27441));
    InMux I__5489 (
            .O(N__27455),
            .I(N__27441));
    InMux I__5488 (
            .O(N__27454),
            .I(N__27430));
    InMux I__5487 (
            .O(N__27453),
            .I(N__27430));
    InMux I__5486 (
            .O(N__27452),
            .I(N__27430));
    InMux I__5485 (
            .O(N__27451),
            .I(N__27421));
    InMux I__5484 (
            .O(N__27450),
            .I(N__27421));
    InMux I__5483 (
            .O(N__27449),
            .I(N__27421));
    InMux I__5482 (
            .O(N__27448),
            .I(N__27421));
    LocalMux I__5481 (
            .O(N__27441),
            .I(N__27415));
    InMux I__5480 (
            .O(N__27440),
            .I(N__27406));
    InMux I__5479 (
            .O(N__27439),
            .I(N__27406));
    InMux I__5478 (
            .O(N__27438),
            .I(N__27406));
    InMux I__5477 (
            .O(N__27437),
            .I(N__27406));
    LocalMux I__5476 (
            .O(N__27430),
            .I(N__27403));
    LocalMux I__5475 (
            .O(N__27421),
            .I(N__27400));
    InMux I__5474 (
            .O(N__27420),
            .I(N__27395));
    InMux I__5473 (
            .O(N__27419),
            .I(N__27395));
    InMux I__5472 (
            .O(N__27418),
            .I(N__27392));
    Span4Mux_h I__5471 (
            .O(N__27415),
            .I(N__27389));
    LocalMux I__5470 (
            .O(N__27406),
            .I(N__27382));
    Span4Mux_h I__5469 (
            .O(N__27403),
            .I(N__27382));
    Span4Mux_h I__5468 (
            .O(N__27400),
            .I(N__27382));
    LocalMux I__5467 (
            .O(N__27395),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    LocalMux I__5466 (
            .O(N__27392),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__5465 (
            .O(N__27389),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    Odrv4 I__5464 (
            .O(N__27382),
            .I(\b2v_inst11.count_0_sqmuxa_i ));
    CascadeMux I__5463 (
            .O(N__27373),
            .I(\b2v_inst11.count_0_sqmuxa_i_cascade_ ));
    InMux I__5462 (
            .O(N__27370),
            .I(N__27367));
    LocalMux I__5461 (
            .O(N__27367),
            .I(\b2v_inst11.count_1_0 ));
    InMux I__5460 (
            .O(N__27364),
            .I(N__27360));
    InMux I__5459 (
            .O(N__27363),
            .I(N__27357));
    LocalMux I__5458 (
            .O(N__27360),
            .I(\b2v_inst36.un2_count_1_axb_1 ));
    LocalMux I__5457 (
            .O(N__27357),
            .I(\b2v_inst36.un2_count_1_axb_1 ));
    CascadeMux I__5456 (
            .O(N__27352),
            .I(N__27345));
    InMux I__5455 (
            .O(N__27351),
            .I(N__27340));
    InMux I__5454 (
            .O(N__27350),
            .I(N__27340));
    InMux I__5453 (
            .O(N__27349),
            .I(N__27335));
    InMux I__5452 (
            .O(N__27348),
            .I(N__27335));
    InMux I__5451 (
            .O(N__27345),
            .I(N__27332));
    LocalMux I__5450 (
            .O(N__27340),
            .I(\b2v_inst36.countZ0Z_0 ));
    LocalMux I__5449 (
            .O(N__27335),
            .I(\b2v_inst36.countZ0Z_0 ));
    LocalMux I__5448 (
            .O(N__27332),
            .I(\b2v_inst36.countZ0Z_0 ));
    InMux I__5447 (
            .O(N__27325),
            .I(N__27322));
    LocalMux I__5446 (
            .O(N__27322),
            .I(\b2v_inst11.un79_clk_100khzlt6 ));
    CascadeMux I__5445 (
            .O(N__27319),
            .I(\b2v_inst11.un79_clk_100khzlto15_4_cascade_ ));
    InMux I__5444 (
            .O(N__27316),
            .I(N__27313));
    LocalMux I__5443 (
            .O(N__27313),
            .I(\b2v_inst11.un79_clk_100khzlto15_7 ));
    CascadeMux I__5442 (
            .O(N__27310),
            .I(\b2v_inst11.count_RNIZ0Z_13_cascade_ ));
    CascadeMux I__5441 (
            .O(N__27307),
            .I(\b2v_inst11.countZ0Z_0_cascade_ ));
    CascadeMux I__5440 (
            .O(N__27304),
            .I(\b2v_inst11.count_1_1_cascade_ ));
    CascadeMux I__5439 (
            .O(N__27301),
            .I(\b2v_inst11.countZ0Z_1_cascade_ ));
    InMux I__5438 (
            .O(N__27298),
            .I(N__27295));
    LocalMux I__5437 (
            .O(N__27295),
            .I(\b2v_inst11.count_0_1 ));
    InMux I__5436 (
            .O(N__27292),
            .I(N__27289));
    LocalMux I__5435 (
            .O(N__27289),
            .I(\b2v_inst11.count_0_0 ));
    InMux I__5434 (
            .O(N__27286),
            .I(N__27282));
    CascadeMux I__5433 (
            .O(N__27285),
            .I(N__27279));
    LocalMux I__5432 (
            .O(N__27282),
            .I(N__27276));
    InMux I__5431 (
            .O(N__27279),
            .I(N__27273));
    Span4Mux_h I__5430 (
            .O(N__27276),
            .I(N__27268));
    LocalMux I__5429 (
            .O(N__27273),
            .I(N__27268));
    Span4Mux_v I__5428 (
            .O(N__27268),
            .I(N__27265));
    Span4Mux_h I__5427 (
            .O(N__27265),
            .I(N__27262));
    Span4Mux_v I__5426 (
            .O(N__27262),
            .I(N__27259));
    Odrv4 I__5425 (
            .O(N__27259),
            .I(b2v_inst11_dutycycle_set_1));
    CascadeMux I__5424 (
            .O(N__27256),
            .I(N__27253));
    InMux I__5423 (
            .O(N__27253),
            .I(N__27247));
    InMux I__5422 (
            .O(N__27252),
            .I(N__27247));
    LocalMux I__5421 (
            .O(N__27247),
            .I(\b2v_inst11.count_1_3 ));
    InMux I__5420 (
            .O(N__27244),
            .I(N__27241));
    LocalMux I__5419 (
            .O(N__27241),
            .I(\b2v_inst11.count_0_3 ));
    CascadeMux I__5418 (
            .O(N__27238),
            .I(N__27235));
    InMux I__5417 (
            .O(N__27235),
            .I(N__27229));
    InMux I__5416 (
            .O(N__27234),
            .I(N__27229));
    LocalMux I__5415 (
            .O(N__27229),
            .I(\b2v_inst11.count_1_13 ));
    InMux I__5414 (
            .O(N__27226),
            .I(N__27223));
    LocalMux I__5413 (
            .O(N__27223),
            .I(\b2v_inst11.count_0_13 ));
    CascadeMux I__5412 (
            .O(N__27220),
            .I(N__27217));
    InMux I__5411 (
            .O(N__27217),
            .I(N__27211));
    InMux I__5410 (
            .O(N__27216),
            .I(N__27211));
    LocalMux I__5409 (
            .O(N__27211),
            .I(\b2v_inst11.count_1_4 ));
    InMux I__5408 (
            .O(N__27208),
            .I(N__27205));
    LocalMux I__5407 (
            .O(N__27205),
            .I(\b2v_inst11.count_0_4 ));
    CascadeMux I__5406 (
            .O(N__27202),
            .I(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ));
    InMux I__5405 (
            .O(N__27199),
            .I(N__27196));
    LocalMux I__5404 (
            .O(N__27196),
            .I(N__27193));
    Span4Mux_v I__5403 (
            .O(N__27193),
            .I(N__27190));
    Odrv4 I__5402 (
            .O(N__27190),
            .I(\b2v_inst11.g2_0_0 ));
    InMux I__5401 (
            .O(N__27187),
            .I(N__27184));
    LocalMux I__5400 (
            .O(N__27184),
            .I(b2v_inst11_un1_dutycycle_164_0));
    CascadeMux I__5399 (
            .O(N__27181),
            .I(N__27178));
    InMux I__5398 (
            .O(N__27178),
            .I(N__27172));
    InMux I__5397 (
            .O(N__27177),
            .I(N__27172));
    LocalMux I__5396 (
            .O(N__27172),
            .I(N__27169));
    Odrv12 I__5395 (
            .O(N__27169),
            .I(\b2v_inst5.N_6 ));
    CascadeMux I__5394 (
            .O(N__27166),
            .I(b2v_inst11_un1_dutycycle_164_0_cascade_));
    InMux I__5393 (
            .O(N__27163),
            .I(N__27160));
    LocalMux I__5392 (
            .O(N__27160),
            .I(N__27157));
    Span4Mux_h I__5391 (
            .O(N__27157),
            .I(N__27154));
    Odrv4 I__5390 (
            .O(N__27154),
            .I(\b2v_inst5.N_13 ));
    CascadeMux I__5389 (
            .O(N__27151),
            .I(N__27143));
    CascadeMux I__5388 (
            .O(N__27150),
            .I(N__27139));
    CascadeMux I__5387 (
            .O(N__27149),
            .I(N__27136));
    CascadeMux I__5386 (
            .O(N__27148),
            .I(N__27133));
    InMux I__5385 (
            .O(N__27147),
            .I(N__27126));
    CascadeMux I__5384 (
            .O(N__27146),
            .I(N__27123));
    InMux I__5383 (
            .O(N__27143),
            .I(N__27120));
    InMux I__5382 (
            .O(N__27142),
            .I(N__27117));
    InMux I__5381 (
            .O(N__27139),
            .I(N__27114));
    InMux I__5380 (
            .O(N__27136),
            .I(N__27109));
    InMux I__5379 (
            .O(N__27133),
            .I(N__27109));
    CascadeMux I__5378 (
            .O(N__27132),
            .I(N__27105));
    CascadeMux I__5377 (
            .O(N__27131),
            .I(N__27097));
    CascadeMux I__5376 (
            .O(N__27130),
            .I(N__27093));
    CascadeMux I__5375 (
            .O(N__27129),
            .I(N__27089));
    LocalMux I__5374 (
            .O(N__27126),
            .I(N__27085));
    InMux I__5373 (
            .O(N__27123),
            .I(N__27082));
    LocalMux I__5372 (
            .O(N__27120),
            .I(N__27079));
    LocalMux I__5371 (
            .O(N__27117),
            .I(N__27075));
    LocalMux I__5370 (
            .O(N__27114),
            .I(N__27070));
    LocalMux I__5369 (
            .O(N__27109),
            .I(N__27070));
    InMux I__5368 (
            .O(N__27108),
            .I(N__27065));
    InMux I__5367 (
            .O(N__27105),
            .I(N__27065));
    CascadeMux I__5366 (
            .O(N__27104),
            .I(N__27060));
    CascadeMux I__5365 (
            .O(N__27103),
            .I(N__27055));
    InMux I__5364 (
            .O(N__27102),
            .I(N__27051));
    InMux I__5363 (
            .O(N__27101),
            .I(N__27034));
    InMux I__5362 (
            .O(N__27100),
            .I(N__27034));
    InMux I__5361 (
            .O(N__27097),
            .I(N__27034));
    InMux I__5360 (
            .O(N__27096),
            .I(N__27034));
    InMux I__5359 (
            .O(N__27093),
            .I(N__27034));
    InMux I__5358 (
            .O(N__27092),
            .I(N__27034));
    InMux I__5357 (
            .O(N__27089),
            .I(N__27034));
    InMux I__5356 (
            .O(N__27088),
            .I(N__27034));
    Span4Mux_v I__5355 (
            .O(N__27085),
            .I(N__27029));
    LocalMux I__5354 (
            .O(N__27082),
            .I(N__27029));
    Span4Mux_v I__5353 (
            .O(N__27079),
            .I(N__27026));
    InMux I__5352 (
            .O(N__27078),
            .I(N__27023));
    Span4Mux_v I__5351 (
            .O(N__27075),
            .I(N__27018));
    Span4Mux_v I__5350 (
            .O(N__27070),
            .I(N__27018));
    LocalMux I__5349 (
            .O(N__27065),
            .I(N__27015));
    InMux I__5348 (
            .O(N__27064),
            .I(N__27010));
    InMux I__5347 (
            .O(N__27063),
            .I(N__27010));
    InMux I__5346 (
            .O(N__27060),
            .I(N__26999));
    InMux I__5345 (
            .O(N__27059),
            .I(N__26999));
    InMux I__5344 (
            .O(N__27058),
            .I(N__26999));
    InMux I__5343 (
            .O(N__27055),
            .I(N__26999));
    InMux I__5342 (
            .O(N__27054),
            .I(N__26999));
    LocalMux I__5341 (
            .O(N__27051),
            .I(N__26992));
    LocalMux I__5340 (
            .O(N__27034),
            .I(N__26992));
    Span4Mux_v I__5339 (
            .O(N__27029),
            .I(N__26992));
    Odrv4 I__5338 (
            .O(N__27026),
            .I(\b2v_inst11.N_3060_i ));
    LocalMux I__5337 (
            .O(N__27023),
            .I(\b2v_inst11.N_3060_i ));
    Odrv4 I__5336 (
            .O(N__27018),
            .I(\b2v_inst11.N_3060_i ));
    Odrv4 I__5335 (
            .O(N__27015),
            .I(\b2v_inst11.N_3060_i ));
    LocalMux I__5334 (
            .O(N__27010),
            .I(\b2v_inst11.N_3060_i ));
    LocalMux I__5333 (
            .O(N__26999),
            .I(\b2v_inst11.N_3060_i ));
    Odrv4 I__5332 (
            .O(N__26992),
            .I(\b2v_inst11.N_3060_i ));
    InMux I__5331 (
            .O(N__26977),
            .I(N__26971));
    InMux I__5330 (
            .O(N__26976),
            .I(N__26971));
    LocalMux I__5329 (
            .O(N__26971),
            .I(N__26968));
    Span4Mux_h I__5328 (
            .O(N__26968),
            .I(N__26965));
    Odrv4 I__5327 (
            .O(N__26965),
            .I(\b2v_inst11.un1_dutycycle_96_0_a3_1 ));
    InMux I__5326 (
            .O(N__26962),
            .I(N__26959));
    LocalMux I__5325 (
            .O(N__26959),
            .I(N__26956));
    Span4Mux_h I__5324 (
            .O(N__26956),
            .I(N__26953));
    Span4Mux_v I__5323 (
            .O(N__26953),
            .I(N__26950));
    Odrv4 I__5322 (
            .O(N__26950),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_7 ));
    CascadeMux I__5321 (
            .O(N__26947),
            .I(N__26944));
    InMux I__5320 (
            .O(N__26944),
            .I(N__26938));
    InMux I__5319 (
            .O(N__26943),
            .I(N__26935));
    InMux I__5318 (
            .O(N__26942),
            .I(N__26932));
    InMux I__5317 (
            .O(N__26941),
            .I(N__26928));
    LocalMux I__5316 (
            .O(N__26938),
            .I(N__26925));
    LocalMux I__5315 (
            .O(N__26935),
            .I(N__26922));
    LocalMux I__5314 (
            .O(N__26932),
            .I(N__26919));
    CascadeMux I__5313 (
            .O(N__26931),
            .I(N__26916));
    LocalMux I__5312 (
            .O(N__26928),
            .I(N__26912));
    Span4Mux_v I__5311 (
            .O(N__26925),
            .I(N__26909));
    Span4Mux_h I__5310 (
            .O(N__26922),
            .I(N__26904));
    Span4Mux_v I__5309 (
            .O(N__26919),
            .I(N__26904));
    InMux I__5308 (
            .O(N__26916),
            .I(N__26899));
    InMux I__5307 (
            .O(N__26915),
            .I(N__26899));
    Span4Mux_h I__5306 (
            .O(N__26912),
            .I(N__26896));
    Odrv4 I__5305 (
            .O(N__26909),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__5304 (
            .O(N__26904),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    LocalMux I__5303 (
            .O(N__26899),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__5302 (
            .O(N__26896),
            .I(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    CascadeMux I__5301 (
            .O(N__26887),
            .I(N__26883));
    InMux I__5300 (
            .O(N__26886),
            .I(N__26880));
    InMux I__5299 (
            .O(N__26883),
            .I(N__26877));
    LocalMux I__5298 (
            .O(N__26880),
            .I(N__26873));
    LocalMux I__5297 (
            .O(N__26877),
            .I(N__26870));
    InMux I__5296 (
            .O(N__26876),
            .I(N__26867));
    Span4Mux_v I__5295 (
            .O(N__26873),
            .I(N__26864));
    Span4Mux_h I__5294 (
            .O(N__26870),
            .I(N__26861));
    LocalMux I__5293 (
            .O(N__26867),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5 ));
    Odrv4 I__5292 (
            .O(N__26864),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5 ));
    Odrv4 I__5291 (
            .O(N__26861),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5 ));
    InMux I__5290 (
            .O(N__26854),
            .I(N__26848));
    InMux I__5289 (
            .O(N__26853),
            .I(N__26848));
    LocalMux I__5288 (
            .O(N__26848),
            .I(N_73_mux_i_i_o3_1_1));
    CascadeMux I__5287 (
            .O(N__26845),
            .I(N__26839));
    CascadeMux I__5286 (
            .O(N__26844),
            .I(N__26827));
    CascadeMux I__5285 (
            .O(N__26843),
            .I(N__26824));
    CascadeMux I__5284 (
            .O(N__26842),
            .I(N__26820));
    InMux I__5283 (
            .O(N__26839),
            .I(N__26817));
    InMux I__5282 (
            .O(N__26838),
            .I(N__26812));
    InMux I__5281 (
            .O(N__26837),
            .I(N__26812));
    CascadeMux I__5280 (
            .O(N__26836),
            .I(N__26809));
    InMux I__5279 (
            .O(N__26835),
            .I(N__26801));
    InMux I__5278 (
            .O(N__26834),
            .I(N__26801));
    InMux I__5277 (
            .O(N__26833),
            .I(N__26801));
    CascadeMux I__5276 (
            .O(N__26832),
            .I(N__26795));
    CascadeMux I__5275 (
            .O(N__26831),
            .I(N__26792));
    InMux I__5274 (
            .O(N__26830),
            .I(N__26784));
    InMux I__5273 (
            .O(N__26827),
            .I(N__26784));
    InMux I__5272 (
            .O(N__26824),
            .I(N__26781));
    CascadeMux I__5271 (
            .O(N__26823),
            .I(N__26778));
    InMux I__5270 (
            .O(N__26820),
            .I(N__26773));
    LocalMux I__5269 (
            .O(N__26817),
            .I(N__26768));
    LocalMux I__5268 (
            .O(N__26812),
            .I(N__26768));
    InMux I__5267 (
            .O(N__26809),
            .I(N__26763));
    InMux I__5266 (
            .O(N__26808),
            .I(N__26763));
    LocalMux I__5265 (
            .O(N__26801),
            .I(N__26760));
    InMux I__5264 (
            .O(N__26800),
            .I(N__26751));
    InMux I__5263 (
            .O(N__26799),
            .I(N__26751));
    InMux I__5262 (
            .O(N__26798),
            .I(N__26751));
    InMux I__5261 (
            .O(N__26795),
            .I(N__26751));
    InMux I__5260 (
            .O(N__26792),
            .I(N__26745));
    InMux I__5259 (
            .O(N__26791),
            .I(N__26745));
    InMux I__5258 (
            .O(N__26790),
            .I(N__26740));
    InMux I__5257 (
            .O(N__26789),
            .I(N__26740));
    LocalMux I__5256 (
            .O(N__26784),
            .I(N__26737));
    LocalMux I__5255 (
            .O(N__26781),
            .I(N__26734));
    InMux I__5254 (
            .O(N__26778),
            .I(N__26731));
    InMux I__5253 (
            .O(N__26777),
            .I(N__26726));
    InMux I__5252 (
            .O(N__26776),
            .I(N__26726));
    LocalMux I__5251 (
            .O(N__26773),
            .I(N__26723));
    Span4Mux_v I__5250 (
            .O(N__26768),
            .I(N__26718));
    LocalMux I__5249 (
            .O(N__26763),
            .I(N__26718));
    Span4Mux_h I__5248 (
            .O(N__26760),
            .I(N__26713));
    LocalMux I__5247 (
            .O(N__26751),
            .I(N__26713));
    CascadeMux I__5246 (
            .O(N__26750),
            .I(N__26709));
    LocalMux I__5245 (
            .O(N__26745),
            .I(N__26706));
    LocalMux I__5244 (
            .O(N__26740),
            .I(N__26703));
    Span4Mux_h I__5243 (
            .O(N__26737),
            .I(N__26700));
    Span4Mux_v I__5242 (
            .O(N__26734),
            .I(N__26693));
    LocalMux I__5241 (
            .O(N__26731),
            .I(N__26693));
    LocalMux I__5240 (
            .O(N__26726),
            .I(N__26693));
    Span4Mux_h I__5239 (
            .O(N__26723),
            .I(N__26688));
    Span4Mux_h I__5238 (
            .O(N__26718),
            .I(N__26688));
    Span4Mux_v I__5237 (
            .O(N__26713),
            .I(N__26685));
    InMux I__5236 (
            .O(N__26712),
            .I(N__26680));
    InMux I__5235 (
            .O(N__26709),
            .I(N__26680));
    Odrv12 I__5234 (
            .O(N__26706),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__5233 (
            .O(N__26703),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__5232 (
            .O(N__26700),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__5231 (
            .O(N__26693),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__5230 (
            .O(N__26688),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    Odrv4 I__5229 (
            .O(N__26685),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    LocalMux I__5228 (
            .O(N__26680),
            .I(\b2v_inst11.dutycycleZ1Z_3 ));
    CascadeMux I__5227 (
            .O(N__26665),
            .I(N__26662));
    InMux I__5226 (
            .O(N__26662),
            .I(N__26659));
    LocalMux I__5225 (
            .O(N__26659),
            .I(N__26656));
    Span4Mux_h I__5224 (
            .O(N__26656),
            .I(N__26653));
    Odrv4 I__5223 (
            .O(N__26653),
            .I(\b2v_inst11.g3_0_1 ));
    InMux I__5222 (
            .O(N__26650),
            .I(N__26638));
    InMux I__5221 (
            .O(N__26649),
            .I(N__26629));
    InMux I__5220 (
            .O(N__26648),
            .I(N__26626));
    InMux I__5219 (
            .O(N__26647),
            .I(N__26623));
    InMux I__5218 (
            .O(N__26646),
            .I(N__26616));
    InMux I__5217 (
            .O(N__26645),
            .I(N__26616));
    InMux I__5216 (
            .O(N__26644),
            .I(N__26616));
    InMux I__5215 (
            .O(N__26643),
            .I(N__26613));
    InMux I__5214 (
            .O(N__26642),
            .I(N__26608));
    CascadeMux I__5213 (
            .O(N__26641),
            .I(N__26605));
    LocalMux I__5212 (
            .O(N__26638),
            .I(N__26602));
    InMux I__5211 (
            .O(N__26637),
            .I(N__26597));
    InMux I__5210 (
            .O(N__26636),
            .I(N__26597));
    InMux I__5209 (
            .O(N__26635),
            .I(N__26594));
    InMux I__5208 (
            .O(N__26634),
            .I(N__26591));
    CascadeMux I__5207 (
            .O(N__26633),
            .I(N__26588));
    InMux I__5206 (
            .O(N__26632),
            .I(N__26584));
    LocalMux I__5205 (
            .O(N__26629),
            .I(N__26579));
    LocalMux I__5204 (
            .O(N__26626),
            .I(N__26579));
    LocalMux I__5203 (
            .O(N__26623),
            .I(N__26576));
    LocalMux I__5202 (
            .O(N__26616),
            .I(N__26571));
    LocalMux I__5201 (
            .O(N__26613),
            .I(N__26571));
    InMux I__5200 (
            .O(N__26612),
            .I(N__26563));
    InMux I__5199 (
            .O(N__26611),
            .I(N__26563));
    LocalMux I__5198 (
            .O(N__26608),
            .I(N__26560));
    InMux I__5197 (
            .O(N__26605),
            .I(N__26557));
    Span4Mux_v I__5196 (
            .O(N__26602),
            .I(N__26552));
    LocalMux I__5195 (
            .O(N__26597),
            .I(N__26552));
    LocalMux I__5194 (
            .O(N__26594),
            .I(N__26547));
    LocalMux I__5193 (
            .O(N__26591),
            .I(N__26547));
    InMux I__5192 (
            .O(N__26588),
            .I(N__26542));
    InMux I__5191 (
            .O(N__26587),
            .I(N__26542));
    LocalMux I__5190 (
            .O(N__26584),
            .I(N__26539));
    Span4Mux_v I__5189 (
            .O(N__26579),
            .I(N__26534));
    Span4Mux_v I__5188 (
            .O(N__26576),
            .I(N__26534));
    Span4Mux_v I__5187 (
            .O(N__26571),
            .I(N__26531));
    InMux I__5186 (
            .O(N__26570),
            .I(N__26526));
    InMux I__5185 (
            .O(N__26569),
            .I(N__26526));
    InMux I__5184 (
            .O(N__26568),
            .I(N__26523));
    LocalMux I__5183 (
            .O(N__26563),
            .I(N__26520));
    Span4Mux_s3_v I__5182 (
            .O(N__26560),
            .I(N__26517));
    LocalMux I__5181 (
            .O(N__26557),
            .I(N__26508));
    Span4Mux_h I__5180 (
            .O(N__26552),
            .I(N__26508));
    Span4Mux_v I__5179 (
            .O(N__26547),
            .I(N__26508));
    LocalMux I__5178 (
            .O(N__26542),
            .I(N__26508));
    Span4Mux_v I__5177 (
            .O(N__26539),
            .I(N__26505));
    Sp12to4 I__5176 (
            .O(N__26534),
            .I(N__26496));
    Sp12to4 I__5175 (
            .O(N__26531),
            .I(N__26496));
    LocalMux I__5174 (
            .O(N__26526),
            .I(N__26496));
    LocalMux I__5173 (
            .O(N__26523),
            .I(N__26496));
    Span4Mux_v I__5172 (
            .O(N__26520),
            .I(N__26489));
    Span4Mux_h I__5171 (
            .O(N__26517),
            .I(N__26489));
    Span4Mux_h I__5170 (
            .O(N__26508),
            .I(N__26489));
    Odrv4 I__5169 (
            .O(N__26505),
            .I(\b2v_inst11.N_3038_i ));
    Odrv12 I__5168 (
            .O(N__26496),
            .I(\b2v_inst11.N_3038_i ));
    Odrv4 I__5167 (
            .O(N__26489),
            .I(\b2v_inst11.N_3038_i ));
    InMux I__5166 (
            .O(N__26482),
            .I(N__26478));
    InMux I__5165 (
            .O(N__26481),
            .I(N__26475));
    LocalMux I__5164 (
            .O(N__26478),
            .I(g3_0_4));
    LocalMux I__5163 (
            .O(N__26475),
            .I(g3_0_4));
    CascadeMux I__5162 (
            .O(N__26470),
            .I(N__26467));
    InMux I__5161 (
            .O(N__26467),
            .I(N__26461));
    InMux I__5160 (
            .O(N__26466),
            .I(N__26461));
    LocalMux I__5159 (
            .O(N__26461),
            .I(\b2v_inst11.count_1_12 ));
    InMux I__5158 (
            .O(N__26458),
            .I(N__26455));
    LocalMux I__5157 (
            .O(N__26455),
            .I(\b2v_inst11.count_0_12 ));
    InMux I__5156 (
            .O(N__26452),
            .I(N__26442));
    CascadeMux I__5155 (
            .O(N__26451),
            .I(N__26439));
    InMux I__5154 (
            .O(N__26450),
            .I(N__26427));
    InMux I__5153 (
            .O(N__26449),
            .I(N__26427));
    InMux I__5152 (
            .O(N__26448),
            .I(N__26422));
    InMux I__5151 (
            .O(N__26447),
            .I(N__26415));
    InMux I__5150 (
            .O(N__26446),
            .I(N__26415));
    InMux I__5149 (
            .O(N__26445),
            .I(N__26415));
    LocalMux I__5148 (
            .O(N__26442),
            .I(N__26412));
    InMux I__5147 (
            .O(N__26439),
            .I(N__26409));
    InMux I__5146 (
            .O(N__26438),
            .I(N__26406));
    InMux I__5145 (
            .O(N__26437),
            .I(N__26403));
    InMux I__5144 (
            .O(N__26436),
            .I(N__26398));
    InMux I__5143 (
            .O(N__26435),
            .I(N__26398));
    InMux I__5142 (
            .O(N__26434),
            .I(N__26391));
    InMux I__5141 (
            .O(N__26433),
            .I(N__26391));
    InMux I__5140 (
            .O(N__26432),
            .I(N__26391));
    LocalMux I__5139 (
            .O(N__26427),
            .I(N__26388));
    InMux I__5138 (
            .O(N__26426),
            .I(N__26383));
    InMux I__5137 (
            .O(N__26425),
            .I(N__26383));
    LocalMux I__5136 (
            .O(N__26422),
            .I(N__26380));
    LocalMux I__5135 (
            .O(N__26415),
            .I(N__26375));
    Span4Mux_h I__5134 (
            .O(N__26412),
            .I(N__26375));
    LocalMux I__5133 (
            .O(N__26409),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__5132 (
            .O(N__26406),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__5131 (
            .O(N__26403),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__5130 (
            .O(N__26398),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__5129 (
            .O(N__26391),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__5128 (
            .O(N__26388),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    LocalMux I__5127 (
            .O(N__26383),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__5126 (
            .O(N__26380),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    Odrv4 I__5125 (
            .O(N__26375),
            .I(\b2v_inst11.dutycycleZ0Z_1 ));
    InMux I__5124 (
            .O(N__26356),
            .I(N__26353));
    LocalMux I__5123 (
            .O(N__26353),
            .I(\b2v_inst11.un1_dutycycle_53_50_1_i_0_1 ));
    InMux I__5122 (
            .O(N__26350),
            .I(N__26347));
    LocalMux I__5121 (
            .O(N__26347),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_1 ));
    CascadeMux I__5120 (
            .O(N__26344),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_1_cascade_ ));
    CascadeMux I__5119 (
            .O(N__26341),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_3_cascade_ ));
    CascadeMux I__5118 (
            .O(N__26338),
            .I(N__26330));
    InMux I__5117 (
            .O(N__26337),
            .I(N__26323));
    CascadeMux I__5116 (
            .O(N__26336),
            .I(N__26320));
    InMux I__5115 (
            .O(N__26335),
            .I(N__26317));
    InMux I__5114 (
            .O(N__26334),
            .I(N__26310));
    InMux I__5113 (
            .O(N__26333),
            .I(N__26310));
    InMux I__5112 (
            .O(N__26330),
            .I(N__26310));
    InMux I__5111 (
            .O(N__26329),
            .I(N__26305));
    InMux I__5110 (
            .O(N__26328),
            .I(N__26302));
    CascadeMux I__5109 (
            .O(N__26327),
            .I(N__26296));
    InMux I__5108 (
            .O(N__26326),
            .I(N__26293));
    LocalMux I__5107 (
            .O(N__26323),
            .I(N__26290));
    InMux I__5106 (
            .O(N__26320),
            .I(N__26287));
    LocalMux I__5105 (
            .O(N__26317),
            .I(N__26284));
    LocalMux I__5104 (
            .O(N__26310),
            .I(N__26281));
    CascadeMux I__5103 (
            .O(N__26309),
            .I(N__26277));
    InMux I__5102 (
            .O(N__26308),
            .I(N__26272));
    LocalMux I__5101 (
            .O(N__26305),
            .I(N__26269));
    LocalMux I__5100 (
            .O(N__26302),
            .I(N__26266));
    InMux I__5099 (
            .O(N__26301),
            .I(N__26257));
    InMux I__5098 (
            .O(N__26300),
            .I(N__26257));
    InMux I__5097 (
            .O(N__26299),
            .I(N__26257));
    InMux I__5096 (
            .O(N__26296),
            .I(N__26257));
    LocalMux I__5095 (
            .O(N__26293),
            .I(N__26254));
    Span4Mux_v I__5094 (
            .O(N__26290),
            .I(N__26251));
    LocalMux I__5093 (
            .O(N__26287),
            .I(N__26244));
    Span4Mux_v I__5092 (
            .O(N__26284),
            .I(N__26244));
    Span4Mux_h I__5091 (
            .O(N__26281),
            .I(N__26244));
    InMux I__5090 (
            .O(N__26280),
            .I(N__26241));
    InMux I__5089 (
            .O(N__26277),
            .I(N__26238));
    InMux I__5088 (
            .O(N__26276),
            .I(N__26233));
    InMux I__5087 (
            .O(N__26275),
            .I(N__26233));
    LocalMux I__5086 (
            .O(N__26272),
            .I(N__26228));
    Span4Mux_h I__5085 (
            .O(N__26269),
            .I(N__26228));
    Span4Mux_h I__5084 (
            .O(N__26266),
            .I(N__26221));
    LocalMux I__5083 (
            .O(N__26257),
            .I(N__26221));
    Span4Mux_h I__5082 (
            .O(N__26254),
            .I(N__26221));
    Odrv4 I__5081 (
            .O(N__26251),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__5080 (
            .O(N__26244),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__5079 (
            .O(N__26241),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__5078 (
            .O(N__26238),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    LocalMux I__5077 (
            .O(N__26233),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__5076 (
            .O(N__26228),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    Odrv4 I__5075 (
            .O(N__26221),
            .I(\b2v_inst11.dutycycleZ0Z_5 ));
    InMux I__5074 (
            .O(N__26206),
            .I(N__26203));
    LocalMux I__5073 (
            .O(N__26203),
            .I(N__26200));
    Odrv4 I__5072 (
            .O(N__26200),
            .I(\b2v_inst11.m6_0_1 ));
    CascadeMux I__5071 (
            .O(N__26197),
            .I(N__26193));
    CascadeMux I__5070 (
            .O(N__26196),
            .I(N__26185));
    InMux I__5069 (
            .O(N__26193),
            .I(N__26180));
    InMux I__5068 (
            .O(N__26192),
            .I(N__26171));
    InMux I__5067 (
            .O(N__26191),
            .I(N__26171));
    InMux I__5066 (
            .O(N__26190),
            .I(N__26171));
    InMux I__5065 (
            .O(N__26189),
            .I(N__26168));
    InMux I__5064 (
            .O(N__26188),
            .I(N__26161));
    InMux I__5063 (
            .O(N__26185),
            .I(N__26158));
    InMux I__5062 (
            .O(N__26184),
            .I(N__26148));
    InMux I__5061 (
            .O(N__26183),
            .I(N__26148));
    LocalMux I__5060 (
            .O(N__26180),
            .I(N__26145));
    InMux I__5059 (
            .O(N__26179),
            .I(N__26140));
    InMux I__5058 (
            .O(N__26178),
            .I(N__26140));
    LocalMux I__5057 (
            .O(N__26171),
            .I(N__26137));
    LocalMux I__5056 (
            .O(N__26168),
            .I(N__26134));
    InMux I__5055 (
            .O(N__26167),
            .I(N__26125));
    InMux I__5054 (
            .O(N__26166),
            .I(N__26125));
    InMux I__5053 (
            .O(N__26165),
            .I(N__26125));
    InMux I__5052 (
            .O(N__26164),
            .I(N__26125));
    LocalMux I__5051 (
            .O(N__26161),
            .I(N__26122));
    LocalMux I__5050 (
            .O(N__26158),
            .I(N__26119));
    InMux I__5049 (
            .O(N__26157),
            .I(N__26116));
    InMux I__5048 (
            .O(N__26156),
            .I(N__26107));
    InMux I__5047 (
            .O(N__26155),
            .I(N__26107));
    InMux I__5046 (
            .O(N__26154),
            .I(N__26107));
    InMux I__5045 (
            .O(N__26153),
            .I(N__26107));
    LocalMux I__5044 (
            .O(N__26148),
            .I(N__26104));
    Span4Mux_v I__5043 (
            .O(N__26145),
            .I(N__26099));
    LocalMux I__5042 (
            .O(N__26140),
            .I(N__26096));
    Span4Mux_v I__5041 (
            .O(N__26137),
            .I(N__26087));
    Span4Mux_v I__5040 (
            .O(N__26134),
            .I(N__26087));
    LocalMux I__5039 (
            .O(N__26125),
            .I(N__26087));
    Span4Mux_v I__5038 (
            .O(N__26122),
            .I(N__26087));
    Span4Mux_v I__5037 (
            .O(N__26119),
            .I(N__26084));
    LocalMux I__5036 (
            .O(N__26116),
            .I(N__26077));
    LocalMux I__5035 (
            .O(N__26107),
            .I(N__26077));
    Span4Mux_h I__5034 (
            .O(N__26104),
            .I(N__26077));
    InMux I__5033 (
            .O(N__26103),
            .I(N__26072));
    InMux I__5032 (
            .O(N__26102),
            .I(N__26072));
    Odrv4 I__5031 (
            .O(N__26099),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv12 I__5030 (
            .O(N__26096),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5029 (
            .O(N__26087),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5028 (
            .O(N__26084),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    Odrv4 I__5027 (
            .O(N__26077),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    LocalMux I__5026 (
            .O(N__26072),
            .I(\b2v_inst11.dutycycleZ1Z_6 ));
    InMux I__5025 (
            .O(N__26059),
            .I(N__26056));
    LocalMux I__5024 (
            .O(N__26056),
            .I(\b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_0_1 ));
    InMux I__5023 (
            .O(N__26053),
            .I(N__26050));
    LocalMux I__5022 (
            .O(N__26050),
            .I(N__26047));
    Span4Mux_h I__5021 (
            .O(N__26047),
            .I(N__26044));
    Odrv4 I__5020 (
            .O(N__26044),
            .I(N_18));
    InMux I__5019 (
            .O(N__26041),
            .I(N__26038));
    LocalMux I__5018 (
            .O(N__26038),
            .I(\b2v_inst11.N_15_mux ));
    InMux I__5017 (
            .O(N__26035),
            .I(N__26032));
    LocalMux I__5016 (
            .O(N__26032),
            .I(\b2v_inst11.i6_mux_i_1 ));
    InMux I__5015 (
            .O(N__26029),
            .I(N__26026));
    LocalMux I__5014 (
            .O(N__26026),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_11 ));
    InMux I__5013 (
            .O(N__26023),
            .I(N__26017));
    InMux I__5012 (
            .O(N__26022),
            .I(N__26017));
    LocalMux I__5011 (
            .O(N__26017),
            .I(N__26014));
    Span4Mux_h I__5010 (
            .O(N__26014),
            .I(N__26011));
    Odrv4 I__5009 (
            .O(N__26011),
            .I(\b2v_inst11.dutycycle_RNI9R6T4Z0Z_12 ));
    CascadeMux I__5008 (
            .O(N__26008),
            .I(N__26005));
    InMux I__5007 (
            .O(N__26005),
            .I(N__25999));
    InMux I__5006 (
            .O(N__26004),
            .I(N__25999));
    LocalMux I__5005 (
            .O(N__25999),
            .I(N__25996));
    Odrv12 I__5004 (
            .O(N__25996),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5 ));
    CascadeMux I__5003 (
            .O(N__25993),
            .I(N__25990));
    InMux I__5002 (
            .O(N__25990),
            .I(N__25984));
    InMux I__5001 (
            .O(N__25989),
            .I(N__25984));
    LocalMux I__5000 (
            .O(N__25984),
            .I(\b2v_inst11.dutycycleZ1Z_12 ));
    SRMux I__4999 (
            .O(N__25981),
            .I(N__25977));
    SRMux I__4998 (
            .O(N__25980),
            .I(N__25973));
    LocalMux I__4997 (
            .O(N__25977),
            .I(N__25969));
    SRMux I__4996 (
            .O(N__25976),
            .I(N__25966));
    LocalMux I__4995 (
            .O(N__25973),
            .I(N__25963));
    SRMux I__4994 (
            .O(N__25972),
            .I(N__25960));
    Span4Mux_h I__4993 (
            .O(N__25969),
            .I(N__25955));
    LocalMux I__4992 (
            .O(N__25966),
            .I(N__25955));
    Span4Mux_h I__4991 (
            .O(N__25963),
            .I(N__25952));
    LocalMux I__4990 (
            .O(N__25960),
            .I(N__25949));
    Span4Mux_v I__4989 (
            .O(N__25955),
            .I(N__25938));
    Span4Mux_h I__4988 (
            .O(N__25952),
            .I(N__25938));
    Span4Mux_h I__4987 (
            .O(N__25949),
            .I(N__25938));
    SRMux I__4986 (
            .O(N__25948),
            .I(N__25934));
    SRMux I__4985 (
            .O(N__25947),
            .I(N__25931));
    SRMux I__4984 (
            .O(N__25946),
            .I(N__25928));
    SRMux I__4983 (
            .O(N__25945),
            .I(N__25925));
    Span4Mux_v I__4982 (
            .O(N__25938),
            .I(N__25922));
    SRMux I__4981 (
            .O(N__25937),
            .I(N__25919));
    LocalMux I__4980 (
            .O(N__25934),
            .I(N__25916));
    LocalMux I__4979 (
            .O(N__25931),
            .I(N__25909));
    LocalMux I__4978 (
            .O(N__25928),
            .I(N__25909));
    LocalMux I__4977 (
            .O(N__25925),
            .I(N__25909));
    IoSpan4Mux I__4976 (
            .O(N__25922),
            .I(N__25904));
    LocalMux I__4975 (
            .O(N__25919),
            .I(N__25904));
    Span4Mux_h I__4974 (
            .O(N__25916),
            .I(N__25901));
    Span4Mux_v I__4973 (
            .O(N__25909),
            .I(N__25898));
    Span4Mux_s3_v I__4972 (
            .O(N__25904),
            .I(N__25894));
    Span4Mux_h I__4971 (
            .O(N__25901),
            .I(N__25891));
    Sp12to4 I__4970 (
            .O(N__25898),
            .I(N__25888));
    SRMux I__4969 (
            .O(N__25897),
            .I(N__25885));
    Span4Mux_h I__4968 (
            .O(N__25894),
            .I(N__25882));
    Odrv4 I__4967 (
            .O(N__25891),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv12 I__4966 (
            .O(N__25888),
            .I(\b2v_inst11.N_224_iZ0 ));
    LocalMux I__4965 (
            .O(N__25885),
            .I(\b2v_inst11.N_224_iZ0 ));
    Odrv4 I__4964 (
            .O(N__25882),
            .I(\b2v_inst11.N_224_iZ0 ));
    InMux I__4963 (
            .O(N__25873),
            .I(N__25867));
    InMux I__4962 (
            .O(N__25872),
            .I(N__25867));
    LocalMux I__4961 (
            .O(N__25867),
            .I(\b2v_inst11.dutycycleZ0Z_15 ));
    InMux I__4960 (
            .O(N__25864),
            .I(N__25854));
    InMux I__4959 (
            .O(N__25863),
            .I(N__25844));
    InMux I__4958 (
            .O(N__25862),
            .I(N__25844));
    InMux I__4957 (
            .O(N__25861),
            .I(N__25844));
    InMux I__4956 (
            .O(N__25860),
            .I(N__25844));
    InMux I__4955 (
            .O(N__25859),
            .I(N__25841));
    InMux I__4954 (
            .O(N__25858),
            .I(N__25831));
    CascadeMux I__4953 (
            .O(N__25857),
            .I(N__25827));
    LocalMux I__4952 (
            .O(N__25854),
            .I(N__25820));
    CascadeMux I__4951 (
            .O(N__25853),
            .I(N__25812));
    LocalMux I__4950 (
            .O(N__25844),
            .I(N__25808));
    LocalMux I__4949 (
            .O(N__25841),
            .I(N__25805));
    InMux I__4948 (
            .O(N__25840),
            .I(N__25802));
    InMux I__4947 (
            .O(N__25839),
            .I(N__25789));
    InMux I__4946 (
            .O(N__25838),
            .I(N__25789));
    InMux I__4945 (
            .O(N__25837),
            .I(N__25789));
    InMux I__4944 (
            .O(N__25836),
            .I(N__25789));
    InMux I__4943 (
            .O(N__25835),
            .I(N__25789));
    InMux I__4942 (
            .O(N__25834),
            .I(N__25789));
    LocalMux I__4941 (
            .O(N__25831),
            .I(N__25786));
    InMux I__4940 (
            .O(N__25830),
            .I(N__25777));
    InMux I__4939 (
            .O(N__25827),
            .I(N__25777));
    InMux I__4938 (
            .O(N__25826),
            .I(N__25777));
    InMux I__4937 (
            .O(N__25825),
            .I(N__25777));
    InMux I__4936 (
            .O(N__25824),
            .I(N__25772));
    InMux I__4935 (
            .O(N__25823),
            .I(N__25772));
    Span4Mux_v I__4934 (
            .O(N__25820),
            .I(N__25769));
    InMux I__4933 (
            .O(N__25819),
            .I(N__25758));
    InMux I__4932 (
            .O(N__25818),
            .I(N__25758));
    InMux I__4931 (
            .O(N__25817),
            .I(N__25758));
    InMux I__4930 (
            .O(N__25816),
            .I(N__25758));
    InMux I__4929 (
            .O(N__25815),
            .I(N__25758));
    InMux I__4928 (
            .O(N__25812),
            .I(N__25753));
    InMux I__4927 (
            .O(N__25811),
            .I(N__25753));
    Span4Mux_h I__4926 (
            .O(N__25808),
            .I(N__25746));
    Span4Mux_h I__4925 (
            .O(N__25805),
            .I(N__25746));
    LocalMux I__4924 (
            .O(N__25802),
            .I(N__25746));
    LocalMux I__4923 (
            .O(N__25789),
            .I(N__25739));
    Span12Mux_s6_v I__4922 (
            .O(N__25786),
            .I(N__25739));
    LocalMux I__4921 (
            .O(N__25777),
            .I(N__25739));
    LocalMux I__4920 (
            .O(N__25772),
            .I(N__25736));
    Odrv4 I__4919 (
            .O(N__25769),
            .I(func_state_RNIVS8U1_3_1));
    LocalMux I__4918 (
            .O(N__25758),
            .I(func_state_RNIVS8U1_3_1));
    LocalMux I__4917 (
            .O(N__25753),
            .I(func_state_RNIVS8U1_3_1));
    Odrv4 I__4916 (
            .O(N__25746),
            .I(func_state_RNIVS8U1_3_1));
    Odrv12 I__4915 (
            .O(N__25739),
            .I(func_state_RNIVS8U1_3_1));
    Odrv4 I__4914 (
            .O(N__25736),
            .I(func_state_RNIVS8U1_3_1));
    CascadeMux I__4913 (
            .O(N__25723),
            .I(N__25720));
    InMux I__4912 (
            .O(N__25720),
            .I(N__25714));
    InMux I__4911 (
            .O(N__25719),
            .I(N__25714));
    LocalMux I__4910 (
            .O(N__25714),
            .I(N__25711));
    Span4Mux_h I__4909 (
            .O(N__25711),
            .I(N__25708));
    Odrv4 I__4908 (
            .O(N__25708),
            .I(\b2v_inst11.dutycycle_en_12 ));
    InMux I__4907 (
            .O(N__25705),
            .I(N__25699));
    InMux I__4906 (
            .O(N__25704),
            .I(N__25699));
    LocalMux I__4905 (
            .O(N__25699),
            .I(N__25696));
    Odrv4 I__4904 (
            .O(N__25696),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ));
    InMux I__4903 (
            .O(N__25693),
            .I(N__25690));
    LocalMux I__4902 (
            .O(N__25690),
            .I(N__25687));
    Span4Mux_v I__4901 (
            .O(N__25687),
            .I(N__25684));
    Odrv4 I__4900 (
            .O(N__25684),
            .I(\b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_3_1 ));
    CascadeMux I__4899 (
            .O(N__25681),
            .I(\b2v_inst11.un1_dutycycle_53_50_1_i_i_1_cascade_ ));
    CascadeMux I__4898 (
            .O(N__25678),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ));
    InMux I__4897 (
            .O(N__25675),
            .I(N__25672));
    LocalMux I__4896 (
            .O(N__25672),
            .I(\b2v_inst11.mult1_un110_sum_i ));
    InMux I__4895 (
            .O(N__25669),
            .I(N__25666));
    LocalMux I__4894 (
            .O(N__25666),
            .I(\b2v_inst5.un12_clk_100khz_13 ));
    InMux I__4893 (
            .O(N__25663),
            .I(N__25660));
    LocalMux I__4892 (
            .O(N__25660),
            .I(\b2v_inst11.un1_dutycycle_53_axb_11 ));
    CascadeMux I__4891 (
            .O(N__25657),
            .I(\b2v_inst11.i7_mux_cascade_ ));
    CascadeMux I__4890 (
            .O(N__25654),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_11_cascade_ ));
    InMux I__4889 (
            .O(N__25651),
            .I(N__25648));
    LocalMux I__4888 (
            .O(N__25648),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_9 ));
    CascadeMux I__4887 (
            .O(N__25645),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_8_cascade_ ));
    InMux I__4886 (
            .O(N__25642),
            .I(N__25639));
    LocalMux I__4885 (
            .O(N__25639),
            .I(\b2v_inst11.mult1_un117_sum_cry_4_s ));
    InMux I__4884 (
            .O(N__25636),
            .I(\b2v_inst11.mult1_un117_sum_cry_3 ));
    CascadeMux I__4883 (
            .O(N__25633),
            .I(N__25630));
    InMux I__4882 (
            .O(N__25630),
            .I(N__25627));
    LocalMux I__4881 (
            .O(N__25627),
            .I(\b2v_inst11.mult1_un117_sum_cry_5_s ));
    InMux I__4880 (
            .O(N__25624),
            .I(\b2v_inst11.mult1_un117_sum_cry_4 ));
    InMux I__4879 (
            .O(N__25621),
            .I(N__25618));
    LocalMux I__4878 (
            .O(N__25618),
            .I(\b2v_inst11.mult1_un117_sum_cry_6_s ));
    InMux I__4877 (
            .O(N__25615),
            .I(\b2v_inst11.mult1_un117_sum_cry_5 ));
    CascadeMux I__4876 (
            .O(N__25612),
            .I(N__25609));
    InMux I__4875 (
            .O(N__25609),
            .I(N__25606));
    LocalMux I__4874 (
            .O(N__25606),
            .I(\b2v_inst11.mult1_un124_sum_axb_8 ));
    InMux I__4873 (
            .O(N__25603),
            .I(\b2v_inst11.mult1_un117_sum_cry_6 ));
    InMux I__4872 (
            .O(N__25600),
            .I(\b2v_inst11.mult1_un117_sum_cry_7 ));
    CascadeMux I__4871 (
            .O(N__25597),
            .I(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ));
    CascadeMux I__4870 (
            .O(N__25594),
            .I(N__25590));
    CascadeMux I__4869 (
            .O(N__25593),
            .I(N__25586));
    InMux I__4868 (
            .O(N__25590),
            .I(N__25579));
    InMux I__4867 (
            .O(N__25589),
            .I(N__25579));
    InMux I__4866 (
            .O(N__25586),
            .I(N__25579));
    LocalMux I__4865 (
            .O(N__25579),
            .I(\b2v_inst11.mult1_un117_sum_i_0_8 ));
    InMux I__4864 (
            .O(N__25576),
            .I(N__25573));
    LocalMux I__4863 (
            .O(N__25573),
            .I(N__25570));
    Span4Mux_h I__4862 (
            .O(N__25570),
            .I(N__25566));
    InMux I__4861 (
            .O(N__25569),
            .I(N__25563));
    Span4Mux_v I__4860 (
            .O(N__25566),
            .I(N__25560));
    LocalMux I__4859 (
            .O(N__25563),
            .I(\b2v_inst5.curr_stateZ0Z_1 ));
    Odrv4 I__4858 (
            .O(N__25560),
            .I(\b2v_inst5.curr_stateZ0Z_1 ));
    CascadeMux I__4857 (
            .O(N__25555),
            .I(N__25552));
    InMux I__4856 (
            .O(N__25552),
            .I(N__25549));
    LocalMux I__4855 (
            .O(N__25549),
            .I(N__25544));
    InMux I__4854 (
            .O(N__25548),
            .I(N__25539));
    InMux I__4853 (
            .O(N__25547),
            .I(N__25539));
    Span4Mux_v I__4852 (
            .O(N__25544),
            .I(N__25534));
    LocalMux I__4851 (
            .O(N__25539),
            .I(N__25534));
    Span4Mux_v I__4850 (
            .O(N__25534),
            .I(N__25531));
    Odrv4 I__4849 (
            .O(N__25531),
            .I(N_413));
    InMux I__4848 (
            .O(N__25528),
            .I(N__25525));
    LocalMux I__4847 (
            .O(N__25525),
            .I(\b2v_inst11.mult1_un138_sum_axb_8 ));
    InMux I__4846 (
            .O(N__25522),
            .I(\b2v_inst11.mult1_un138_sum_cry_7 ));
    CascadeMux I__4845 (
            .O(N__25519),
            .I(N__25514));
    CascadeMux I__4844 (
            .O(N__25518),
            .I(N__25511));
    CascadeMux I__4843 (
            .O(N__25517),
            .I(N__25508));
    InMux I__4842 (
            .O(N__25514),
            .I(N__25505));
    InMux I__4841 (
            .O(N__25511),
            .I(N__25500));
    InMux I__4840 (
            .O(N__25508),
            .I(N__25500));
    LocalMux I__4839 (
            .O(N__25505),
            .I(\b2v_inst11.mult1_un131_sum_i_0_8 ));
    LocalMux I__4838 (
            .O(N__25500),
            .I(\b2v_inst11.mult1_un131_sum_i_0_8 ));
    InMux I__4837 (
            .O(N__25495),
            .I(N__25492));
    LocalMux I__4836 (
            .O(N__25492),
            .I(\b2v_inst11.mult1_un117_sum_i ));
    InMux I__4835 (
            .O(N__25489),
            .I(N__25486));
    LocalMux I__4834 (
            .O(N__25486),
            .I(\b2v_inst11.mult1_un131_sum_i ));
    CascadeMux I__4833 (
            .O(N__25483),
            .I(N__25479));
    CascadeMux I__4832 (
            .O(N__25482),
            .I(N__25476));
    InMux I__4831 (
            .O(N__25479),
            .I(N__25470));
    InMux I__4830 (
            .O(N__25476),
            .I(N__25465));
    InMux I__4829 (
            .O(N__25475),
            .I(N__25465));
    InMux I__4828 (
            .O(N__25474),
            .I(N__25462));
    InMux I__4827 (
            .O(N__25473),
            .I(N__25459));
    LocalMux I__4826 (
            .O(N__25470),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__4825 (
            .O(N__25465),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__4824 (
            .O(N__25462),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    LocalMux I__4823 (
            .O(N__25459),
            .I(\b2v_inst11.mult1_un131_sum_s_8 ));
    InMux I__4822 (
            .O(N__25450),
            .I(N__25447));
    LocalMux I__4821 (
            .O(N__25447),
            .I(\b2v_inst11.mult1_un124_sum_i ));
    InMux I__4820 (
            .O(N__25444),
            .I(N__25441));
    LocalMux I__4819 (
            .O(N__25441),
            .I(N__25438));
    Odrv4 I__4818 (
            .O(N__25438),
            .I(\b2v_inst11.mult1_un145_sum_i ));
    CascadeMux I__4817 (
            .O(N__25435),
            .I(N__25432));
    InMux I__4816 (
            .O(N__25432),
            .I(N__25429));
    LocalMux I__4815 (
            .O(N__25429),
            .I(\b2v_inst11.mult1_un117_sum_cry_3_s ));
    InMux I__4814 (
            .O(N__25426),
            .I(\b2v_inst11.mult1_un117_sum_cry_2 ));
    InMux I__4813 (
            .O(N__25423),
            .I(N__25420));
    LocalMux I__4812 (
            .O(N__25420),
            .I(N__25417));
    Odrv4 I__4811 (
            .O(N__25417),
            .I(\b2v_inst5.count_1_12 ));
    InMux I__4810 (
            .O(N__25414),
            .I(N__25411));
    LocalMux I__4809 (
            .O(N__25411),
            .I(\b2v_inst5.count_1_14 ));
    InMux I__4808 (
            .O(N__25408),
            .I(\b2v_inst11.mult1_un138_sum_cry_2 ));
    InMux I__4807 (
            .O(N__25405),
            .I(N__25402));
    LocalMux I__4806 (
            .O(N__25402),
            .I(\b2v_inst11.mult1_un131_sum_cry_3_s ));
    InMux I__4805 (
            .O(N__25399),
            .I(\b2v_inst11.mult1_un138_sum_cry_3 ));
    InMux I__4804 (
            .O(N__25396),
            .I(N__25393));
    LocalMux I__4803 (
            .O(N__25393),
            .I(\b2v_inst11.mult1_un131_sum_cry_4_s ));
    InMux I__4802 (
            .O(N__25390),
            .I(\b2v_inst11.mult1_un138_sum_cry_4 ));
    InMux I__4801 (
            .O(N__25387),
            .I(N__25384));
    LocalMux I__4800 (
            .O(N__25384),
            .I(\b2v_inst11.mult1_un131_sum_cry_5_s ));
    InMux I__4799 (
            .O(N__25381),
            .I(\b2v_inst11.mult1_un138_sum_cry_5 ));
    InMux I__4798 (
            .O(N__25378),
            .I(N__25375));
    LocalMux I__4797 (
            .O(N__25375),
            .I(\b2v_inst11.mult1_un131_sum_cry_6_s ));
    InMux I__4796 (
            .O(N__25372),
            .I(\b2v_inst11.mult1_un138_sum_cry_6 ));
    CascadeMux I__4795 (
            .O(N__25369),
            .I(N__25366));
    InMux I__4794 (
            .O(N__25366),
            .I(N__25357));
    InMux I__4793 (
            .O(N__25365),
            .I(N__25357));
    InMux I__4792 (
            .O(N__25364),
            .I(N__25357));
    LocalMux I__4791 (
            .O(N__25357),
            .I(\b2v_inst36.N_2939_i ));
    CascadeMux I__4790 (
            .O(N__25354),
            .I(N__25348));
    CascadeMux I__4789 (
            .O(N__25353),
            .I(N__25344));
    CascadeMux I__4788 (
            .O(N__25352),
            .I(N__25341));
    CascadeMux I__4787 (
            .O(N__25351),
            .I(N__25337));
    InMux I__4786 (
            .O(N__25348),
            .I(N__25325));
    InMux I__4785 (
            .O(N__25347),
            .I(N__25325));
    InMux I__4784 (
            .O(N__25344),
            .I(N__25325));
    InMux I__4783 (
            .O(N__25341),
            .I(N__25325));
    InMux I__4782 (
            .O(N__25340),
            .I(N__25325));
    InMux I__4781 (
            .O(N__25337),
            .I(N__25320));
    InMux I__4780 (
            .O(N__25336),
            .I(N__25320));
    LocalMux I__4779 (
            .O(N__25325),
            .I(N__25317));
    LocalMux I__4778 (
            .O(N__25320),
            .I(N__25314));
    Span4Mux_h I__4777 (
            .O(N__25317),
            .I(N__25311));
    Span4Mux_v I__4776 (
            .O(N__25314),
            .I(N__25308));
    Sp12to4 I__4775 (
            .O(N__25311),
            .I(N__25305));
    Span4Mux_v I__4774 (
            .O(N__25308),
            .I(N__25302));
    Span12Mux_v I__4773 (
            .O(N__25305),
            .I(N__25299));
    Span4Mux_v I__4772 (
            .O(N__25302),
            .I(N__25296));
    Odrv12 I__4771 (
            .O(N__25299),
            .I(V33DSW_OK_c));
    Odrv4 I__4770 (
            .O(N__25296),
            .I(V33DSW_OK_c));
    InMux I__4769 (
            .O(N__25291),
            .I(N__25280));
    InMux I__4768 (
            .O(N__25290),
            .I(N__25280));
    InMux I__4767 (
            .O(N__25289),
            .I(N__25269));
    InMux I__4766 (
            .O(N__25288),
            .I(N__25269));
    InMux I__4765 (
            .O(N__25287),
            .I(N__25269));
    InMux I__4764 (
            .O(N__25286),
            .I(N__25269));
    InMux I__4763 (
            .O(N__25285),
            .I(N__25269));
    LocalMux I__4762 (
            .O(N__25280),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    LocalMux I__4761 (
            .O(N__25269),
            .I(\b2v_inst36.curr_stateZ0Z_1 ));
    CascadeMux I__4760 (
            .O(N__25264),
            .I(\b2v_inst36.count_rst_7_cascade_ ));
    CascadeMux I__4759 (
            .O(N__25261),
            .I(\b2v_inst36.N_2942_i_cascade_ ));
    InMux I__4758 (
            .O(N__25258),
            .I(N__25254));
    InMux I__4757 (
            .O(N__25257),
            .I(N__25251));
    LocalMux I__4756 (
            .O(N__25254),
            .I(N__25246));
    LocalMux I__4755 (
            .O(N__25251),
            .I(N__25246));
    Span4Mux_h I__4754 (
            .O(N__25246),
            .I(N__25243));
    Odrv4 I__4753 (
            .O(N__25243),
            .I(\b2v_inst200.countZ0Z_9 ));
    InMux I__4752 (
            .O(N__25240),
            .I(N__25234));
    InMux I__4751 (
            .O(N__25239),
            .I(N__25234));
    LocalMux I__4750 (
            .O(N__25234),
            .I(N__25231));
    Span4Mux_h I__4749 (
            .O(N__25231),
            .I(N__25228));
    Odrv4 I__4748 (
            .O(N__25228),
            .I(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ));
    InMux I__4747 (
            .O(N__25225),
            .I(N__25222));
    LocalMux I__4746 (
            .O(N__25222),
            .I(\b2v_inst200.count_3_9 ));
    InMux I__4745 (
            .O(N__25219),
            .I(N__25199));
    InMux I__4744 (
            .O(N__25218),
            .I(N__25192));
    InMux I__4743 (
            .O(N__25217),
            .I(N__25192));
    InMux I__4742 (
            .O(N__25216),
            .I(N__25192));
    InMux I__4741 (
            .O(N__25215),
            .I(N__25185));
    InMux I__4740 (
            .O(N__25214),
            .I(N__25185));
    InMux I__4739 (
            .O(N__25213),
            .I(N__25185));
    InMux I__4738 (
            .O(N__25212),
            .I(N__25178));
    InMux I__4737 (
            .O(N__25211),
            .I(N__25178));
    InMux I__4736 (
            .O(N__25210),
            .I(N__25178));
    InMux I__4735 (
            .O(N__25209),
            .I(N__25169));
    InMux I__4734 (
            .O(N__25208),
            .I(N__25169));
    InMux I__4733 (
            .O(N__25207),
            .I(N__25169));
    InMux I__4732 (
            .O(N__25206),
            .I(N__25169));
    InMux I__4731 (
            .O(N__25205),
            .I(N__25162));
    InMux I__4730 (
            .O(N__25204),
            .I(N__25162));
    InMux I__4729 (
            .O(N__25203),
            .I(N__25162));
    InMux I__4728 (
            .O(N__25202),
            .I(N__25159));
    LocalMux I__4727 (
            .O(N__25199),
            .I(N__25150));
    LocalMux I__4726 (
            .O(N__25192),
            .I(N__25147));
    LocalMux I__4725 (
            .O(N__25185),
            .I(N__25144));
    LocalMux I__4724 (
            .O(N__25178),
            .I(N__25141));
    LocalMux I__4723 (
            .O(N__25169),
            .I(N__25138));
    LocalMux I__4722 (
            .O(N__25162),
            .I(N__25135));
    LocalMux I__4721 (
            .O(N__25159),
            .I(N__25132));
    CEMux I__4720 (
            .O(N__25158),
            .I(N__25105));
    CEMux I__4719 (
            .O(N__25157),
            .I(N__25105));
    CEMux I__4718 (
            .O(N__25156),
            .I(N__25105));
    CEMux I__4717 (
            .O(N__25155),
            .I(N__25105));
    CEMux I__4716 (
            .O(N__25154),
            .I(N__25105));
    CEMux I__4715 (
            .O(N__25153),
            .I(N__25105));
    Glb2LocalMux I__4714 (
            .O(N__25150),
            .I(N__25105));
    Glb2LocalMux I__4713 (
            .O(N__25147),
            .I(N__25105));
    Glb2LocalMux I__4712 (
            .O(N__25144),
            .I(N__25105));
    Glb2LocalMux I__4711 (
            .O(N__25141),
            .I(N__25105));
    Glb2LocalMux I__4710 (
            .O(N__25138),
            .I(N__25105));
    Glb2LocalMux I__4709 (
            .O(N__25135),
            .I(N__25105));
    Glb2LocalMux I__4708 (
            .O(N__25132),
            .I(N__25105));
    GlobalMux I__4707 (
            .O(N__25105),
            .I(N__25102));
    gio2CtrlBuf I__4706 (
            .O(N__25102),
            .I(\b2v_inst200.count_en_g ));
    InMux I__4705 (
            .O(N__25099),
            .I(N__25096));
    LocalMux I__4704 (
            .O(N__25096),
            .I(N__25093));
    Odrv4 I__4703 (
            .O(N__25093),
            .I(\b2v_inst36.count_2_14 ));
    InMux I__4702 (
            .O(N__25090),
            .I(N__25087));
    LocalMux I__4701 (
            .O(N__25087),
            .I(\b2v_inst5.count_1_11 ));
    CascadeMux I__4700 (
            .O(N__25084),
            .I(\b2v_inst36.count_rst_3_cascade_ ));
    CascadeMux I__4699 (
            .O(N__25081),
            .I(\b2v_inst36.countZ0Z_11_cascade_ ));
    InMux I__4698 (
            .O(N__25078),
            .I(N__25075));
    LocalMux I__4697 (
            .O(N__25075),
            .I(\b2v_inst36.count_2_11 ));
    CascadeMux I__4696 (
            .O(N__25072),
            .I(\b2v_inst36.count_rst_12_cascade_ ));
    CascadeMux I__4695 (
            .O(N__25069),
            .I(\b2v_inst36.countZ0Z_2_cascade_ ));
    InMux I__4694 (
            .O(N__25066),
            .I(N__25063));
    LocalMux I__4693 (
            .O(N__25063),
            .I(\b2v_inst36.count_2_2 ));
    InMux I__4692 (
            .O(N__25060),
            .I(N__25057));
    LocalMux I__4691 (
            .O(N__25057),
            .I(\b2v_inst36.curr_state_7_1 ));
    CascadeMux I__4690 (
            .O(N__25054),
            .I(\b2v_inst36.curr_stateZ0Z_1_cascade_ ));
    InMux I__4689 (
            .O(N__25051),
            .I(N__25048));
    LocalMux I__4688 (
            .O(N__25048),
            .I(\b2v_inst36.curr_state_0_1 ));
    CascadeMux I__4687 (
            .O(N__25045),
            .I(\b2v_inst36.countZ0Z_1_cascade_ ));
    InMux I__4686 (
            .O(N__25042),
            .I(N__25039));
    LocalMux I__4685 (
            .O(N__25039),
            .I(N__25036));
    Odrv4 I__4684 (
            .O(N__25036),
            .I(\b2v_inst36.un12_clk_100khz_9 ));
    CascadeMux I__4683 (
            .O(N__25033),
            .I(\b2v_inst36.un12_clk_100khz_10_cascade_ ));
    InMux I__4682 (
            .O(N__25030),
            .I(N__25027));
    LocalMux I__4681 (
            .O(N__25027),
            .I(\b2v_inst36.count_2_0 ));
    CascadeMux I__4680 (
            .O(N__25024),
            .I(\b2v_inst36.countZ0Z_0_cascade_ ));
    InMux I__4679 (
            .O(N__25021),
            .I(N__25018));
    LocalMux I__4678 (
            .O(N__25018),
            .I(\b2v_inst36.count_rst_13 ));
    CascadeMux I__4677 (
            .O(N__25015),
            .I(\b2v_inst36.count_rst_13_cascade_ ));
    CascadeMux I__4676 (
            .O(N__25012),
            .I(\b2v_inst36.un2_count_1_axb_1_cascade_ ));
    InMux I__4675 (
            .O(N__25009),
            .I(N__25003));
    InMux I__4674 (
            .O(N__25008),
            .I(N__25003));
    LocalMux I__4673 (
            .O(N__25003),
            .I(\b2v_inst36.count_2_1 ));
    InMux I__4672 (
            .O(N__25000),
            .I(N__24997));
    LocalMux I__4671 (
            .O(N__24997),
            .I(\b2v_inst36.un12_clk_100khz_8 ));
    InMux I__4670 (
            .O(N__24994),
            .I(N__24991));
    LocalMux I__4669 (
            .O(N__24991),
            .I(\b2v_inst36.count_rst_14 ));
    CascadeMux I__4668 (
            .O(N__24988),
            .I(N__24985));
    InMux I__4667 (
            .O(N__24985),
            .I(N__24979));
    InMux I__4666 (
            .O(N__24984),
            .I(N__24979));
    LocalMux I__4665 (
            .O(N__24979),
            .I(N__24976));
    Odrv4 I__4664 (
            .O(N__24976),
            .I(\b2v_inst11.count_1_6 ));
    InMux I__4663 (
            .O(N__24973),
            .I(N__24970));
    LocalMux I__4662 (
            .O(N__24970),
            .I(\b2v_inst11.count_0_6 ));
    CascadeMux I__4661 (
            .O(N__24967),
            .I(N__24964));
    InMux I__4660 (
            .O(N__24964),
            .I(N__24958));
    InMux I__4659 (
            .O(N__24963),
            .I(N__24958));
    LocalMux I__4658 (
            .O(N__24958),
            .I(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ));
    InMux I__4657 (
            .O(N__24955),
            .I(N__24952));
    LocalMux I__4656 (
            .O(N__24952),
            .I(\b2v_inst11.count_0_15 ));
    CascadeMux I__4655 (
            .O(N__24949),
            .I(\b2v_inst11.pwm_out_en_cascade_ ));
    IoInMux I__4654 (
            .O(N__24946),
            .I(N__24943));
    LocalMux I__4653 (
            .O(N__24943),
            .I(PWRBTN_LED_c));
    InMux I__4652 (
            .O(N__24940),
            .I(N__24937));
    LocalMux I__4651 (
            .O(N__24937),
            .I(\b2v_inst11.pwm_out_1_sqmuxa_0 ));
    InMux I__4650 (
            .O(N__24934),
            .I(N__24928));
    CascadeMux I__4649 (
            .O(N__24933),
            .I(N__24925));
    CascadeMux I__4648 (
            .O(N__24932),
            .I(N__24921));
    InMux I__4647 (
            .O(N__24931),
            .I(N__24917));
    LocalMux I__4646 (
            .O(N__24928),
            .I(N__24914));
    InMux I__4645 (
            .O(N__24925),
            .I(N__24911));
    InMux I__4644 (
            .O(N__24924),
            .I(N__24908));
    InMux I__4643 (
            .O(N__24921),
            .I(N__24905));
    InMux I__4642 (
            .O(N__24920),
            .I(N__24902));
    LocalMux I__4641 (
            .O(N__24917),
            .I(N__24895));
    Span4Mux_h I__4640 (
            .O(N__24914),
            .I(N__24895));
    LocalMux I__4639 (
            .O(N__24911),
            .I(N__24890));
    LocalMux I__4638 (
            .O(N__24908),
            .I(N__24890));
    LocalMux I__4637 (
            .O(N__24905),
            .I(N__24885));
    LocalMux I__4636 (
            .O(N__24902),
            .I(N__24885));
    InMux I__4635 (
            .O(N__24901),
            .I(N__24880));
    InMux I__4634 (
            .O(N__24900),
            .I(N__24880));
    Span4Mux_v I__4633 (
            .O(N__24895),
            .I(N__24875));
    Span4Mux_h I__4632 (
            .O(N__24890),
            .I(N__24875));
    Span4Mux_h I__4631 (
            .O(N__24885),
            .I(N__24872));
    LocalMux I__4630 (
            .O(N__24880),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    Odrv4 I__4629 (
            .O(N__24875),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    Odrv4 I__4628 (
            .O(N__24872),
            .I(SYNTHESIZED_WIRE_1keep_3_rep1));
    CascadeMux I__4627 (
            .O(N__24865),
            .I(N__24861));
    CascadeMux I__4626 (
            .O(N__24864),
            .I(N__24858));
    InMux I__4625 (
            .O(N__24861),
            .I(N__24850));
    InMux I__4624 (
            .O(N__24858),
            .I(N__24850));
    InMux I__4623 (
            .O(N__24857),
            .I(N__24850));
    LocalMux I__4622 (
            .O(N__24850),
            .I(N__24846));
    InMux I__4621 (
            .O(N__24849),
            .I(N__24842));
    Span4Mux_v I__4620 (
            .O(N__24846),
            .I(N__24832));
    InMux I__4619 (
            .O(N__24845),
            .I(N__24829));
    LocalMux I__4618 (
            .O(N__24842),
            .I(N__24826));
    InMux I__4617 (
            .O(N__24841),
            .I(N__24815));
    InMux I__4616 (
            .O(N__24840),
            .I(N__24815));
    InMux I__4615 (
            .O(N__24839),
            .I(N__24815));
    InMux I__4614 (
            .O(N__24838),
            .I(N__24815));
    InMux I__4613 (
            .O(N__24837),
            .I(N__24815));
    InMux I__4612 (
            .O(N__24836),
            .I(N__24810));
    InMux I__4611 (
            .O(N__24835),
            .I(N__24810));
    Span4Mux_v I__4610 (
            .O(N__24832),
            .I(N__24805));
    LocalMux I__4609 (
            .O(N__24829),
            .I(N__24805));
    Span4Mux_v I__4608 (
            .O(N__24826),
            .I(N__24802));
    LocalMux I__4607 (
            .O(N__24815),
            .I(N__24797));
    LocalMux I__4606 (
            .O(N__24810),
            .I(N__24797));
    Span4Mux_h I__4605 (
            .O(N__24805),
            .I(N__24794));
    Odrv4 I__4604 (
            .O(N__24802),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv12 I__4603 (
            .O(N__24797),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    Odrv4 I__4602 (
            .O(N__24794),
            .I(b2v_inst20_un4_counter_7_THRU_CO));
    CascadeMux I__4601 (
            .O(N__24787),
            .I(N__24784));
    InMux I__4600 (
            .O(N__24784),
            .I(N__24778));
    InMux I__4599 (
            .O(N__24783),
            .I(N__24778));
    LocalMux I__4598 (
            .O(N__24778),
            .I(\b2v_inst11.count_1_11 ));
    InMux I__4597 (
            .O(N__24775),
            .I(\b2v_inst11.un1_count_cry_10 ));
    InMux I__4596 (
            .O(N__24772),
            .I(\b2v_inst11.un1_count_cry_11 ));
    InMux I__4595 (
            .O(N__24769),
            .I(\b2v_inst11.un1_count_cry_12 ));
    InMux I__4594 (
            .O(N__24766),
            .I(\b2v_inst11.un1_count_cry_13 ));
    InMux I__4593 (
            .O(N__24763),
            .I(\b2v_inst11.un1_count_cry_14 ));
    CascadeMux I__4592 (
            .O(N__24760),
            .I(N__24757));
    InMux I__4591 (
            .O(N__24757),
            .I(N__24751));
    InMux I__4590 (
            .O(N__24756),
            .I(N__24751));
    LocalMux I__4589 (
            .O(N__24751),
            .I(N__24748));
    Odrv4 I__4588 (
            .O(N__24748),
            .I(\b2v_inst11.count_1_5 ));
    InMux I__4587 (
            .O(N__24745),
            .I(N__24742));
    LocalMux I__4586 (
            .O(N__24742),
            .I(\b2v_inst11.count_0_5 ));
    InMux I__4585 (
            .O(N__24739),
            .I(N__24735));
    InMux I__4584 (
            .O(N__24738),
            .I(N__24732));
    LocalMux I__4583 (
            .O(N__24735),
            .I(\b2v_inst11.count_1_14 ));
    LocalMux I__4582 (
            .O(N__24732),
            .I(\b2v_inst11.count_1_14 ));
    InMux I__4581 (
            .O(N__24727),
            .I(N__24724));
    LocalMux I__4580 (
            .O(N__24724),
            .I(\b2v_inst11.count_0_14 ));
    CascadeMux I__4579 (
            .O(N__24721),
            .I(N__24717));
    InMux I__4578 (
            .O(N__24720),
            .I(N__24712));
    InMux I__4577 (
            .O(N__24717),
            .I(N__24712));
    LocalMux I__4576 (
            .O(N__24712),
            .I(N__24709));
    Odrv4 I__4575 (
            .O(N__24709),
            .I(\b2v_inst11.count_1_2 ));
    InMux I__4574 (
            .O(N__24706),
            .I(\b2v_inst11.un1_count_cry_1 ));
    InMux I__4573 (
            .O(N__24703),
            .I(\b2v_inst11.un1_count_cry_2 ));
    InMux I__4572 (
            .O(N__24700),
            .I(\b2v_inst11.un1_count_cry_3 ));
    InMux I__4571 (
            .O(N__24697),
            .I(\b2v_inst11.un1_count_cry_4 ));
    InMux I__4570 (
            .O(N__24694),
            .I(\b2v_inst11.un1_count_cry_5 ));
    InMux I__4569 (
            .O(N__24691),
            .I(N__24685));
    InMux I__4568 (
            .O(N__24690),
            .I(N__24685));
    LocalMux I__4567 (
            .O(N__24685),
            .I(N__24682));
    Odrv4 I__4566 (
            .O(N__24682),
            .I(\b2v_inst11.count_1_7 ));
    InMux I__4565 (
            .O(N__24679),
            .I(\b2v_inst11.un1_count_cry_6 ));
    InMux I__4564 (
            .O(N__24676),
            .I(\b2v_inst11.un1_count_cry_7 ));
    CascadeMux I__4563 (
            .O(N__24673),
            .I(N__24670));
    InMux I__4562 (
            .O(N__24670),
            .I(N__24664));
    InMux I__4561 (
            .O(N__24669),
            .I(N__24664));
    LocalMux I__4560 (
            .O(N__24664),
            .I(\b2v_inst11.count_1_9 ));
    InMux I__4559 (
            .O(N__24661),
            .I(bfn_7_14_0_));
    CascadeMux I__4558 (
            .O(N__24658),
            .I(N__24654));
    InMux I__4557 (
            .O(N__24657),
            .I(N__24649));
    InMux I__4556 (
            .O(N__24654),
            .I(N__24649));
    LocalMux I__4555 (
            .O(N__24649),
            .I(\b2v_inst11.count_1_10 ));
    InMux I__4554 (
            .O(N__24646),
            .I(\b2v_inst11.un1_count_cry_9 ));
    InMux I__4553 (
            .O(N__24643),
            .I(N__24634));
    InMux I__4552 (
            .O(N__24642),
            .I(N__24631));
    InMux I__4551 (
            .O(N__24641),
            .I(N__24626));
    InMux I__4550 (
            .O(N__24640),
            .I(N__24626));
    InMux I__4549 (
            .O(N__24639),
            .I(N__24623));
    InMux I__4548 (
            .O(N__24638),
            .I(N__24619));
    InMux I__4547 (
            .O(N__24637),
            .I(N__24616));
    LocalMux I__4546 (
            .O(N__24634),
            .I(N__24607));
    LocalMux I__4545 (
            .O(N__24631),
            .I(N__24607));
    LocalMux I__4544 (
            .O(N__24626),
            .I(N__24607));
    LocalMux I__4543 (
            .O(N__24623),
            .I(N__24607));
    InMux I__4542 (
            .O(N__24622),
            .I(N__24601));
    LocalMux I__4541 (
            .O(N__24619),
            .I(N__24596));
    LocalMux I__4540 (
            .O(N__24616),
            .I(N__24596));
    Span4Mux_v I__4539 (
            .O(N__24607),
            .I(N__24593));
    InMux I__4538 (
            .O(N__24606),
            .I(N__24588));
    InMux I__4537 (
            .O(N__24605),
            .I(N__24588));
    CascadeMux I__4536 (
            .O(N__24604),
            .I(N__24583));
    LocalMux I__4535 (
            .O(N__24601),
            .I(N__24577));
    Span4Mux_h I__4534 (
            .O(N__24596),
            .I(N__24574));
    Sp12to4 I__4533 (
            .O(N__24593),
            .I(N__24569));
    LocalMux I__4532 (
            .O(N__24588),
            .I(N__24569));
    InMux I__4531 (
            .O(N__24587),
            .I(N__24566));
    InMux I__4530 (
            .O(N__24586),
            .I(N__24563));
    InMux I__4529 (
            .O(N__24583),
            .I(N__24555));
    InMux I__4528 (
            .O(N__24582),
            .I(N__24555));
    InMux I__4527 (
            .O(N__24581),
            .I(N__24555));
    InMux I__4526 (
            .O(N__24580),
            .I(N__24552));
    Sp12to4 I__4525 (
            .O(N__24577),
            .I(N__24549));
    Span4Mux_v I__4524 (
            .O(N__24574),
            .I(N__24546));
    Span12Mux_s4_h I__4523 (
            .O(N__24569),
            .I(N__24539));
    LocalMux I__4522 (
            .O(N__24566),
            .I(N__24539));
    LocalMux I__4521 (
            .O(N__24563),
            .I(N__24539));
    InMux I__4520 (
            .O(N__24562),
            .I(N__24536));
    LocalMux I__4519 (
            .O(N__24555),
            .I(N__24531));
    LocalMux I__4518 (
            .O(N__24552),
            .I(N__24531));
    Odrv12 I__4517 (
            .O(N__24549),
            .I(GPIO_FPGA_SoC_4_c));
    Odrv4 I__4516 (
            .O(N__24546),
            .I(GPIO_FPGA_SoC_4_c));
    Odrv12 I__4515 (
            .O(N__24539),
            .I(GPIO_FPGA_SoC_4_c));
    LocalMux I__4514 (
            .O(N__24536),
            .I(GPIO_FPGA_SoC_4_c));
    Odrv4 I__4513 (
            .O(N__24531),
            .I(GPIO_FPGA_SoC_4_c));
    CascadeMux I__4512 (
            .O(N__24520),
            .I(N__24516));
    CascadeMux I__4511 (
            .O(N__24519),
            .I(N__24507));
    InMux I__4510 (
            .O(N__24516),
            .I(N__24504));
    CascadeMux I__4509 (
            .O(N__24515),
            .I(N__24501));
    InMux I__4508 (
            .O(N__24514),
            .I(N__24497));
    CascadeMux I__4507 (
            .O(N__24513),
            .I(N__24494));
    InMux I__4506 (
            .O(N__24512),
            .I(N__24491));
    InMux I__4505 (
            .O(N__24511),
            .I(N__24488));
    InMux I__4504 (
            .O(N__24510),
            .I(N__24485));
    InMux I__4503 (
            .O(N__24507),
            .I(N__24481));
    LocalMux I__4502 (
            .O(N__24504),
            .I(N__24478));
    InMux I__4501 (
            .O(N__24501),
            .I(N__24473));
    InMux I__4500 (
            .O(N__24500),
            .I(N__24473));
    LocalMux I__4499 (
            .O(N__24497),
            .I(N__24470));
    InMux I__4498 (
            .O(N__24494),
            .I(N__24466));
    LocalMux I__4497 (
            .O(N__24491),
            .I(N__24461));
    LocalMux I__4496 (
            .O(N__24488),
            .I(N__24461));
    LocalMux I__4495 (
            .O(N__24485),
            .I(N__24458));
    InMux I__4494 (
            .O(N__24484),
            .I(N__24455));
    LocalMux I__4493 (
            .O(N__24481),
            .I(N__24452));
    Span4Mux_h I__4492 (
            .O(N__24478),
            .I(N__24449));
    LocalMux I__4491 (
            .O(N__24473),
            .I(N__24446));
    Span4Mux_v I__4490 (
            .O(N__24470),
            .I(N__24443));
    InMux I__4489 (
            .O(N__24469),
            .I(N__24440));
    LocalMux I__4488 (
            .O(N__24466),
            .I(N__24437));
    Span4Mux_v I__4487 (
            .O(N__24461),
            .I(N__24434));
    Span4Mux_s2_v I__4486 (
            .O(N__24458),
            .I(N__24429));
    LocalMux I__4485 (
            .O(N__24455),
            .I(N__24429));
    Span4Mux_v I__4484 (
            .O(N__24452),
            .I(N__24426));
    Span4Mux_v I__4483 (
            .O(N__24449),
            .I(N__24415));
    Span4Mux_s2_h I__4482 (
            .O(N__24446),
            .I(N__24415));
    Span4Mux_h I__4481 (
            .O(N__24443),
            .I(N__24415));
    LocalMux I__4480 (
            .O(N__24440),
            .I(N__24415));
    Span4Mux_h I__4479 (
            .O(N__24437),
            .I(N__24415));
    Span4Mux_h I__4478 (
            .O(N__24434),
            .I(N__24410));
    Span4Mux_v I__4477 (
            .O(N__24429),
            .I(N__24410));
    Span4Mux_s2_h I__4476 (
            .O(N__24426),
            .I(N__24405));
    Span4Mux_v I__4475 (
            .O(N__24415),
            .I(N__24405));
    Odrv4 I__4474 (
            .O(N__24410),
            .I(N_161));
    Odrv4 I__4473 (
            .O(N__24405),
            .I(N_161));
    CascadeMux I__4472 (
            .O(N__24400),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ));
    InMux I__4471 (
            .O(N__24397),
            .I(N__24376));
    InMux I__4470 (
            .O(N__24396),
            .I(N__24376));
    InMux I__4469 (
            .O(N__24395),
            .I(N__24376));
    InMux I__4468 (
            .O(N__24394),
            .I(N__24376));
    InMux I__4467 (
            .O(N__24393),
            .I(N__24376));
    InMux I__4466 (
            .O(N__24392),
            .I(N__24371));
    InMux I__4465 (
            .O(N__24391),
            .I(N__24371));
    InMux I__4464 (
            .O(N__24390),
            .I(N__24367));
    InMux I__4463 (
            .O(N__24389),
            .I(N__24362));
    InMux I__4462 (
            .O(N__24388),
            .I(N__24358));
    InMux I__4461 (
            .O(N__24387),
            .I(N__24355));
    LocalMux I__4460 (
            .O(N__24376),
            .I(N__24350));
    LocalMux I__4459 (
            .O(N__24371),
            .I(N__24350));
    InMux I__4458 (
            .O(N__24370),
            .I(N__24347));
    LocalMux I__4457 (
            .O(N__24367),
            .I(N__24344));
    InMux I__4456 (
            .O(N__24366),
            .I(N__24341));
    InMux I__4455 (
            .O(N__24365),
            .I(N__24338));
    LocalMux I__4454 (
            .O(N__24362),
            .I(N__24335));
    InMux I__4453 (
            .O(N__24361),
            .I(N__24332));
    LocalMux I__4452 (
            .O(N__24358),
            .I(N__24325));
    LocalMux I__4451 (
            .O(N__24355),
            .I(N__24320));
    Span4Mux_h I__4450 (
            .O(N__24350),
            .I(N__24320));
    LocalMux I__4449 (
            .O(N__24347),
            .I(N__24314));
    Span4Mux_v I__4448 (
            .O(N__24344),
            .I(N__24309));
    LocalMux I__4447 (
            .O(N__24341),
            .I(N__24309));
    LocalMux I__4446 (
            .O(N__24338),
            .I(N__24305));
    Span4Mux_v I__4445 (
            .O(N__24335),
            .I(N__24300));
    LocalMux I__4444 (
            .O(N__24332),
            .I(N__24300));
    InMux I__4443 (
            .O(N__24331),
            .I(N__24297));
    InMux I__4442 (
            .O(N__24330),
            .I(N__24290));
    InMux I__4441 (
            .O(N__24329),
            .I(N__24290));
    InMux I__4440 (
            .O(N__24328),
            .I(N__24290));
    Span4Mux_v I__4439 (
            .O(N__24325),
            .I(N__24285));
    Span4Mux_v I__4438 (
            .O(N__24320),
            .I(N__24285));
    InMux I__4437 (
            .O(N__24319),
            .I(N__24278));
    InMux I__4436 (
            .O(N__24318),
            .I(N__24278));
    InMux I__4435 (
            .O(N__24317),
            .I(N__24278));
    Span4Mux_h I__4434 (
            .O(N__24314),
            .I(N__24275));
    Span4Mux_v I__4433 (
            .O(N__24309),
            .I(N__24272));
    InMux I__4432 (
            .O(N__24308),
            .I(N__24269));
    Span4Mux_v I__4431 (
            .O(N__24305),
            .I(N__24266));
    Span4Mux_h I__4430 (
            .O(N__24300),
            .I(N__24259));
    LocalMux I__4429 (
            .O(N__24297),
            .I(N__24259));
    LocalMux I__4428 (
            .O(N__24290),
            .I(N__24259));
    Span4Mux_v I__4427 (
            .O(N__24285),
            .I(N__24254));
    LocalMux I__4426 (
            .O(N__24278),
            .I(N__24254));
    Span4Mux_v I__4425 (
            .O(N__24275),
            .I(N__24251));
    Span4Mux_v I__4424 (
            .O(N__24272),
            .I(N__24246));
    LocalMux I__4423 (
            .O(N__24269),
            .I(N__24246));
    Span4Mux_v I__4422 (
            .O(N__24266),
            .I(N__24241));
    Span4Mux_v I__4421 (
            .O(N__24259),
            .I(N__24241));
    Span4Mux_h I__4420 (
            .O(N__24254),
            .I(N__24238));
    Span4Mux_h I__4419 (
            .O(N__24251),
            .I(N__24233));
    Span4Mux_h I__4418 (
            .O(N__24246),
            .I(N__24233));
    Odrv4 I__4417 (
            .O(N__24241),
            .I(SLP_S3n_c));
    Odrv4 I__4416 (
            .O(N__24238),
            .I(SLP_S3n_c));
    Odrv4 I__4415 (
            .O(N__24233),
            .I(SLP_S3n_c));
    InMux I__4414 (
            .O(N__24226),
            .I(N__24223));
    LocalMux I__4413 (
            .O(N__24223),
            .I(N__24220));
    Odrv4 I__4412 (
            .O(N__24220),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_c_RNIZ0 ));
    CascadeMux I__4411 (
            .O(N__24217),
            .I(N__24214));
    InMux I__4410 (
            .O(N__24214),
            .I(N__24208));
    InMux I__4409 (
            .O(N__24213),
            .I(N__24205));
    InMux I__4408 (
            .O(N__24212),
            .I(N__24202));
    InMux I__4407 (
            .O(N__24211),
            .I(N__24199));
    LocalMux I__4406 (
            .O(N__24208),
            .I(N__24196));
    LocalMux I__4405 (
            .O(N__24205),
            .I(N__24191));
    LocalMux I__4404 (
            .O(N__24202),
            .I(N__24191));
    LocalMux I__4403 (
            .O(N__24199),
            .I(N__24187));
    Span4Mux_h I__4402 (
            .O(N__24196),
            .I(N__24184));
    Span4Mux_v I__4401 (
            .O(N__24191),
            .I(N__24181));
    InMux I__4400 (
            .O(N__24190),
            .I(N__24178));
    Span4Mux_s3_h I__4399 (
            .O(N__24187),
            .I(N__24175));
    Odrv4 I__4398 (
            .O(N__24184),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    Odrv4 I__4397 (
            .O(N__24181),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    LocalMux I__4396 (
            .O(N__24178),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    Odrv4 I__4395 (
            .O(N__24175),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1 ));
    CascadeMux I__4394 (
            .O(N__24166),
            .I(N__24163));
    InMux I__4393 (
            .O(N__24163),
            .I(N__24156));
    InMux I__4392 (
            .O(N__24162),
            .I(N__24156));
    CascadeMux I__4391 (
            .O(N__24161),
            .I(N__24152));
    LocalMux I__4390 (
            .O(N__24156),
            .I(N__24145));
    InMux I__4389 (
            .O(N__24155),
            .I(N__24142));
    InMux I__4388 (
            .O(N__24152),
            .I(N__24133));
    InMux I__4387 (
            .O(N__24151),
            .I(N__24133));
    InMux I__4386 (
            .O(N__24150),
            .I(N__24133));
    InMux I__4385 (
            .O(N__24149),
            .I(N__24133));
    CascadeMux I__4384 (
            .O(N__24148),
            .I(N__24129));
    Span4Mux_s3_h I__4383 (
            .O(N__24145),
            .I(N__24120));
    LocalMux I__4382 (
            .O(N__24142),
            .I(N__24120));
    LocalMux I__4381 (
            .O(N__24133),
            .I(N__24117));
    InMux I__4380 (
            .O(N__24132),
            .I(N__24114));
    InMux I__4379 (
            .O(N__24129),
            .I(N__24108));
    CascadeMux I__4378 (
            .O(N__24128),
            .I(N__24105));
    InMux I__4377 (
            .O(N__24127),
            .I(N__24097));
    InMux I__4376 (
            .O(N__24126),
            .I(N__24094));
    InMux I__4375 (
            .O(N__24125),
            .I(N__24091));
    Span4Mux_h I__4374 (
            .O(N__24120),
            .I(N__24086));
    Span4Mux_s3_h I__4373 (
            .O(N__24117),
            .I(N__24086));
    LocalMux I__4372 (
            .O(N__24114),
            .I(N__24083));
    InMux I__4371 (
            .O(N__24113),
            .I(N__24076));
    InMux I__4370 (
            .O(N__24112),
            .I(N__24076));
    InMux I__4369 (
            .O(N__24111),
            .I(N__24076));
    LocalMux I__4368 (
            .O(N__24108),
            .I(N__24073));
    InMux I__4367 (
            .O(N__24105),
            .I(N__24066));
    InMux I__4366 (
            .O(N__24104),
            .I(N__24066));
    InMux I__4365 (
            .O(N__24103),
            .I(N__24066));
    InMux I__4364 (
            .O(N__24102),
            .I(N__24063));
    CascadeMux I__4363 (
            .O(N__24101),
            .I(N__24060));
    CascadeMux I__4362 (
            .O(N__24100),
            .I(N__24057));
    LocalMux I__4361 (
            .O(N__24097),
            .I(N__24053));
    LocalMux I__4360 (
            .O(N__24094),
            .I(N__24047));
    LocalMux I__4359 (
            .O(N__24091),
            .I(N__24047));
    Span4Mux_v I__4358 (
            .O(N__24086),
            .I(N__24040));
    Span4Mux_s3_h I__4357 (
            .O(N__24083),
            .I(N__24040));
    LocalMux I__4356 (
            .O(N__24076),
            .I(N__24040));
    Span4Mux_s3_h I__4355 (
            .O(N__24073),
            .I(N__24035));
    LocalMux I__4354 (
            .O(N__24066),
            .I(N__24035));
    LocalMux I__4353 (
            .O(N__24063),
            .I(N__24032));
    InMux I__4352 (
            .O(N__24060),
            .I(N__24029));
    InMux I__4351 (
            .O(N__24057),
            .I(N__24026));
    CascadeMux I__4350 (
            .O(N__24056),
            .I(N__24022));
    Span4Mux_s3_h I__4349 (
            .O(N__24053),
            .I(N__24018));
    InMux I__4348 (
            .O(N__24052),
            .I(N__24015));
    Span4Mux_h I__4347 (
            .O(N__24047),
            .I(N__24012));
    Span4Mux_h I__4346 (
            .O(N__24040),
            .I(N__24009));
    Span4Mux_v I__4345 (
            .O(N__24035),
            .I(N__24000));
    Span4Mux_h I__4344 (
            .O(N__24032),
            .I(N__24000));
    LocalMux I__4343 (
            .O(N__24029),
            .I(N__24000));
    LocalMux I__4342 (
            .O(N__24026),
            .I(N__24000));
    InMux I__4341 (
            .O(N__24025),
            .I(N__23995));
    InMux I__4340 (
            .O(N__24022),
            .I(N__23995));
    InMux I__4339 (
            .O(N__24021),
            .I(N__23992));
    Sp12to4 I__4338 (
            .O(N__24018),
            .I(N__23986));
    LocalMux I__4337 (
            .O(N__24015),
            .I(N__23986));
    Span4Mux_v I__4336 (
            .O(N__24012),
            .I(N__23983));
    Span4Mux_v I__4335 (
            .O(N__24009),
            .I(N__23980));
    Span4Mux_v I__4334 (
            .O(N__24000),
            .I(N__23975));
    LocalMux I__4333 (
            .O(N__23995),
            .I(N__23975));
    LocalMux I__4332 (
            .O(N__23992),
            .I(N__23972));
    InMux I__4331 (
            .O(N__23991),
            .I(N__23969));
    Odrv12 I__4330 (
            .O(N__23986),
            .I(SLP_S4n_c));
    Odrv4 I__4329 (
            .O(N__23983),
            .I(SLP_S4n_c));
    Odrv4 I__4328 (
            .O(N__23980),
            .I(SLP_S4n_c));
    Odrv4 I__4327 (
            .O(N__23975),
            .I(SLP_S4n_c));
    Odrv12 I__4326 (
            .O(N__23972),
            .I(SLP_S4n_c));
    LocalMux I__4325 (
            .O(N__23969),
            .I(SLP_S4n_c));
    CascadeMux I__4324 (
            .O(N__23956),
            .I(\b2v_inst11.g1_0_0_cascade_ ));
    InMux I__4323 (
            .O(N__23953),
            .I(N__23950));
    LocalMux I__4322 (
            .O(N__23950),
            .I(\b2v_inst11.N_295 ));
    CascadeMux I__4321 (
            .O(N__23947),
            .I(N__23944));
    InMux I__4320 (
            .O(N__23944),
            .I(N__23941));
    LocalMux I__4319 (
            .O(N__23941),
            .I(\b2v_inst11.g1 ));
    CascadeMux I__4318 (
            .O(N__23938),
            .I(\b2v_inst11.g1_cascade_ ));
    InMux I__4317 (
            .O(N__23935),
            .I(N__23929));
    InMux I__4316 (
            .O(N__23934),
            .I(N__23929));
    LocalMux I__4315 (
            .O(N__23929),
            .I(N__23926));
    Span4Mux_v I__4314 (
            .O(N__23926),
            .I(N__23923));
    Odrv4 I__4313 (
            .O(N__23923),
            .I(\b2v_inst11.g1_0 ));
    InMux I__4312 (
            .O(N__23920),
            .I(N__23914));
    InMux I__4311 (
            .O(N__23919),
            .I(N__23914));
    LocalMux I__4310 (
            .O(N__23914),
            .I(\b2v_inst11.dutycycleZ0Z_2 ));
    IoInMux I__4309 (
            .O(N__23911),
            .I(N__23908));
    LocalMux I__4308 (
            .O(N__23908),
            .I(N__23900));
    CascadeMux I__4307 (
            .O(N__23907),
            .I(N__23896));
    CascadeMux I__4306 (
            .O(N__23906),
            .I(N__23891));
    CascadeMux I__4305 (
            .O(N__23905),
            .I(N__23888));
    InMux I__4304 (
            .O(N__23904),
            .I(N__23881));
    InMux I__4303 (
            .O(N__23903),
            .I(N__23881));
    IoSpan4Mux I__4302 (
            .O(N__23900),
            .I(N__23871));
    InMux I__4301 (
            .O(N__23899),
            .I(N__23866));
    InMux I__4300 (
            .O(N__23896),
            .I(N__23866));
    InMux I__4299 (
            .O(N__23895),
            .I(N__23861));
    InMux I__4298 (
            .O(N__23894),
            .I(N__23861));
    InMux I__4297 (
            .O(N__23891),
            .I(N__23858));
    InMux I__4296 (
            .O(N__23888),
            .I(N__23854));
    InMux I__4295 (
            .O(N__23887),
            .I(N__23847));
    InMux I__4294 (
            .O(N__23886),
            .I(N__23847));
    LocalMux I__4293 (
            .O(N__23881),
            .I(N__23844));
    InMux I__4292 (
            .O(N__23880),
            .I(N__23841));
    InMux I__4291 (
            .O(N__23879),
            .I(N__23838));
    InMux I__4290 (
            .O(N__23878),
            .I(N__23830));
    InMux I__4289 (
            .O(N__23877),
            .I(N__23830));
    InMux I__4288 (
            .O(N__23876),
            .I(N__23825));
    InMux I__4287 (
            .O(N__23875),
            .I(N__23825));
    InMux I__4286 (
            .O(N__23874),
            .I(N__23822));
    Span4Mux_s0_h I__4285 (
            .O(N__23871),
            .I(N__23817));
    LocalMux I__4284 (
            .O(N__23866),
            .I(N__23817));
    LocalMux I__4283 (
            .O(N__23861),
            .I(N__23812));
    LocalMux I__4282 (
            .O(N__23858),
            .I(N__23812));
    InMux I__4281 (
            .O(N__23857),
            .I(N__23809));
    LocalMux I__4280 (
            .O(N__23854),
            .I(N__23806));
    InMux I__4279 (
            .O(N__23853),
            .I(N__23803));
    InMux I__4278 (
            .O(N__23852),
            .I(N__23800));
    LocalMux I__4277 (
            .O(N__23847),
            .I(N__23793));
    Span4Mux_v I__4276 (
            .O(N__23844),
            .I(N__23793));
    LocalMux I__4275 (
            .O(N__23841),
            .I(N__23793));
    LocalMux I__4274 (
            .O(N__23838),
            .I(N__23789));
    InMux I__4273 (
            .O(N__23837),
            .I(N__23782));
    InMux I__4272 (
            .O(N__23836),
            .I(N__23782));
    InMux I__4271 (
            .O(N__23835),
            .I(N__23782));
    LocalMux I__4270 (
            .O(N__23830),
            .I(N__23779));
    LocalMux I__4269 (
            .O(N__23825),
            .I(N__23776));
    LocalMux I__4268 (
            .O(N__23822),
            .I(N__23767));
    Span4Mux_h I__4267 (
            .O(N__23817),
            .I(N__23767));
    Span4Mux_v I__4266 (
            .O(N__23812),
            .I(N__23767));
    LocalMux I__4265 (
            .O(N__23809),
            .I(N__23767));
    Span4Mux_v I__4264 (
            .O(N__23806),
            .I(N__23758));
    LocalMux I__4263 (
            .O(N__23803),
            .I(N__23758));
    LocalMux I__4262 (
            .O(N__23800),
            .I(N__23758));
    Span4Mux_h I__4261 (
            .O(N__23793),
            .I(N__23758));
    InMux I__4260 (
            .O(N__23792),
            .I(N__23754));
    Span4Mux_v I__4259 (
            .O(N__23789),
            .I(N__23751));
    LocalMux I__4258 (
            .O(N__23782),
            .I(N__23748));
    Span4Mux_h I__4257 (
            .O(N__23779),
            .I(N__23745));
    Span4Mux_h I__4256 (
            .O(N__23776),
            .I(N__23738));
    Span4Mux_v I__4255 (
            .O(N__23767),
            .I(N__23738));
    Span4Mux_v I__4254 (
            .O(N__23758),
            .I(N__23738));
    InMux I__4253 (
            .O(N__23757),
            .I(N__23735));
    LocalMux I__4252 (
            .O(N__23754),
            .I(RSMRSTn_fast_RNIGMH81));
    Odrv4 I__4251 (
            .O(N__23751),
            .I(RSMRSTn_fast_RNIGMH81));
    Odrv12 I__4250 (
            .O(N__23748),
            .I(RSMRSTn_fast_RNIGMH81));
    Odrv4 I__4249 (
            .O(N__23745),
            .I(RSMRSTn_fast_RNIGMH81));
    Odrv4 I__4248 (
            .O(N__23738),
            .I(RSMRSTn_fast_RNIGMH81));
    LocalMux I__4247 (
            .O(N__23735),
            .I(RSMRSTn_fast_RNIGMH81));
    InMux I__4246 (
            .O(N__23722),
            .I(N__23717));
    InMux I__4245 (
            .O(N__23721),
            .I(N__23711));
    CascadeMux I__4244 (
            .O(N__23720),
            .I(N__23706));
    LocalMux I__4243 (
            .O(N__23717),
            .I(N__23690));
    InMux I__4242 (
            .O(N__23716),
            .I(N__23687));
    InMux I__4241 (
            .O(N__23715),
            .I(N__23684));
    InMux I__4240 (
            .O(N__23714),
            .I(N__23681));
    LocalMux I__4239 (
            .O(N__23711),
            .I(N__23678));
    InMux I__4238 (
            .O(N__23710),
            .I(N__23673));
    InMux I__4237 (
            .O(N__23709),
            .I(N__23673));
    InMux I__4236 (
            .O(N__23706),
            .I(N__23664));
    InMux I__4235 (
            .O(N__23705),
            .I(N__23664));
    InMux I__4234 (
            .O(N__23704),
            .I(N__23664));
    InMux I__4233 (
            .O(N__23703),
            .I(N__23657));
    InMux I__4232 (
            .O(N__23702),
            .I(N__23657));
    InMux I__4231 (
            .O(N__23701),
            .I(N__23657));
    InMux I__4230 (
            .O(N__23700),
            .I(N__23650));
    InMux I__4229 (
            .O(N__23699),
            .I(N__23650));
    InMux I__4228 (
            .O(N__23698),
            .I(N__23647));
    InMux I__4227 (
            .O(N__23697),
            .I(N__23640));
    InMux I__4226 (
            .O(N__23696),
            .I(N__23640));
    InMux I__4225 (
            .O(N__23695),
            .I(N__23640));
    InMux I__4224 (
            .O(N__23694),
            .I(N__23633));
    InMux I__4223 (
            .O(N__23693),
            .I(N__23633));
    Span4Mux_h I__4222 (
            .O(N__23690),
            .I(N__23619));
    LocalMux I__4221 (
            .O(N__23687),
            .I(N__23619));
    LocalMux I__4220 (
            .O(N__23684),
            .I(N__23619));
    LocalMux I__4219 (
            .O(N__23681),
            .I(N__23619));
    Span4Mux_v I__4218 (
            .O(N__23678),
            .I(N__23619));
    LocalMux I__4217 (
            .O(N__23673),
            .I(N__23619));
    InMux I__4216 (
            .O(N__23672),
            .I(N__23612));
    InMux I__4215 (
            .O(N__23671),
            .I(N__23612));
    LocalMux I__4214 (
            .O(N__23664),
            .I(N__23607));
    LocalMux I__4213 (
            .O(N__23657),
            .I(N__23607));
    InMux I__4212 (
            .O(N__23656),
            .I(N__23602));
    InMux I__4211 (
            .O(N__23655),
            .I(N__23602));
    LocalMux I__4210 (
            .O(N__23650),
            .I(N__23599));
    LocalMux I__4209 (
            .O(N__23647),
            .I(N__23596));
    LocalMux I__4208 (
            .O(N__23640),
            .I(N__23593));
    InMux I__4207 (
            .O(N__23639),
            .I(N__23588));
    InMux I__4206 (
            .O(N__23638),
            .I(N__23588));
    LocalMux I__4205 (
            .O(N__23633),
            .I(N__23584));
    InMux I__4204 (
            .O(N__23632),
            .I(N__23581));
    Span4Mux_v I__4203 (
            .O(N__23619),
            .I(N__23578));
    InMux I__4202 (
            .O(N__23618),
            .I(N__23573));
    InMux I__4201 (
            .O(N__23617),
            .I(N__23573));
    LocalMux I__4200 (
            .O(N__23612),
            .I(N__23568));
    Span12Mux_s11_v I__4199 (
            .O(N__23607),
            .I(N__23568));
    LocalMux I__4198 (
            .O(N__23602),
            .I(N__23563));
    Span4Mux_s3_h I__4197 (
            .O(N__23599),
            .I(N__23563));
    Span4Mux_s3_h I__4196 (
            .O(N__23596),
            .I(N__23560));
    Span4Mux_s3_h I__4195 (
            .O(N__23593),
            .I(N__23555));
    LocalMux I__4194 (
            .O(N__23588),
            .I(N__23555));
    InMux I__4193 (
            .O(N__23587),
            .I(N__23552));
    Odrv12 I__4192 (
            .O(N__23584),
            .I(func_state_RNI6BE8E_0_1));
    LocalMux I__4191 (
            .O(N__23581),
            .I(func_state_RNI6BE8E_0_1));
    Odrv4 I__4190 (
            .O(N__23578),
            .I(func_state_RNI6BE8E_0_1));
    LocalMux I__4189 (
            .O(N__23573),
            .I(func_state_RNI6BE8E_0_1));
    Odrv12 I__4188 (
            .O(N__23568),
            .I(func_state_RNI6BE8E_0_1));
    Odrv4 I__4187 (
            .O(N__23563),
            .I(func_state_RNI6BE8E_0_1));
    Odrv4 I__4186 (
            .O(N__23560),
            .I(func_state_RNI6BE8E_0_1));
    Odrv4 I__4185 (
            .O(N__23555),
            .I(func_state_RNI6BE8E_0_1));
    LocalMux I__4184 (
            .O(N__23552),
            .I(func_state_RNI6BE8E_0_1));
    CascadeMux I__4183 (
            .O(N__23533),
            .I(N__23528));
    CascadeMux I__4182 (
            .O(N__23532),
            .I(N__23525));
    CascadeMux I__4181 (
            .O(N__23531),
            .I(N__23522));
    InMux I__4180 (
            .O(N__23528),
            .I(N__23514));
    InMux I__4179 (
            .O(N__23525),
            .I(N__23514));
    InMux I__4178 (
            .O(N__23522),
            .I(N__23511));
    CascadeMux I__4177 (
            .O(N__23521),
            .I(N__23506));
    CascadeMux I__4176 (
            .O(N__23520),
            .I(N__23503));
    CascadeMux I__4175 (
            .O(N__23519),
            .I(N__23500));
    LocalMux I__4174 (
            .O(N__23514),
            .I(N__23496));
    LocalMux I__4173 (
            .O(N__23511),
            .I(N__23493));
    InMux I__4172 (
            .O(N__23510),
            .I(N__23490));
    InMux I__4171 (
            .O(N__23509),
            .I(N__23487));
    InMux I__4170 (
            .O(N__23506),
            .I(N__23484));
    InMux I__4169 (
            .O(N__23503),
            .I(N__23479));
    InMux I__4168 (
            .O(N__23500),
            .I(N__23476));
    InMux I__4167 (
            .O(N__23499),
            .I(N__23473));
    Span4Mux_h I__4166 (
            .O(N__23496),
            .I(N__23469));
    Span4Mux_h I__4165 (
            .O(N__23493),
            .I(N__23462));
    LocalMux I__4164 (
            .O(N__23490),
            .I(N__23462));
    LocalMux I__4163 (
            .O(N__23487),
            .I(N__23462));
    LocalMux I__4162 (
            .O(N__23484),
            .I(N__23459));
    InMux I__4161 (
            .O(N__23483),
            .I(N__23456));
    InMux I__4160 (
            .O(N__23482),
            .I(N__23453));
    LocalMux I__4159 (
            .O(N__23479),
            .I(N__23447));
    LocalMux I__4158 (
            .O(N__23476),
            .I(N__23447));
    LocalMux I__4157 (
            .O(N__23473),
            .I(N__23444));
    InMux I__4156 (
            .O(N__23472),
            .I(N__23441));
    Span4Mux_v I__4155 (
            .O(N__23469),
            .I(N__23430));
    Span4Mux_v I__4154 (
            .O(N__23462),
            .I(N__23430));
    Span4Mux_v I__4153 (
            .O(N__23459),
            .I(N__23430));
    LocalMux I__4152 (
            .O(N__23456),
            .I(N__23430));
    LocalMux I__4151 (
            .O(N__23453),
            .I(N__23430));
    InMux I__4150 (
            .O(N__23452),
            .I(N__23427));
    Span4Mux_h I__4149 (
            .O(N__23447),
            .I(N__23423));
    Span4Mux_h I__4148 (
            .O(N__23444),
            .I(N__23420));
    LocalMux I__4147 (
            .O(N__23441),
            .I(N__23417));
    Span4Mux_h I__4146 (
            .O(N__23430),
            .I(N__23414));
    LocalMux I__4145 (
            .O(N__23427),
            .I(N__23411));
    InMux I__4144 (
            .O(N__23426),
            .I(N__23408));
    Odrv4 I__4143 (
            .O(N__23423),
            .I(b2v_inst11_dutycycle_1_0_iv_0_o3_out));
    Odrv4 I__4142 (
            .O(N__23420),
            .I(b2v_inst11_dutycycle_1_0_iv_0_o3_out));
    Odrv12 I__4141 (
            .O(N__23417),
            .I(b2v_inst11_dutycycle_1_0_iv_0_o3_out));
    Odrv4 I__4140 (
            .O(N__23414),
            .I(b2v_inst11_dutycycle_1_0_iv_0_o3_out));
    Odrv12 I__4139 (
            .O(N__23411),
            .I(b2v_inst11_dutycycle_1_0_iv_0_o3_out));
    LocalMux I__4138 (
            .O(N__23408),
            .I(b2v_inst11_dutycycle_1_0_iv_0_o3_out));
    CascadeMux I__4137 (
            .O(N__23395),
            .I(N__23392));
    InMux I__4136 (
            .O(N__23392),
            .I(N__23383));
    InMux I__4135 (
            .O(N__23391),
            .I(N__23383));
    CascadeMux I__4134 (
            .O(N__23390),
            .I(N__23377));
    InMux I__4133 (
            .O(N__23389),
            .I(N__23370));
    InMux I__4132 (
            .O(N__23388),
            .I(N__23370));
    LocalMux I__4131 (
            .O(N__23383),
            .I(N__23367));
    InMux I__4130 (
            .O(N__23382),
            .I(N__23360));
    InMux I__4129 (
            .O(N__23381),
            .I(N__23360));
    InMux I__4128 (
            .O(N__23380),
            .I(N__23357));
    InMux I__4127 (
            .O(N__23377),
            .I(N__23353));
    InMux I__4126 (
            .O(N__23376),
            .I(N__23350));
    CascadeMux I__4125 (
            .O(N__23375),
            .I(N__23346));
    LocalMux I__4124 (
            .O(N__23370),
            .I(N__23343));
    Span4Mux_v I__4123 (
            .O(N__23367),
            .I(N__23340));
    InMux I__4122 (
            .O(N__23366),
            .I(N__23335));
    InMux I__4121 (
            .O(N__23365),
            .I(N__23335));
    LocalMux I__4120 (
            .O(N__23360),
            .I(N__23332));
    LocalMux I__4119 (
            .O(N__23357),
            .I(N__23329));
    InMux I__4118 (
            .O(N__23356),
            .I(N__23326));
    LocalMux I__4117 (
            .O(N__23353),
            .I(N__23323));
    LocalMux I__4116 (
            .O(N__23350),
            .I(N__23319));
    InMux I__4115 (
            .O(N__23349),
            .I(N__23316));
    InMux I__4114 (
            .O(N__23346),
            .I(N__23313));
    Span4Mux_v I__4113 (
            .O(N__23343),
            .I(N__23310));
    Span4Mux_h I__4112 (
            .O(N__23340),
            .I(N__23305));
    LocalMux I__4111 (
            .O(N__23335),
            .I(N__23305));
    Span4Mux_s3_h I__4110 (
            .O(N__23332),
            .I(N__23298));
    Span4Mux_h I__4109 (
            .O(N__23329),
            .I(N__23298));
    LocalMux I__4108 (
            .O(N__23326),
            .I(N__23298));
    Span4Mux_s3_h I__4107 (
            .O(N__23323),
            .I(N__23295));
    InMux I__4106 (
            .O(N__23322),
            .I(N__23292));
    Odrv12 I__4105 (
            .O(N__23319),
            .I(func_state_RNI_4_0));
    LocalMux I__4104 (
            .O(N__23316),
            .I(func_state_RNI_4_0));
    LocalMux I__4103 (
            .O(N__23313),
            .I(func_state_RNI_4_0));
    Odrv4 I__4102 (
            .O(N__23310),
            .I(func_state_RNI_4_0));
    Odrv4 I__4101 (
            .O(N__23305),
            .I(func_state_RNI_4_0));
    Odrv4 I__4100 (
            .O(N__23298),
            .I(func_state_RNI_4_0));
    Odrv4 I__4099 (
            .O(N__23295),
            .I(func_state_RNI_4_0));
    LocalMux I__4098 (
            .O(N__23292),
            .I(func_state_RNI_4_0));
    CascadeMux I__4097 (
            .O(N__23275),
            .I(N__23272));
    InMux I__4096 (
            .O(N__23272),
            .I(N__23266));
    InMux I__4095 (
            .O(N__23271),
            .I(N__23266));
    LocalMux I__4094 (
            .O(N__23266),
            .I(\b2v_inst11.dutycycleZ0Z_13 ));
    CascadeMux I__4093 (
            .O(N__23263),
            .I(\b2v_inst11.dutycycleZ0Z_5_cascade_ ));
    InMux I__4092 (
            .O(N__23260),
            .I(N__23256));
    InMux I__4091 (
            .O(N__23259),
            .I(N__23253));
    LocalMux I__4090 (
            .O(N__23256),
            .I(N__23248));
    LocalMux I__4089 (
            .O(N__23253),
            .I(N__23248));
    Span4Mux_h I__4088 (
            .O(N__23248),
            .I(N__23245));
    Odrv4 I__4087 (
            .O(N__23245),
            .I(\b2v_inst11.N_326_N ));
    InMux I__4086 (
            .O(N__23242),
            .I(N__23236));
    InMux I__4085 (
            .O(N__23241),
            .I(N__23236));
    LocalMux I__4084 (
            .O(N__23236),
            .I(N__23226));
    InMux I__4083 (
            .O(N__23235),
            .I(N__23221));
    InMux I__4082 (
            .O(N__23234),
            .I(N__23221));
    InMux I__4081 (
            .O(N__23233),
            .I(N__23216));
    InMux I__4080 (
            .O(N__23232),
            .I(N__23216));
    InMux I__4079 (
            .O(N__23231),
            .I(N__23211));
    InMux I__4078 (
            .O(N__23230),
            .I(N__23211));
    InMux I__4077 (
            .O(N__23229),
            .I(N__23208));
    Span4Mux_v I__4076 (
            .O(N__23226),
            .I(N__23205));
    LocalMux I__4075 (
            .O(N__23221),
            .I(N__23200));
    LocalMux I__4074 (
            .O(N__23216),
            .I(N__23200));
    LocalMux I__4073 (
            .O(N__23211),
            .I(N__23195));
    LocalMux I__4072 (
            .O(N__23208),
            .I(N__23195));
    Span4Mux_v I__4071 (
            .O(N__23205),
            .I(N__23192));
    Span4Mux_h I__4070 (
            .O(N__23200),
            .I(N__23187));
    Span4Mux_v I__4069 (
            .O(N__23195),
            .I(N__23187));
    Odrv4 I__4068 (
            .O(N__23192),
            .I(\b2v_inst11.N_140_N ));
    Odrv4 I__4067 (
            .O(N__23187),
            .I(\b2v_inst11.N_140_N ));
    InMux I__4066 (
            .O(N__23182),
            .I(N__23176));
    InMux I__4065 (
            .O(N__23181),
            .I(N__23168));
    InMux I__4064 (
            .O(N__23180),
            .I(N__23168));
    CascadeMux I__4063 (
            .O(N__23179),
            .I(N__23161));
    LocalMux I__4062 (
            .O(N__23176),
            .I(N__23158));
    InMux I__4061 (
            .O(N__23175),
            .I(N__23154));
    InMux I__4060 (
            .O(N__23174),
            .I(N__23149));
    InMux I__4059 (
            .O(N__23173),
            .I(N__23149));
    LocalMux I__4058 (
            .O(N__23168),
            .I(N__23146));
    InMux I__4057 (
            .O(N__23167),
            .I(N__23143));
    InMux I__4056 (
            .O(N__23166),
            .I(N__23136));
    InMux I__4055 (
            .O(N__23165),
            .I(N__23136));
    InMux I__4054 (
            .O(N__23164),
            .I(N__23136));
    InMux I__4053 (
            .O(N__23161),
            .I(N__23133));
    Span4Mux_v I__4052 (
            .O(N__23158),
            .I(N__23129));
    InMux I__4051 (
            .O(N__23157),
            .I(N__23126));
    LocalMux I__4050 (
            .O(N__23154),
            .I(N__23116));
    LocalMux I__4049 (
            .O(N__23149),
            .I(N__23116));
    Span4Mux_v I__4048 (
            .O(N__23146),
            .I(N__23116));
    LocalMux I__4047 (
            .O(N__23143),
            .I(N__23116));
    LocalMux I__4046 (
            .O(N__23136),
            .I(N__23113));
    LocalMux I__4045 (
            .O(N__23133),
            .I(N__23110));
    InMux I__4044 (
            .O(N__23132),
            .I(N__23107));
    Span4Mux_h I__4043 (
            .O(N__23129),
            .I(N__23102));
    LocalMux I__4042 (
            .O(N__23126),
            .I(N__23102));
    InMux I__4041 (
            .O(N__23125),
            .I(N__23099));
    Span4Mux_h I__4040 (
            .O(N__23116),
            .I(N__23092));
    Span4Mux_s3_h I__4039 (
            .O(N__23113),
            .I(N__23092));
    Span4Mux_s3_h I__4038 (
            .O(N__23110),
            .I(N__23092));
    LocalMux I__4037 (
            .O(N__23107),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__4036 (
            .O(N__23102),
            .I(\b2v_inst11.N_425 ));
    LocalMux I__4035 (
            .O(N__23099),
            .I(\b2v_inst11.N_425 ));
    Odrv4 I__4034 (
            .O(N__23092),
            .I(\b2v_inst11.N_425 ));
    CascadeMux I__4033 (
            .O(N__23083),
            .I(\b2v_inst11.N_154_N_cascade_ ));
    CascadeMux I__4032 (
            .O(N__23080),
            .I(\b2v_inst11.dutycycle_en_4_cascade_ ));
    InMux I__4031 (
            .O(N__23077),
            .I(N__23071));
    InMux I__4030 (
            .O(N__23076),
            .I(N__23071));
    LocalMux I__4029 (
            .O(N__23071),
            .I(\b2v_inst11.dutycycle_e_1_8 ));
    InMux I__4028 (
            .O(N__23068),
            .I(N__23062));
    InMux I__4027 (
            .O(N__23067),
            .I(N__23048));
    InMux I__4026 (
            .O(N__23066),
            .I(N__23038));
    InMux I__4025 (
            .O(N__23065),
            .I(N__23038));
    LocalMux I__4024 (
            .O(N__23062),
            .I(N__23035));
    InMux I__4023 (
            .O(N__23061),
            .I(N__23032));
    InMux I__4022 (
            .O(N__23060),
            .I(N__23027));
    InMux I__4021 (
            .O(N__23059),
            .I(N__23027));
    CascadeMux I__4020 (
            .O(N__23058),
            .I(N__23022));
    InMux I__4019 (
            .O(N__23057),
            .I(N__23019));
    InMux I__4018 (
            .O(N__23056),
            .I(N__23012));
    InMux I__4017 (
            .O(N__23055),
            .I(N__23012));
    InMux I__4016 (
            .O(N__23054),
            .I(N__23012));
    InMux I__4015 (
            .O(N__23053),
            .I(N__23005));
    InMux I__4014 (
            .O(N__23052),
            .I(N__23005));
    InMux I__4013 (
            .O(N__23051),
            .I(N__23005));
    LocalMux I__4012 (
            .O(N__23048),
            .I(N__23002));
    InMux I__4011 (
            .O(N__23047),
            .I(N__22997));
    InMux I__4010 (
            .O(N__23046),
            .I(N__22997));
    InMux I__4009 (
            .O(N__23045),
            .I(N__22992));
    InMux I__4008 (
            .O(N__23044),
            .I(N__22992));
    CascadeMux I__4007 (
            .O(N__23043),
            .I(N__22988));
    LocalMux I__4006 (
            .O(N__23038),
            .I(N__22983));
    Span4Mux_s3_h I__4005 (
            .O(N__23035),
            .I(N__22976));
    LocalMux I__4004 (
            .O(N__23032),
            .I(N__22976));
    LocalMux I__4003 (
            .O(N__23027),
            .I(N__22976));
    InMux I__4002 (
            .O(N__23026),
            .I(N__22971));
    InMux I__4001 (
            .O(N__23025),
            .I(N__22971));
    InMux I__4000 (
            .O(N__23022),
            .I(N__22968));
    LocalMux I__3999 (
            .O(N__23019),
            .I(N__22961));
    LocalMux I__3998 (
            .O(N__23012),
            .I(N__22961));
    LocalMux I__3997 (
            .O(N__23005),
            .I(N__22961));
    Span4Mux_h I__3996 (
            .O(N__23002),
            .I(N__22954));
    LocalMux I__3995 (
            .O(N__22997),
            .I(N__22954));
    LocalMux I__3994 (
            .O(N__22992),
            .I(N__22954));
    InMux I__3993 (
            .O(N__22991),
            .I(N__22947));
    InMux I__3992 (
            .O(N__22988),
            .I(N__22947));
    InMux I__3991 (
            .O(N__22987),
            .I(N__22947));
    InMux I__3990 (
            .O(N__22986),
            .I(N__22944));
    Span4Mux_v I__3989 (
            .O(N__22983),
            .I(N__22937));
    Span4Mux_v I__3988 (
            .O(N__22976),
            .I(N__22937));
    LocalMux I__3987 (
            .O(N__22971),
            .I(N__22937));
    LocalMux I__3986 (
            .O(N__22968),
            .I(N__22930));
    Span4Mux_h I__3985 (
            .O(N__22961),
            .I(N__22930));
    Span4Mux_v I__3984 (
            .O(N__22954),
            .I(N__22930));
    LocalMux I__3983 (
            .O(N__22947),
            .I(N__22925));
    LocalMux I__3982 (
            .O(N__22944),
            .I(N__22925));
    Span4Mux_h I__3981 (
            .O(N__22937),
            .I(N__22922));
    Odrv4 I__3980 (
            .O(N__22930),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv12 I__3979 (
            .O(N__22925),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    Odrv4 I__3978 (
            .O(N__22922),
            .I(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ));
    InMux I__3977 (
            .O(N__22915),
            .I(N__22912));
    LocalMux I__3976 (
            .O(N__22912),
            .I(\b2v_inst11.dutycycle_en_4 ));
    InMux I__3975 (
            .O(N__22909),
            .I(N__22903));
    InMux I__3974 (
            .O(N__22908),
            .I(N__22903));
    LocalMux I__3973 (
            .O(N__22903),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69 ));
    CascadeMux I__3972 (
            .O(N__22900),
            .I(N__22897));
    InMux I__3971 (
            .O(N__22897),
            .I(N__22893));
    InMux I__3970 (
            .O(N__22896),
            .I(N__22890));
    LocalMux I__3969 (
            .O(N__22893),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    LocalMux I__3968 (
            .O(N__22890),
            .I(\b2v_inst11.dutycycleZ0Z_10 ));
    CascadeMux I__3967 (
            .O(N__22885),
            .I(N__22882));
    InMux I__3966 (
            .O(N__22882),
            .I(N__22873));
    InMux I__3965 (
            .O(N__22881),
            .I(N__22873));
    InMux I__3964 (
            .O(N__22880),
            .I(N__22873));
    LocalMux I__3963 (
            .O(N__22873),
            .I(\b2v_inst11.dutycycleZ1Z_8 ));
    InMux I__3962 (
            .O(N__22870),
            .I(N__22867));
    LocalMux I__3961 (
            .O(N__22867),
            .I(N__22864));
    Odrv4 I__3960 (
            .O(N__22864),
            .I(\b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49 ));
    CascadeMux I__3959 (
            .O(N__22861),
            .I(N__22858));
    InMux I__3958 (
            .O(N__22858),
            .I(N__22852));
    InMux I__3957 (
            .O(N__22857),
            .I(N__22852));
    LocalMux I__3956 (
            .O(N__22852),
            .I(\b2v_inst11.dutycycle_RNI1KT13Z0Z_8 ));
    InMux I__3955 (
            .O(N__22849),
            .I(N__22846));
    LocalMux I__3954 (
            .O(N__22846),
            .I(\b2v_inst11.dutycycle_RNI_1Z0Z_3 ));
    CascadeMux I__3953 (
            .O(N__22843),
            .I(\b2v_inst11.dutycycleZ0Z_8_cascade_ ));
    CascadeMux I__3952 (
            .O(N__22840),
            .I(\b2v_inst11.N_153_N_cascade_ ));
    CascadeMux I__3951 (
            .O(N__22837),
            .I(\b2v_inst11.N_156_N_cascade_ ));
    InMux I__3950 (
            .O(N__22834),
            .I(N__22831));
    LocalMux I__3949 (
            .O(N__22831),
            .I(\b2v_inst11.dutycycle_e_1_9 ));
    CascadeMux I__3948 (
            .O(N__22828),
            .I(N__22825));
    InMux I__3947 (
            .O(N__22825),
            .I(N__22821));
    InMux I__3946 (
            .O(N__22824),
            .I(N__22818));
    LocalMux I__3945 (
            .O(N__22821),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ));
    LocalMux I__3944 (
            .O(N__22818),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ));
    CascadeMux I__3943 (
            .O(N__22813),
            .I(\b2v_inst11.dutycycle_e_1_9_cascade_ ));
    InMux I__3942 (
            .O(N__22810),
            .I(N__22804));
    InMux I__3941 (
            .O(N__22809),
            .I(N__22804));
    LocalMux I__3940 (
            .O(N__22804),
            .I(\b2v_inst11.dutycycleZ1Z_9 ));
    CascadeMux I__3939 (
            .O(N__22801),
            .I(N__22798));
    InMux I__3938 (
            .O(N__22798),
            .I(N__22792));
    InMux I__3937 (
            .O(N__22797),
            .I(N__22792));
    LocalMux I__3936 (
            .O(N__22792),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ));
    InMux I__3935 (
            .O(N__22789),
            .I(N__22783));
    InMux I__3934 (
            .O(N__22788),
            .I(N__22783));
    LocalMux I__3933 (
            .O(N__22783),
            .I(\b2v_inst11.dutycycle_en_10 ));
    InMux I__3932 (
            .O(N__22780),
            .I(N__22777));
    LocalMux I__3931 (
            .O(N__22777),
            .I(\b2v_inst5.count_rst_10 ));
    CascadeMux I__3930 (
            .O(N__22774),
            .I(\b2v_inst5.countZ0Z_8_cascade_ ));
    InMux I__3929 (
            .O(N__22771),
            .I(N__22765));
    InMux I__3928 (
            .O(N__22770),
            .I(N__22765));
    LocalMux I__3927 (
            .O(N__22765),
            .I(\b2v_inst5.count_1_4 ));
    CascadeMux I__3926 (
            .O(N__22762),
            .I(\b2v_inst5.un12_clk_100khz_7_cascade_ ));
    CascadeMux I__3925 (
            .O(N__22759),
            .I(\b2v_inst11.N_8_1_cascade_ ));
    InMux I__3924 (
            .O(N__22756),
            .I(N__22753));
    LocalMux I__3923 (
            .O(N__22753),
            .I(N__22750));
    Span4Mux_v I__3922 (
            .O(N__22750),
            .I(N__22747));
    Odrv4 I__3921 (
            .O(N__22747),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_8 ));
    CascadeMux I__3920 (
            .O(N__22744),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_ ));
    InMux I__3919 (
            .O(N__22741),
            .I(N__22738));
    LocalMux I__3918 (
            .O(N__22738),
            .I(N__22734));
    InMux I__3917 (
            .O(N__22737),
            .I(N__22731));
    Odrv4 I__3916 (
            .O(N__22734),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ));
    LocalMux I__3915 (
            .O(N__22731),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ));
    InMux I__3914 (
            .O(N__22726),
            .I(N__22723));
    LocalMux I__3913 (
            .O(N__22723),
            .I(N__22720));
    Odrv4 I__3912 (
            .O(N__22720),
            .I(\b2v_inst11.dutycycle_en_11 ));
    CascadeMux I__3911 (
            .O(N__22717),
            .I(N__22714));
    InMux I__3910 (
            .O(N__22714),
            .I(N__22711));
    LocalMux I__3909 (
            .O(N__22711),
            .I(N__22707));
    InMux I__3908 (
            .O(N__22710),
            .I(N__22704));
    Span4Mux_h I__3907 (
            .O(N__22707),
            .I(N__22701));
    LocalMux I__3906 (
            .O(N__22704),
            .I(\b2v_inst11.dutycycleZ0Z_14 ));
    Odrv4 I__3905 (
            .O(N__22701),
            .I(\b2v_inst11.dutycycleZ0Z_14 ));
    CascadeMux I__3904 (
            .O(N__22696),
            .I(\b2v_inst11.dutycycleZ0Z_12_cascade_ ));
    InMux I__3903 (
            .O(N__22693),
            .I(N__22690));
    LocalMux I__3902 (
            .O(N__22690),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ));
    InMux I__3901 (
            .O(N__22687),
            .I(N__22683));
    InMux I__3900 (
            .O(N__22686),
            .I(N__22680));
    LocalMux I__3899 (
            .O(N__22683),
            .I(N__22677));
    LocalMux I__3898 (
            .O(N__22680),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_9 ));
    Odrv4 I__3897 (
            .O(N__22677),
            .I(\b2v_inst11.dutycycle_RNI_4Z0Z_9 ));
    InMux I__3896 (
            .O(N__22672),
            .I(N__22668));
    InMux I__3895 (
            .O(N__22671),
            .I(N__22665));
    LocalMux I__3894 (
            .O(N__22668),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    LocalMux I__3893 (
            .O(N__22665),
            .I(\b2v_inst11.mult1_un124_sum_cry_3_s ));
    CascadeMux I__3892 (
            .O(N__22660),
            .I(N__22657));
    InMux I__3891 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__3890 (
            .O(N__22654),
            .I(N__22651));
    Odrv4 I__3889 (
            .O(N__22651),
            .I(\b2v_inst11.mult1_un131_sum_axb_4_l_fx ));
    InMux I__3888 (
            .O(N__22648),
            .I(N__22645));
    LocalMux I__3887 (
            .O(N__22645),
            .I(\b2v_inst11.g0_13_1 ));
    CascadeMux I__3886 (
            .O(N__22642),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_9_cascade_ ));
    InMux I__3885 (
            .O(N__22639),
            .I(N__22636));
    LocalMux I__3884 (
            .O(N__22636),
            .I(N__22633));
    Span4Mux_v I__3883 (
            .O(N__22633),
            .I(N__22630));
    Odrv4 I__3882 (
            .O(N__22630),
            .I(\b2v_inst200.count_RNIC03N_6Z0Z_0 ));
    InMux I__3881 (
            .O(N__22627),
            .I(N__22624));
    LocalMux I__3880 (
            .O(N__22624),
            .I(N__22620));
    InMux I__3879 (
            .O(N__22623),
            .I(N__22617));
    Span4Mux_v I__3878 (
            .O(N__22620),
            .I(N__22614));
    LocalMux I__3877 (
            .O(N__22617),
            .I(N__22611));
    Span4Mux_v I__3876 (
            .O(N__22614),
            .I(N__22608));
    Span12Mux_s5_h I__3875 (
            .O(N__22611),
            .I(N__22605));
    Odrv4 I__3874 (
            .O(N__22608),
            .I(N_411));
    Odrv12 I__3873 (
            .O(N__22605),
            .I(N_411));
    CascadeMux I__3872 (
            .O(N__22600),
            .I(N__22597));
    InMux I__3871 (
            .O(N__22597),
            .I(N__22590));
    InMux I__3870 (
            .O(N__22596),
            .I(N__22590));
    InMux I__3869 (
            .O(N__22595),
            .I(N__22587));
    LocalMux I__3868 (
            .O(N__22590),
            .I(N__22582));
    LocalMux I__3867 (
            .O(N__22587),
            .I(N__22582));
    Span4Mux_h I__3866 (
            .O(N__22582),
            .I(N__22579));
    Span4Mux_v I__3865 (
            .O(N__22579),
            .I(N__22576));
    Span4Mux_v I__3864 (
            .O(N__22576),
            .I(N__22573));
    Odrv4 I__3863 (
            .O(N__22573),
            .I(\b2v_inst200.m11_0_a3_0 ));
    CascadeMux I__3862 (
            .O(N__22570),
            .I(\b2v_inst5.count_rst_10_cascade_ ));
    CascadeMux I__3861 (
            .O(N__22567),
            .I(\b2v_inst5.un2_count_1_axb_4_cascade_ ));
    InMux I__3860 (
            .O(N__22564),
            .I(N__22561));
    LocalMux I__3859 (
            .O(N__22561),
            .I(\b2v_inst5.count_1_8 ));
    CascadeMux I__3858 (
            .O(N__22558),
            .I(N__22555));
    InMux I__3857 (
            .O(N__22555),
            .I(N__22552));
    LocalMux I__3856 (
            .O(N__22552),
            .I(\b2v_inst11.mult1_un124_sum_cry_4_s ));
    InMux I__3855 (
            .O(N__22549),
            .I(\b2v_inst11.mult1_un124_sum_cry_3 ));
    InMux I__3854 (
            .O(N__22546),
            .I(N__22543));
    LocalMux I__3853 (
            .O(N__22543),
            .I(\b2v_inst11.mult1_un124_sum_cry_5_s ));
    InMux I__3852 (
            .O(N__22540),
            .I(\b2v_inst11.mult1_un124_sum_cry_4 ));
    InMux I__3851 (
            .O(N__22537),
            .I(N__22531));
    InMux I__3850 (
            .O(N__22536),
            .I(N__22531));
    LocalMux I__3849 (
            .O(N__22531),
            .I(\b2v_inst11.mult1_un124_sum_cry_6_s ));
    InMux I__3848 (
            .O(N__22528),
            .I(\b2v_inst11.mult1_un124_sum_cry_5 ));
    CascadeMux I__3847 (
            .O(N__22525),
            .I(N__22522));
    InMux I__3846 (
            .O(N__22522),
            .I(N__22519));
    LocalMux I__3845 (
            .O(N__22519),
            .I(\b2v_inst11.mult1_un131_sum_axb_8 ));
    InMux I__3844 (
            .O(N__22516),
            .I(\b2v_inst11.mult1_un124_sum_cry_6 ));
    InMux I__3843 (
            .O(N__22513),
            .I(\b2v_inst11.mult1_un124_sum_cry_7 ));
    CascadeMux I__3842 (
            .O(N__22510),
            .I(\b2v_inst11.mult1_un124_sum_s_8_cascade_ ));
    CascadeMux I__3841 (
            .O(N__22507),
            .I(N__22504));
    InMux I__3840 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__3839 (
            .O(N__22501),
            .I(\b2v_inst11.mult1_un124_sum_i_0_8 ));
    InMux I__3838 (
            .O(N__22498),
            .I(N__22493));
    InMux I__3837 (
            .O(N__22497),
            .I(N__22490));
    InMux I__3836 (
            .O(N__22496),
            .I(N__22487));
    LocalMux I__3835 (
            .O(N__22493),
            .I(N__22484));
    LocalMux I__3834 (
            .O(N__22490),
            .I(N__22480));
    LocalMux I__3833 (
            .O(N__22487),
            .I(N__22477));
    Sp12to4 I__3832 (
            .O(N__22484),
            .I(N__22474));
    InMux I__3831 (
            .O(N__22483),
            .I(N__22471));
    Span4Mux_h I__3830 (
            .O(N__22480),
            .I(N__22468));
    Span4Mux_h I__3829 (
            .O(N__22477),
            .I(N__22465));
    Odrv12 I__3828 (
            .O(N__22474),
            .I(\b2v_inst11.N_382 ));
    LocalMux I__3827 (
            .O(N__22471),
            .I(\b2v_inst11.N_382 ));
    Odrv4 I__3826 (
            .O(N__22468),
            .I(\b2v_inst11.N_382 ));
    Odrv4 I__3825 (
            .O(N__22465),
            .I(\b2v_inst11.N_382 ));
    CascadeMux I__3824 (
            .O(N__22456),
            .I(N__22453));
    InMux I__3823 (
            .O(N__22453),
            .I(N__22450));
    LocalMux I__3822 (
            .O(N__22450),
            .I(N__22447));
    Odrv4 I__3821 (
            .O(N__22447),
            .I(\b2v_inst11.N_302 ));
    InMux I__3820 (
            .O(N__22444),
            .I(\b2v_inst11.mult1_un131_sum_cry_2 ));
    InMux I__3819 (
            .O(N__22441),
            .I(\b2v_inst11.mult1_un131_sum_cry_3 ));
    InMux I__3818 (
            .O(N__22438),
            .I(\b2v_inst11.mult1_un131_sum_cry_4 ));
    InMux I__3817 (
            .O(N__22435),
            .I(\b2v_inst11.mult1_un131_sum_cry_5 ));
    InMux I__3816 (
            .O(N__22432),
            .I(\b2v_inst11.mult1_un131_sum_cry_6 ));
    InMux I__3815 (
            .O(N__22429),
            .I(\b2v_inst11.mult1_un131_sum_cry_7 ));
    CascadeMux I__3814 (
            .O(N__22426),
            .I(N__22423));
    InMux I__3813 (
            .O(N__22423),
            .I(N__22420));
    LocalMux I__3812 (
            .O(N__22420),
            .I(\b2v_inst11.mult1_un131_sum_axb_7_l_fx ));
    InMux I__3811 (
            .O(N__22417),
            .I(\b2v_inst11.mult1_un124_sum_cry_2 ));
    InMux I__3810 (
            .O(N__22414),
            .I(N__22411));
    LocalMux I__3809 (
            .O(N__22411),
            .I(\b2v_inst36.DSW_PWROK_0 ));
    InMux I__3808 (
            .O(N__22408),
            .I(N__22405));
    LocalMux I__3807 (
            .O(N__22405),
            .I(\b2v_inst36.curr_state_0_0 ));
    CascadeMux I__3806 (
            .O(N__22402),
            .I(\b2v_inst36.curr_state_7_0_cascade_ ));
    CascadeMux I__3805 (
            .O(N__22399),
            .I(N__22394));
    InMux I__3804 (
            .O(N__22398),
            .I(N__22390));
    InMux I__3803 (
            .O(N__22397),
            .I(N__22383));
    InMux I__3802 (
            .O(N__22394),
            .I(N__22383));
    InMux I__3801 (
            .O(N__22393),
            .I(N__22383));
    LocalMux I__3800 (
            .O(N__22390),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    LocalMux I__3799 (
            .O(N__22383),
            .I(\b2v_inst36.curr_stateZ0Z_0 ));
    CascadeMux I__3798 (
            .O(N__22378),
            .I(\b2v_inst36.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__3797 (
            .O(N__22375),
            .I(\b2v_inst36.N_2939_i_cascade_ ));
    InMux I__3796 (
            .O(N__22372),
            .I(N__22369));
    LocalMux I__3795 (
            .O(N__22369),
            .I(\b2v_inst36.count_2_4 ));
    InMux I__3794 (
            .O(N__22366),
            .I(N__22363));
    LocalMux I__3793 (
            .O(N__22363),
            .I(\b2v_inst36.count_2_9 ));
    InMux I__3792 (
            .O(N__22360),
            .I(N__22357));
    LocalMux I__3791 (
            .O(N__22357),
            .I(\b2v_inst36.count_2_12 ));
    CascadeMux I__3790 (
            .O(N__22354),
            .I(\b2v_inst36.curr_state_RNI8TT2Z0Z_0_cascade_ ));
    IoInMux I__3789 (
            .O(N__22351),
            .I(N__22348));
    LocalMux I__3788 (
            .O(N__22348),
            .I(N__22345));
    IoSpan4Mux I__3787 (
            .O(N__22345),
            .I(N__22342));
    Span4Mux_s2_h I__3786 (
            .O(N__22342),
            .I(N__22339));
    Span4Mux_h I__3785 (
            .O(N__22339),
            .I(N__22336));
    Odrv4 I__3784 (
            .O(N__22336),
            .I(DSW_PWROK_c));
    CascadeMux I__3783 (
            .O(N__22333),
            .I(\b2v_inst200.curr_stateZ0Z_1_cascade_ ));
    InMux I__3782 (
            .O(N__22330),
            .I(N__22326));
    CascadeMux I__3781 (
            .O(N__22329),
            .I(N__22319));
    LocalMux I__3780 (
            .O(N__22326),
            .I(N__22314));
    InMux I__3779 (
            .O(N__22325),
            .I(N__22296));
    InMux I__3778 (
            .O(N__22324),
            .I(N__22296));
    InMux I__3777 (
            .O(N__22323),
            .I(N__22296));
    InMux I__3776 (
            .O(N__22322),
            .I(N__22296));
    InMux I__3775 (
            .O(N__22319),
            .I(N__22296));
    InMux I__3774 (
            .O(N__22318),
            .I(N__22296));
    InMux I__3773 (
            .O(N__22317),
            .I(N__22293));
    Span12Mux_s7_v I__3772 (
            .O(N__22314),
            .I(N__22290));
    InMux I__3771 (
            .O(N__22313),
            .I(N__22287));
    InMux I__3770 (
            .O(N__22312),
            .I(N__22278));
    InMux I__3769 (
            .O(N__22311),
            .I(N__22278));
    InMux I__3768 (
            .O(N__22310),
            .I(N__22278));
    InMux I__3767 (
            .O(N__22309),
            .I(N__22278));
    LocalMux I__3766 (
            .O(N__22296),
            .I(N__22273));
    LocalMux I__3765 (
            .O(N__22293),
            .I(N__22273));
    Odrv12 I__3764 (
            .O(N__22290),
            .I(\b2v_inst200.count_RNI_0_0 ));
    LocalMux I__3763 (
            .O(N__22287),
            .I(\b2v_inst200.count_RNI_0_0 ));
    LocalMux I__3762 (
            .O(N__22278),
            .I(\b2v_inst200.count_RNI_0_0 ));
    Odrv4 I__3761 (
            .O(N__22273),
            .I(\b2v_inst200.count_RNI_0_0 ));
    InMux I__3760 (
            .O(N__22264),
            .I(N__22261));
    LocalMux I__3759 (
            .O(N__22261),
            .I(N__22258));
    Span4Mux_h I__3758 (
            .O(N__22258),
            .I(N__22255));
    Odrv4 I__3757 (
            .O(N__22255),
            .I(GPIO_FPGA_SoC_1_c));
    CascadeMux I__3756 (
            .O(N__22252),
            .I(N_411_cascade_));
    InMux I__3755 (
            .O(N__22249),
            .I(N__22246));
    LocalMux I__3754 (
            .O(N__22246),
            .I(\b2v_inst200.m6_i_0 ));
    CascadeMux I__3753 (
            .O(N__22243),
            .I(\b2v_inst200.m6_i_0_cascade_ ));
    InMux I__3752 (
            .O(N__22240),
            .I(N__22237));
    LocalMux I__3751 (
            .O(N__22237),
            .I(\b2v_inst200.curr_state_3_0 ));
    CascadeMux I__3750 (
            .O(N__22234),
            .I(\b2v_inst200.N_58_cascade_ ));
    InMux I__3749 (
            .O(N__22231),
            .I(N__22220));
    InMux I__3748 (
            .O(N__22230),
            .I(N__22220));
    InMux I__3747 (
            .O(N__22229),
            .I(N__22220));
    InMux I__3746 (
            .O(N__22228),
            .I(N__22215));
    InMux I__3745 (
            .O(N__22227),
            .I(N__22215));
    LocalMux I__3744 (
            .O(N__22220),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    LocalMux I__3743 (
            .O(N__22215),
            .I(\b2v_inst200.curr_stateZ0Z_0 ));
    CascadeMux I__3742 (
            .O(N__22210),
            .I(\b2v_inst200.curr_stateZ0Z_0_cascade_ ));
    InMux I__3741 (
            .O(N__22207),
            .I(N__22201));
    InMux I__3740 (
            .O(N__22206),
            .I(N__22201));
    LocalMux I__3739 (
            .O(N__22201),
            .I(N_412));
    CascadeMux I__3738 (
            .O(N__22198),
            .I(N_412_cascade_));
    CascadeMux I__3737 (
            .O(N__22195),
            .I(N__22187));
    InMux I__3736 (
            .O(N__22194),
            .I(N__22181));
    InMux I__3735 (
            .O(N__22193),
            .I(N__22181));
    InMux I__3734 (
            .O(N__22192),
            .I(N__22176));
    InMux I__3733 (
            .O(N__22191),
            .I(N__22176));
    InMux I__3732 (
            .O(N__22190),
            .I(N__22169));
    InMux I__3731 (
            .O(N__22187),
            .I(N__22169));
    InMux I__3730 (
            .O(N__22186),
            .I(N__22169));
    LocalMux I__3729 (
            .O(N__22181),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__3728 (
            .O(N__22176),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    LocalMux I__3727 (
            .O(N__22169),
            .I(\b2v_inst200.curr_stateZ0Z_1 ));
    InMux I__3726 (
            .O(N__22162),
            .I(N__22159));
    LocalMux I__3725 (
            .O(N__22159),
            .I(\b2v_inst200.curr_state_3_1 ));
    InMux I__3724 (
            .O(N__22156),
            .I(N__22153));
    LocalMux I__3723 (
            .O(N__22153),
            .I(\b2v_inst36.count_2_6 ));
    InMux I__3722 (
            .O(N__22150),
            .I(N__22147));
    LocalMux I__3721 (
            .O(N__22147),
            .I(\b2v_inst11.count_0_9 ));
    InMux I__3720 (
            .O(N__22144),
            .I(N__22141));
    LocalMux I__3719 (
            .O(N__22141),
            .I(\b2v_inst11.count_0_10 ));
    InMux I__3718 (
            .O(N__22138),
            .I(N__22135));
    LocalMux I__3717 (
            .O(N__22135),
            .I(\b2v_inst11.count_0_11 ));
    InMux I__3716 (
            .O(N__22132),
            .I(N__22129));
    LocalMux I__3715 (
            .O(N__22129),
            .I(\b2v_inst11.count_0_2 ));
    CascadeMux I__3714 (
            .O(N__22126),
            .I(\b2v_inst200.N_56_cascade_ ));
    CascadeMux I__3713 (
            .O(N__22123),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1_cascade_ ));
    InMux I__3712 (
            .O(N__22120),
            .I(N__22116));
    InMux I__3711 (
            .O(N__22119),
            .I(N__22110));
    LocalMux I__3710 (
            .O(N__22116),
            .I(N__22107));
    InMux I__3709 (
            .O(N__22115),
            .I(N__22104));
    InMux I__3708 (
            .O(N__22114),
            .I(N__22099));
    InMux I__3707 (
            .O(N__22113),
            .I(N__22099));
    LocalMux I__3706 (
            .O(N__22110),
            .I(N__22090));
    Span4Mux_v I__3705 (
            .O(N__22107),
            .I(N__22087));
    LocalMux I__3704 (
            .O(N__22104),
            .I(N__22084));
    LocalMux I__3703 (
            .O(N__22099),
            .I(N__22081));
    InMux I__3702 (
            .O(N__22098),
            .I(N__22074));
    InMux I__3701 (
            .O(N__22097),
            .I(N__22074));
    InMux I__3700 (
            .O(N__22096),
            .I(N__22074));
    InMux I__3699 (
            .O(N__22095),
            .I(N__22067));
    InMux I__3698 (
            .O(N__22094),
            .I(N__22067));
    InMux I__3697 (
            .O(N__22093),
            .I(N__22067));
    Span4Mux_s2_v I__3696 (
            .O(N__22090),
            .I(N__22060));
    Span4Mux_v I__3695 (
            .O(N__22087),
            .I(N__22060));
    Span4Mux_v I__3694 (
            .O(N__22084),
            .I(N__22055));
    Span4Mux_h I__3693 (
            .O(N__22081),
            .I(N__22055));
    LocalMux I__3692 (
            .O(N__22074),
            .I(N__22050));
    LocalMux I__3691 (
            .O(N__22067),
            .I(N__22050));
    InMux I__3690 (
            .O(N__22066),
            .I(N__22045));
    InMux I__3689 (
            .O(N__22065),
            .I(N__22045));
    Odrv4 I__3688 (
            .O(N__22060),
            .I(b2v_inst5_RSMRSTn_latmux));
    Odrv4 I__3687 (
            .O(N__22055),
            .I(b2v_inst5_RSMRSTn_latmux));
    Odrv4 I__3686 (
            .O(N__22050),
            .I(b2v_inst5_RSMRSTn_latmux));
    LocalMux I__3685 (
            .O(N__22045),
            .I(b2v_inst5_RSMRSTn_latmux));
    InMux I__3684 (
            .O(N__22036),
            .I(N__22032));
    InMux I__3683 (
            .O(N__22035),
            .I(N__22028));
    LocalMux I__3682 (
            .O(N__22032),
            .I(N__22025));
    InMux I__3681 (
            .O(N__22031),
            .I(N__22022));
    LocalMux I__3680 (
            .O(N__22028),
            .I(N__22018));
    Span4Mux_h I__3679 (
            .O(N__22025),
            .I(N__22013));
    LocalMux I__3678 (
            .O(N__22022),
            .I(N__22013));
    CascadeMux I__3677 (
            .O(N__22021),
            .I(N__22010));
    Span12Mux_s5_h I__3676 (
            .O(N__22018),
            .I(N__22006));
    Span4Mux_v I__3675 (
            .O(N__22013),
            .I(N__22003));
    InMux I__3674 (
            .O(N__22010),
            .I(N__21998));
    InMux I__3673 (
            .O(N__22009),
            .I(N__21998));
    Odrv12 I__3672 (
            .O(N__22006),
            .I(b2v_inst5_RSMRSTn_fast));
    Odrv4 I__3671 (
            .O(N__22003),
            .I(b2v_inst5_RSMRSTn_fast));
    LocalMux I__3670 (
            .O(N__21998),
            .I(b2v_inst5_RSMRSTn_fast));
    InMux I__3669 (
            .O(N__21991),
            .I(N__21988));
    LocalMux I__3668 (
            .O(N__21988),
            .I(N__21983));
    InMux I__3667 (
            .O(N__21987),
            .I(N__21980));
    CascadeMux I__3666 (
            .O(N__21986),
            .I(N__21974));
    Span4Mux_s2_v I__3665 (
            .O(N__21983),
            .I(N__21969));
    LocalMux I__3664 (
            .O(N__21980),
            .I(N__21969));
    InMux I__3663 (
            .O(N__21979),
            .I(N__21966));
    InMux I__3662 (
            .O(N__21978),
            .I(N__21959));
    InMux I__3661 (
            .O(N__21977),
            .I(N__21959));
    InMux I__3660 (
            .O(N__21974),
            .I(N__21959));
    Span4Mux_v I__3659 (
            .O(N__21969),
            .I(N__21956));
    LocalMux I__3658 (
            .O(N__21966),
            .I(N__21951));
    LocalMux I__3657 (
            .O(N__21959),
            .I(N__21951));
    Odrv4 I__3656 (
            .O(N__21956),
            .I(RSMRSTn_0));
    Odrv4 I__3655 (
            .O(N__21951),
            .I(RSMRSTn_0));
    InMux I__3654 (
            .O(N__21946),
            .I(N__21939));
    InMux I__3653 (
            .O(N__21945),
            .I(N__21939));
    InMux I__3652 (
            .O(N__21944),
            .I(N__21936));
    LocalMux I__3651 (
            .O(N__21939),
            .I(N__21933));
    LocalMux I__3650 (
            .O(N__21936),
            .I(\b2v_inst5.N_2897_i ));
    Odrv4 I__3649 (
            .O(N__21933),
            .I(\b2v_inst5.N_2897_i ));
    InMux I__3648 (
            .O(N__21928),
            .I(N__21915));
    InMux I__3647 (
            .O(N__21927),
            .I(N__21915));
    InMux I__3646 (
            .O(N__21926),
            .I(N__21915));
    InMux I__3645 (
            .O(N__21925),
            .I(N__21915));
    InMux I__3644 (
            .O(N__21924),
            .I(N__21912));
    LocalMux I__3643 (
            .O(N__21915),
            .I(N__21909));
    LocalMux I__3642 (
            .O(N__21912),
            .I(\b2v_inst5.curr_stateZ0Z_0 ));
    Odrv4 I__3641 (
            .O(N__21909),
            .I(\b2v_inst5.curr_stateZ0Z_0 ));
    InMux I__3640 (
            .O(N__21904),
            .I(N__21889));
    InMux I__3639 (
            .O(N__21903),
            .I(N__21889));
    InMux I__3638 (
            .O(N__21902),
            .I(N__21889));
    InMux I__3637 (
            .O(N__21901),
            .I(N__21889));
    InMux I__3636 (
            .O(N__21900),
            .I(N__21889));
    LocalMux I__3635 (
            .O(N__21889),
            .I(\b2v_inst5.curr_state_RNIZ0Z_1 ));
    CascadeMux I__3634 (
            .O(N__21886),
            .I(\b2v_inst5.N_51_cascade_ ));
    InMux I__3633 (
            .O(N__21883),
            .I(N__21880));
    LocalMux I__3632 (
            .O(N__21880),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_0 ));
    CascadeMux I__3631 (
            .O(N__21877),
            .I(N__21871));
    InMux I__3630 (
            .O(N__21876),
            .I(N__21858));
    InMux I__3629 (
            .O(N__21875),
            .I(N__21858));
    InMux I__3628 (
            .O(N__21874),
            .I(N__21858));
    InMux I__3627 (
            .O(N__21871),
            .I(N__21858));
    InMux I__3626 (
            .O(N__21870),
            .I(N__21858));
    CascadeMux I__3625 (
            .O(N__21869),
            .I(N__21854));
    LocalMux I__3624 (
            .O(N__21858),
            .I(N__21850));
    InMux I__3623 (
            .O(N__21857),
            .I(N__21843));
    InMux I__3622 (
            .O(N__21854),
            .I(N__21843));
    InMux I__3621 (
            .O(N__21853),
            .I(N__21843));
    Span4Mux_v I__3620 (
            .O(N__21850),
            .I(N__21840));
    LocalMux I__3619 (
            .O(N__21843),
            .I(N__21837));
    Odrv4 I__3618 (
            .O(N__21840),
            .I(\b2v_inst11.N_19_i ));
    Odrv4 I__3617 (
            .O(N__21837),
            .I(\b2v_inst11.N_19_i ));
    CascadeMux I__3616 (
            .O(N__21832),
            .I(N__21829));
    InMux I__3615 (
            .O(N__21829),
            .I(N__21826));
    LocalMux I__3614 (
            .O(N__21826),
            .I(\b2v_inst11.N_5572_0 ));
    CascadeMux I__3613 (
            .O(N__21823),
            .I(N__21820));
    InMux I__3612 (
            .O(N__21820),
            .I(N__21814));
    InMux I__3611 (
            .O(N__21819),
            .I(N__21814));
    LocalMux I__3610 (
            .O(N__21814),
            .I(N__21809));
    InMux I__3609 (
            .O(N__21813),
            .I(N__21806));
    InMux I__3608 (
            .O(N__21812),
            .I(N__21803));
    Span4Mux_v I__3607 (
            .O(N__21809),
            .I(N__21798));
    LocalMux I__3606 (
            .O(N__21806),
            .I(N__21798));
    LocalMux I__3605 (
            .O(N__21803),
            .I(N__21795));
    Odrv4 I__3604 (
            .O(N__21798),
            .I(\b2v_inst11.N_172 ));
    Odrv4 I__3603 (
            .O(N__21795),
            .I(\b2v_inst11.N_172 ));
    InMux I__3602 (
            .O(N__21790),
            .I(N__21787));
    LocalMux I__3601 (
            .O(N__21787),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_1 ));
    InMux I__3600 (
            .O(N__21784),
            .I(N__21781));
    LocalMux I__3599 (
            .O(N__21781),
            .I(\b2v_inst11.dutycycle_eena ));
    InMux I__3598 (
            .O(N__21778),
            .I(N__21772));
    InMux I__3597 (
            .O(N__21777),
            .I(N__21772));
    LocalMux I__3596 (
            .O(N__21772),
            .I(\b2v_inst11.dutycycleZ1Z_0 ));
    CascadeMux I__3595 (
            .O(N__21769),
            .I(N__21766));
    InMux I__3594 (
            .O(N__21766),
            .I(N__21762));
    InMux I__3593 (
            .O(N__21765),
            .I(N__21759));
    LocalMux I__3592 (
            .O(N__21762),
            .I(\b2v_inst11.dutycycle_1_0_0 ));
    LocalMux I__3591 (
            .O(N__21759),
            .I(\b2v_inst11.dutycycle_1_0_0 ));
    CascadeMux I__3590 (
            .O(N__21754),
            .I(\b2v_inst11.dutycycle_eena_cascade_ ));
    InMux I__3589 (
            .O(N__21751),
            .I(N__21745));
    InMux I__3588 (
            .O(N__21750),
            .I(N__21745));
    LocalMux I__3587 (
            .O(N__21745),
            .I(\b2v_inst11.N_117_f0_1 ));
    CascadeMux I__3586 (
            .O(N__21742),
            .I(\b2v_inst11.dutycycle_eena_0_cascade_ ));
    CascadeMux I__3585 (
            .O(N__21739),
            .I(\b2v_inst11.dutycycle_cascade_ ));
    InMux I__3584 (
            .O(N__21736),
            .I(N__21730));
    InMux I__3583 (
            .O(N__21735),
            .I(N__21730));
    LocalMux I__3582 (
            .O(N__21730),
            .I(\b2v_inst11.dutycycle_1_0_1 ));
    InMux I__3581 (
            .O(N__21727),
            .I(N__21724));
    LocalMux I__3580 (
            .O(N__21724),
            .I(\b2v_inst11.dutycycle_eena_0 ));
    InMux I__3579 (
            .O(N__21721),
            .I(N__21715));
    InMux I__3578 (
            .O(N__21720),
            .I(N__21715));
    LocalMux I__3577 (
            .O(N__21715),
            .I(\b2v_inst11.dutycycleZ1Z_1 ));
    InMux I__3576 (
            .O(N__21712),
            .I(N__21706));
    InMux I__3575 (
            .O(N__21711),
            .I(N__21706));
    LocalMux I__3574 (
            .O(N__21706),
            .I(\b2v_inst11.dutycycle_0_6 ));
    CascadeMux I__3573 (
            .O(N__21703),
            .I(N__21700));
    InMux I__3572 (
            .O(N__21700),
            .I(N__21694));
    InMux I__3571 (
            .O(N__21699),
            .I(N__21694));
    LocalMux I__3570 (
            .O(N__21694),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQZ0Z6 ));
    InMux I__3569 (
            .O(N__21691),
            .I(N__21685));
    InMux I__3568 (
            .O(N__21690),
            .I(N__21685));
    LocalMux I__3567 (
            .O(N__21685),
            .I(N__21682));
    Span4Mux_h I__3566 (
            .O(N__21682),
            .I(N__21679));
    Odrv4 I__3565 (
            .O(N__21679),
            .I(\b2v_inst11.dutycycle_e_1_6 ));
    InMux I__3564 (
            .O(N__21676),
            .I(N__21673));
    LocalMux I__3563 (
            .O(N__21673),
            .I(N__21669));
    InMux I__3562 (
            .O(N__21672),
            .I(N__21666));
    Span4Mux_v I__3561 (
            .O(N__21669),
            .I(N__21662));
    LocalMux I__3560 (
            .O(N__21666),
            .I(N__21659));
    InMux I__3559 (
            .O(N__21665),
            .I(N__21656));
    Span4Mux_h I__3558 (
            .O(N__21662),
            .I(N__21651));
    Span4Mux_v I__3557 (
            .O(N__21659),
            .I(N__21651));
    LocalMux I__3556 (
            .O(N__21656),
            .I(\b2v_inst11.func_state_RNI_5Z0Z_1 ));
    Odrv4 I__3555 (
            .O(N__21651),
            .I(\b2v_inst11.func_state_RNI_5Z0Z_1 ));
    CascadeMux I__3554 (
            .O(N__21646),
            .I(\b2v_inst11.N_186_cascade_ ));
    InMux I__3553 (
            .O(N__21643),
            .I(N__21640));
    LocalMux I__3552 (
            .O(N__21640),
            .I(N__21637));
    Span4Mux_h I__3551 (
            .O(N__21637),
            .I(N__21634));
    Odrv4 I__3550 (
            .O(N__21634),
            .I(\b2v_inst11.N_426_0 ));
    CascadeMux I__3549 (
            .O(N__21631),
            .I(b2v_inst11_g0_i_m2_i_a6_1_1_cascade_));
    InMux I__3548 (
            .O(N__21628),
            .I(N__21625));
    LocalMux I__3547 (
            .O(N__21625),
            .I(N__21622));
    Span4Mux_h I__3546 (
            .O(N__21622),
            .I(N__21619));
    Span4Mux_v I__3545 (
            .O(N__21619),
            .I(N__21616));
    Odrv4 I__3544 (
            .O(N__21616),
            .I(SLP_S3n_ibuf_RNI9HQHZ0Z3));
    InMux I__3543 (
            .O(N__21613),
            .I(N__21607));
    InMux I__3542 (
            .O(N__21612),
            .I(N__21607));
    LocalMux I__3541 (
            .O(N__21607),
            .I(N__21604));
    Span4Mux_v I__3540 (
            .O(N__21604),
            .I(N__21599));
    InMux I__3539 (
            .O(N__21603),
            .I(N__21594));
    InMux I__3538 (
            .O(N__21602),
            .I(N__21594));
    Odrv4 I__3537 (
            .O(N__21599),
            .I(\b2v_inst11.dutycycle_RNI_9Z0Z_1 ));
    LocalMux I__3536 (
            .O(N__21594),
            .I(\b2v_inst11.dutycycle_RNI_9Z0Z_1 ));
    InMux I__3535 (
            .O(N__21589),
            .I(N__21586));
    LocalMux I__3534 (
            .O(N__21586),
            .I(\b2v_inst11.N_165_0 ));
    CascadeMux I__3533 (
            .O(N__21583),
            .I(\b2v_inst11.g0_i_m2_i_0_1_cascade_ ));
    InMux I__3532 (
            .O(N__21580),
            .I(N__21577));
    LocalMux I__3531 (
            .O(N__21577),
            .I(N_15_i_0_a4_1_0));
    InMux I__3530 (
            .O(N__21574),
            .I(\b2v_inst11.un1_dutycycle_94_cry_12 ));
    InMux I__3529 (
            .O(N__21571),
            .I(\b2v_inst11.un1_dutycycle_94_cry_13 ));
    InMux I__3528 (
            .O(N__21568),
            .I(\b2v_inst11.un1_dutycycle_94_cry_14 ));
    InMux I__3527 (
            .O(N__21565),
            .I(N__21562));
    LocalMux I__3526 (
            .O(N__21562),
            .I(N__21559));
    Odrv4 I__3525 (
            .O(N__21559),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ));
    InMux I__3524 (
            .O(N__21556),
            .I(N__21553));
    LocalMux I__3523 (
            .O(N__21553),
            .I(\b2v_inst11.dutycycle_RNIP7P13Z0Z_4 ));
    CascadeMux I__3522 (
            .O(N__21550),
            .I(N__21546));
    CascadeMux I__3521 (
            .O(N__21549),
            .I(N__21542));
    InMux I__3520 (
            .O(N__21546),
            .I(N__21537));
    InMux I__3519 (
            .O(N__21545),
            .I(N__21537));
    InMux I__3518 (
            .O(N__21542),
            .I(N__21534));
    LocalMux I__3517 (
            .O(N__21537),
            .I(\b2v_inst11.dutycycleZ1Z_4 ));
    LocalMux I__3516 (
            .O(N__21534),
            .I(\b2v_inst11.dutycycleZ1Z_4 ));
    CascadeMux I__3515 (
            .O(N__21529),
            .I(\b2v_inst11.dutycycle_RNIP7P13Z0Z_4_cascade_ ));
    CascadeMux I__3514 (
            .O(N__21526),
            .I(\b2v_inst11.dutycycleZ0Z_7_cascade_ ));
    InMux I__3513 (
            .O(N__21523),
            .I(N__21517));
    InMux I__3512 (
            .O(N__21522),
            .I(N__21517));
    LocalMux I__3511 (
            .O(N__21517),
            .I(\b2v_inst11.dutycycle_e_1_4 ));
    CascadeMux I__3510 (
            .O(N__21514),
            .I(\b2v_inst11.N_158_N_cascade_ ));
    InMux I__3509 (
            .O(N__21511),
            .I(\b2v_inst11.un1_dutycycle_94_cry_3 ));
    InMux I__3508 (
            .O(N__21508),
            .I(N__21505));
    LocalMux I__3507 (
            .O(N__21505),
            .I(N__21502));
    Odrv4 I__3506 (
            .O(N__21502),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19 ));
    InMux I__3505 (
            .O(N__21499),
            .I(\b2v_inst11.un1_dutycycle_94_cry_4_cZ0 ));
    InMux I__3504 (
            .O(N__21496),
            .I(N__21493));
    LocalMux I__3503 (
            .O(N__21493),
            .I(N__21490));
    Span4Mux_h I__3502 (
            .O(N__21490),
            .I(N__21487));
    Odrv4 I__3501 (
            .O(N__21487),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29 ));
    InMux I__3500 (
            .O(N__21484),
            .I(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__3499 (
            .O(N__21481),
            .I(N__21478));
    LocalMux I__3498 (
            .O(N__21478),
            .I(N__21475));
    Span4Mux_h I__3497 (
            .O(N__21475),
            .I(N__21472));
    Odrv4 I__3496 (
            .O(N__21472),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ));
    InMux I__3495 (
            .O(N__21469),
            .I(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ));
    InMux I__3494 (
            .O(N__21466),
            .I(bfn_6_10_0_));
    InMux I__3493 (
            .O(N__21463),
            .I(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ));
    InMux I__3492 (
            .O(N__21460),
            .I(\b2v_inst11.un1_dutycycle_94_cry_9 ));
    InMux I__3491 (
            .O(N__21457),
            .I(N__21451));
    InMux I__3490 (
            .O(N__21456),
            .I(N__21451));
    LocalMux I__3489 (
            .O(N__21451),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5 ));
    InMux I__3488 (
            .O(N__21448),
            .I(\b2v_inst11.un1_dutycycle_94_cry_10_cZ0 ));
    InMux I__3487 (
            .O(N__21445),
            .I(\b2v_inst11.un1_dutycycle_94_cry_11 ));
    CascadeMux I__3486 (
            .O(N__21442),
            .I(\b2v_inst11.un1_dutycycle_53_30_1_0_cascade_ ));
    CascadeMux I__3485 (
            .O(N__21439),
            .I(N__21436));
    InMux I__3484 (
            .O(N__21436),
            .I(N__21433));
    LocalMux I__3483 (
            .O(N__21433),
            .I(\b2v_inst11.dutycycle_RNI_2Z0Z_9 ));
    InMux I__3482 (
            .O(N__21430),
            .I(N__21427));
    LocalMux I__3481 (
            .O(N__21427),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_8 ));
    CascadeMux I__3480 (
            .O(N__21424),
            .I(\b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_ ));
    InMux I__3479 (
            .O(N__21421),
            .I(N__21414));
    InMux I__3478 (
            .O(N__21420),
            .I(N__21414));
    InMux I__3477 (
            .O(N__21419),
            .I(N__21410));
    LocalMux I__3476 (
            .O(N__21414),
            .I(N__21407));
    CascadeMux I__3475 (
            .O(N__21413),
            .I(N__21403));
    LocalMux I__3474 (
            .O(N__21410),
            .I(N__21399));
    Span4Mux_v I__3473 (
            .O(N__21407),
            .I(N__21396));
    InMux I__3472 (
            .O(N__21406),
            .I(N__21391));
    InMux I__3471 (
            .O(N__21403),
            .I(N__21391));
    InMux I__3470 (
            .O(N__21402),
            .I(N__21388));
    Odrv4 I__3469 (
            .O(N__21399),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ));
    Odrv4 I__3468 (
            .O(N__21396),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ));
    LocalMux I__3467 (
            .O(N__21391),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ));
    LocalMux I__3466 (
            .O(N__21388),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ));
    InMux I__3465 (
            .O(N__21379),
            .I(N__21375));
    InMux I__3464 (
            .O(N__21378),
            .I(N__21372));
    LocalMux I__3463 (
            .O(N__21375),
            .I(N__21369));
    LocalMux I__3462 (
            .O(N__21372),
            .I(N__21366));
    Odrv4 I__3461 (
            .O(N__21369),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_1 ));
    Odrv4 I__3460 (
            .O(N__21366),
            .I(\b2v_inst11.dutycycle_RNI_7Z0Z_1 ));
    InMux I__3459 (
            .O(N__21361),
            .I(N__21358));
    LocalMux I__3458 (
            .O(N__21358),
            .I(N__21355));
    Span4Mux_v I__3457 (
            .O(N__21355),
            .I(N__21352));
    Odrv4 I__3456 (
            .O(N__21352),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ));
    InMux I__3455 (
            .O(N__21349),
            .I(\b2v_inst11.un1_dutycycle_94_cry_0 ));
    InMux I__3454 (
            .O(N__21346),
            .I(\b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ));
    InMux I__3453 (
            .O(N__21343),
            .I(N__21340));
    LocalMux I__3452 (
            .O(N__21340),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ));
    InMux I__3451 (
            .O(N__21337),
            .I(\b2v_inst11.un1_dutycycle_94_cry_2 ));
    InMux I__3450 (
            .O(N__21334),
            .I(N__21331));
    LocalMux I__3449 (
            .O(N__21331),
            .I(\b2v_inst11.un2_count_clk_17_0_a2_1_3 ));
    CascadeMux I__3448 (
            .O(N__21328),
            .I(\b2v_inst11.un2_count_clk_17_0_a2_1_2_cascade_ ));
    InMux I__3447 (
            .O(N__21325),
            .I(N__21318));
    InMux I__3446 (
            .O(N__21324),
            .I(N__21318));
    CascadeMux I__3445 (
            .O(N__21323),
            .I(N__21315));
    LocalMux I__3444 (
            .O(N__21318),
            .I(N__21312));
    InMux I__3443 (
            .O(N__21315),
            .I(N__21309));
    Span4Mux_v I__3442 (
            .O(N__21312),
            .I(N__21304));
    LocalMux I__3441 (
            .O(N__21309),
            .I(N__21304));
    Odrv4 I__3440 (
            .O(N__21304),
            .I(\b2v_inst11.N_363 ));
    CascadeMux I__3439 (
            .O(N__21301),
            .I(N__21298));
    InMux I__3438 (
            .O(N__21298),
            .I(N__21294));
    InMux I__3437 (
            .O(N__21297),
            .I(N__21291));
    LocalMux I__3436 (
            .O(N__21294),
            .I(N__21288));
    LocalMux I__3435 (
            .O(N__21291),
            .I(\b2v_inst11.N_360 ));
    Odrv4 I__3434 (
            .O(N__21288),
            .I(\b2v_inst11.N_360 ));
    CascadeMux I__3433 (
            .O(N__21283),
            .I(\b2v_inst11.N_363_cascade_ ));
    InMux I__3432 (
            .O(N__21280),
            .I(N__21277));
    LocalMux I__3431 (
            .O(N__21277),
            .I(\b2v_inst11.N_365 ));
    CascadeMux I__3430 (
            .O(N__21274),
            .I(\b2v_inst11.N_365_cascade_ ));
    InMux I__3429 (
            .O(N__21271),
            .I(N__21268));
    LocalMux I__3428 (
            .O(N__21268),
            .I(N__21265));
    Odrv4 I__3427 (
            .O(N__21265),
            .I(\b2v_inst11.N_293 ));
    InMux I__3426 (
            .O(N__21262),
            .I(\b2v_inst11.mult1_un152_sum_cry_2_c ));
    InMux I__3425 (
            .O(N__21259),
            .I(\b2v_inst11.mult1_un152_sum_cry_3_c ));
    InMux I__3424 (
            .O(N__21256),
            .I(\b2v_inst11.mult1_un152_sum_cry_4_c ));
    InMux I__3423 (
            .O(N__21253),
            .I(\b2v_inst11.mult1_un152_sum_cry_5_c ));
    InMux I__3422 (
            .O(N__21250),
            .I(\b2v_inst11.mult1_un152_sum_cry_6_c ));
    InMux I__3421 (
            .O(N__21247),
            .I(\b2v_inst11.mult1_un152_sum_cry_7 ));
    CascadeMux I__3420 (
            .O(N__21244),
            .I(N__21239));
    CascadeMux I__3419 (
            .O(N__21243),
            .I(N__21236));
    CascadeMux I__3418 (
            .O(N__21242),
            .I(N__21233));
    InMux I__3417 (
            .O(N__21239),
            .I(N__21230));
    InMux I__3416 (
            .O(N__21236),
            .I(N__21225));
    InMux I__3415 (
            .O(N__21233),
            .I(N__21225));
    LocalMux I__3414 (
            .O(N__21230),
            .I(\b2v_inst11.mult1_un145_sum_i_0_8 ));
    LocalMux I__3413 (
            .O(N__21225),
            .I(\b2v_inst11.mult1_un145_sum_i_0_8 ));
    InMux I__3412 (
            .O(N__21220),
            .I(N__21217));
    LocalMux I__3411 (
            .O(N__21217),
            .I(N__21214));
    Span4Mux_v I__3410 (
            .O(N__21214),
            .I(N__21211));
    Span4Mux_v I__3409 (
            .O(N__21211),
            .I(N__21208));
    Span4Mux_h I__3408 (
            .O(N__21208),
            .I(N__21205));
    Odrv4 I__3407 (
            .O(N__21205),
            .I(VDDQ_OK_c));
    InMux I__3406 (
            .O(N__21202),
            .I(N__21196));
    InMux I__3405 (
            .O(N__21201),
            .I(N__21193));
    InMux I__3404 (
            .O(N__21200),
            .I(N__21190));
    InMux I__3403 (
            .O(N__21199),
            .I(N__21187));
    LocalMux I__3402 (
            .O(N__21196),
            .I(N__21184));
    LocalMux I__3401 (
            .O(N__21193),
            .I(N__21181));
    LocalMux I__3400 (
            .O(N__21190),
            .I(N__21178));
    LocalMux I__3399 (
            .O(N__21187),
            .I(N__21174));
    Span4Mux_v I__3398 (
            .O(N__21184),
            .I(N__21169));
    Span4Mux_v I__3397 (
            .O(N__21181),
            .I(N__21169));
    Span4Mux_v I__3396 (
            .O(N__21178),
            .I(N__21166));
    InMux I__3395 (
            .O(N__21177),
            .I(N__21161));
    Span4Mux_v I__3394 (
            .O(N__21174),
            .I(N__21154));
    Span4Mux_v I__3393 (
            .O(N__21169),
            .I(N__21154));
    Span4Mux_v I__3392 (
            .O(N__21166),
            .I(N__21154));
    InMux I__3391 (
            .O(N__21165),
            .I(N__21149));
    InMux I__3390 (
            .O(N__21164),
            .I(N__21149));
    LocalMux I__3389 (
            .O(N__21161),
            .I(VCCST_EN_i_0_o3_0));
    Odrv4 I__3388 (
            .O(N__21154),
            .I(VCCST_EN_i_0_o3_0));
    LocalMux I__3387 (
            .O(N__21149),
            .I(VCCST_EN_i_0_o3_0));
    InMux I__3386 (
            .O(N__21142),
            .I(N__21127));
    InMux I__3385 (
            .O(N__21141),
            .I(N__21127));
    InMux I__3384 (
            .O(N__21140),
            .I(N__21127));
    InMux I__3383 (
            .O(N__21139),
            .I(N__21127));
    InMux I__3382 (
            .O(N__21138),
            .I(N__21127));
    LocalMux I__3381 (
            .O(N__21127),
            .I(N__21124));
    Span12Mux_s6_v I__3380 (
            .O(N__21124),
            .I(N__21121));
    Odrv12 I__3379 (
            .O(N__21121),
            .I(\b2v_inst16.N_208_0 ));
    CascadeMux I__3378 (
            .O(N__21118),
            .I(N__21115));
    InMux I__3377 (
            .O(N__21115),
            .I(N__21112));
    LocalMux I__3376 (
            .O(N__21112),
            .I(N__21109));
    Span4Mux_v I__3375 (
            .O(N__21109),
            .I(N__21105));
    InMux I__3374 (
            .O(N__21108),
            .I(N__21102));
    Odrv4 I__3373 (
            .O(N__21105),
            .I(\b2v_inst11.N_354 ));
    LocalMux I__3372 (
            .O(N__21102),
            .I(\b2v_inst11.N_354 ));
    InMux I__3371 (
            .O(N__21097),
            .I(N__21091));
    InMux I__3370 (
            .O(N__21096),
            .I(N__21091));
    LocalMux I__3369 (
            .O(N__21091),
            .I(\b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29 ));
    CascadeMux I__3368 (
            .O(N__21088),
            .I(N__21085));
    InMux I__3367 (
            .O(N__21085),
            .I(N__21082));
    LocalMux I__3366 (
            .O(N__21082),
            .I(\b2v_inst200.count_3_11 ));
    InMux I__3365 (
            .O(N__21079),
            .I(N__21076));
    LocalMux I__3364 (
            .O(N__21076),
            .I(\b2v_inst200.countZ0Z_11 ));
    InMux I__3363 (
            .O(N__21073),
            .I(N__21069));
    InMux I__3362 (
            .O(N__21072),
            .I(N__21066));
    LocalMux I__3361 (
            .O(N__21069),
            .I(\b2v_inst200.countZ0Z_17 ));
    LocalMux I__3360 (
            .O(N__21066),
            .I(\b2v_inst200.countZ0Z_17 ));
    CascadeMux I__3359 (
            .O(N__21061),
            .I(\b2v_inst200.countZ0Z_11_cascade_ ));
    InMux I__3358 (
            .O(N__21058),
            .I(N__21054));
    InMux I__3357 (
            .O(N__21057),
            .I(N__21051));
    LocalMux I__3356 (
            .O(N__21054),
            .I(\b2v_inst200.countZ0Z_16 ));
    LocalMux I__3355 (
            .O(N__21051),
            .I(\b2v_inst200.countZ0Z_16 ));
    InMux I__3354 (
            .O(N__21046),
            .I(N__21043));
    LocalMux I__3353 (
            .O(N__21043),
            .I(N__21040));
    Odrv4 I__3352 (
            .O(N__21040),
            .I(\b2v_inst200.un25_clk_100khz_9 ));
    InMux I__3351 (
            .O(N__21037),
            .I(N__21034));
    LocalMux I__3350 (
            .O(N__21034),
            .I(N__21031));
    Span4Mux_h I__3349 (
            .O(N__21031),
            .I(N__21028));
    Odrv4 I__3348 (
            .O(N__21028),
            .I(\b2v_inst200.un25_clk_100khz_12 ));
    CascadeMux I__3347 (
            .O(N__21025),
            .I(\b2v_inst200.un25_clk_100khz_13_cascade_ ));
    InMux I__3346 (
            .O(N__21022),
            .I(N__21019));
    LocalMux I__3345 (
            .O(N__21019),
            .I(\b2v_inst200.un25_clk_100khz_14 ));
    CascadeMux I__3344 (
            .O(N__21016),
            .I(\b2v_inst200.count_RNIC03N_6Z0Z_0_cascade_ ));
    InMux I__3343 (
            .O(N__21013),
            .I(N__21007));
    InMux I__3342 (
            .O(N__21012),
            .I(N__21007));
    LocalMux I__3341 (
            .O(N__21007),
            .I(\b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0 ));
    InMux I__3340 (
            .O(N__21004),
            .I(N__21001));
    LocalMux I__3339 (
            .O(N__21001),
            .I(\b2v_inst200.count_3_10 ));
    CascadeMux I__3338 (
            .O(N__20998),
            .I(\b2v_inst200.count_RNI_0_0_cascade_ ));
    CascadeMux I__3337 (
            .O(N__20995),
            .I(N__20991));
    InMux I__3336 (
            .O(N__20994),
            .I(N__20988));
    InMux I__3335 (
            .O(N__20991),
            .I(N__20985));
    LocalMux I__3334 (
            .O(N__20988),
            .I(\b2v_inst200.countZ0Z_10 ));
    LocalMux I__3333 (
            .O(N__20985),
            .I(\b2v_inst200.countZ0Z_10 ));
    InMux I__3332 (
            .O(N__20980),
            .I(N__20977));
    LocalMux I__3331 (
            .O(N__20977),
            .I(N__20974));
    Span4Mux_h I__3330 (
            .O(N__20974),
            .I(N__20970));
    InMux I__3329 (
            .O(N__20973),
            .I(N__20967));
    Odrv4 I__3328 (
            .O(N__20970),
            .I(\b2v_inst16.count_rst_1 ));
    LocalMux I__3327 (
            .O(N__20967),
            .I(\b2v_inst16.count_rst_1 ));
    InMux I__3326 (
            .O(N__20962),
            .I(N__20959));
    LocalMux I__3325 (
            .O(N__20959),
            .I(N__20956));
    Span4Mux_s3_h I__3324 (
            .O(N__20956),
            .I(N__20953));
    Odrv4 I__3323 (
            .O(N__20953),
            .I(\b2v_inst16.count_4_12 ));
    CEMux I__3322 (
            .O(N__20950),
            .I(N__20946));
    CEMux I__3321 (
            .O(N__20949),
            .I(N__20929));
    LocalMux I__3320 (
            .O(N__20946),
            .I(N__20925));
    CEMux I__3319 (
            .O(N__20945),
            .I(N__20922));
    CEMux I__3318 (
            .O(N__20944),
            .I(N__20919));
    CEMux I__3317 (
            .O(N__20943),
            .I(N__20916));
    CEMux I__3316 (
            .O(N__20942),
            .I(N__20907));
    InMux I__3315 (
            .O(N__20941),
            .I(N__20902));
    InMux I__3314 (
            .O(N__20940),
            .I(N__20902));
    InMux I__3313 (
            .O(N__20939),
            .I(N__20897));
    InMux I__3312 (
            .O(N__20938),
            .I(N__20897));
    InMux I__3311 (
            .O(N__20937),
            .I(N__20890));
    InMux I__3310 (
            .O(N__20936),
            .I(N__20890));
    InMux I__3309 (
            .O(N__20935),
            .I(N__20890));
    InMux I__3308 (
            .O(N__20934),
            .I(N__20883));
    InMux I__3307 (
            .O(N__20933),
            .I(N__20883));
    InMux I__3306 (
            .O(N__20932),
            .I(N__20883));
    LocalMux I__3305 (
            .O(N__20929),
            .I(N__20879));
    CEMux I__3304 (
            .O(N__20928),
            .I(N__20876));
    Span4Mux_v I__3303 (
            .O(N__20925),
            .I(N__20873));
    LocalMux I__3302 (
            .O(N__20922),
            .I(N__20870));
    LocalMux I__3301 (
            .O(N__20919),
            .I(N__20867));
    LocalMux I__3300 (
            .O(N__20916),
            .I(N__20864));
    InMux I__3299 (
            .O(N__20915),
            .I(N__20859));
    CEMux I__3298 (
            .O(N__20914),
            .I(N__20859));
    InMux I__3297 (
            .O(N__20913),
            .I(N__20856));
    InMux I__3296 (
            .O(N__20912),
            .I(N__20849));
    InMux I__3295 (
            .O(N__20911),
            .I(N__20849));
    InMux I__3294 (
            .O(N__20910),
            .I(N__20849));
    LocalMux I__3293 (
            .O(N__20907),
            .I(N__20838));
    LocalMux I__3292 (
            .O(N__20902),
            .I(N__20838));
    LocalMux I__3291 (
            .O(N__20897),
            .I(N__20838));
    LocalMux I__3290 (
            .O(N__20890),
            .I(N__20838));
    LocalMux I__3289 (
            .O(N__20883),
            .I(N__20838));
    InMux I__3288 (
            .O(N__20882),
            .I(N__20835));
    Span4Mux_s1_v I__3287 (
            .O(N__20879),
            .I(N__20832));
    LocalMux I__3286 (
            .O(N__20876),
            .I(N__20829));
    Span4Mux_h I__3285 (
            .O(N__20873),
            .I(N__20820));
    Span4Mux_v I__3284 (
            .O(N__20870),
            .I(N__20820));
    Span4Mux_v I__3283 (
            .O(N__20867),
            .I(N__20820));
    Span4Mux_s1_h I__3282 (
            .O(N__20864),
            .I(N__20820));
    LocalMux I__3281 (
            .O(N__20859),
            .I(N__20809));
    LocalMux I__3280 (
            .O(N__20856),
            .I(N__20809));
    LocalMux I__3279 (
            .O(N__20849),
            .I(N__20809));
    Span4Mux_s1_v I__3278 (
            .O(N__20838),
            .I(N__20809));
    LocalMux I__3277 (
            .O(N__20835),
            .I(N__20809));
    Odrv4 I__3276 (
            .O(N__20832),
            .I(\b2v_inst16.count_en ));
    Odrv12 I__3275 (
            .O(N__20829),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__3274 (
            .O(N__20820),
            .I(\b2v_inst16.count_en ));
    Odrv4 I__3273 (
            .O(N__20809),
            .I(\b2v_inst16.count_en ));
    SRMux I__3272 (
            .O(N__20800),
            .I(N__20793));
    SRMux I__3271 (
            .O(N__20799),
            .I(N__20790));
    SRMux I__3270 (
            .O(N__20798),
            .I(N__20786));
    SRMux I__3269 (
            .O(N__20797),
            .I(N__20782));
    SRMux I__3268 (
            .O(N__20796),
            .I(N__20779));
    LocalMux I__3267 (
            .O(N__20793),
            .I(N__20776));
    LocalMux I__3266 (
            .O(N__20790),
            .I(N__20773));
    SRMux I__3265 (
            .O(N__20789),
            .I(N__20770));
    LocalMux I__3264 (
            .O(N__20786),
            .I(N__20767));
    SRMux I__3263 (
            .O(N__20785),
            .I(N__20764));
    LocalMux I__3262 (
            .O(N__20782),
            .I(N__20760));
    LocalMux I__3261 (
            .O(N__20779),
            .I(N__20757));
    Span4Mux_h I__3260 (
            .O(N__20776),
            .I(N__20750));
    Span4Mux_s3_v I__3259 (
            .O(N__20773),
            .I(N__20750));
    LocalMux I__3258 (
            .O(N__20770),
            .I(N__20750));
    Span4Mux_h I__3257 (
            .O(N__20767),
            .I(N__20745));
    LocalMux I__3256 (
            .O(N__20764),
            .I(N__20745));
    SRMux I__3255 (
            .O(N__20763),
            .I(N__20742));
    Span4Mux_s2_v I__3254 (
            .O(N__20760),
            .I(N__20739));
    Span4Mux_h I__3253 (
            .O(N__20757),
            .I(N__20736));
    Span4Mux_h I__3252 (
            .O(N__20750),
            .I(N__20733));
    Span4Mux_v I__3251 (
            .O(N__20745),
            .I(N__20728));
    LocalMux I__3250 (
            .O(N__20742),
            .I(N__20728));
    Span4Mux_h I__3249 (
            .O(N__20739),
            .I(N__20725));
    Span4Mux_s0_h I__3248 (
            .O(N__20736),
            .I(N__20722));
    Span4Mux_s0_h I__3247 (
            .O(N__20733),
            .I(N__20719));
    Span4Mux_h I__3246 (
            .O(N__20728),
            .I(N__20716));
    Odrv4 I__3245 (
            .O(N__20725),
            .I(\b2v_inst16.N_2987_i ));
    Odrv4 I__3244 (
            .O(N__20722),
            .I(\b2v_inst16.N_2987_i ));
    Odrv4 I__3243 (
            .O(N__20719),
            .I(\b2v_inst16.N_2987_i ));
    Odrv4 I__3242 (
            .O(N__20716),
            .I(\b2v_inst16.N_2987_i ));
    InMux I__3241 (
            .O(N__20707),
            .I(N__20703));
    InMux I__3240 (
            .O(N__20706),
            .I(N__20700));
    LocalMux I__3239 (
            .O(N__20703),
            .I(N__20688));
    LocalMux I__3238 (
            .O(N__20700),
            .I(N__20688));
    InMux I__3237 (
            .O(N__20699),
            .I(N__20685));
    InMux I__3236 (
            .O(N__20698),
            .I(N__20682));
    InMux I__3235 (
            .O(N__20697),
            .I(N__20675));
    InMux I__3234 (
            .O(N__20696),
            .I(N__20675));
    InMux I__3233 (
            .O(N__20695),
            .I(N__20675));
    InMux I__3232 (
            .O(N__20694),
            .I(N__20670));
    InMux I__3231 (
            .O(N__20693),
            .I(N__20670));
    Span4Mux_v I__3230 (
            .O(N__20688),
            .I(N__20659));
    LocalMux I__3229 (
            .O(N__20685),
            .I(N__20659));
    LocalMux I__3228 (
            .O(N__20682),
            .I(N__20659));
    LocalMux I__3227 (
            .O(N__20675),
            .I(N__20659));
    LocalMux I__3226 (
            .O(N__20670),
            .I(N__20659));
    Span4Mux_v I__3225 (
            .O(N__20659),
            .I(N__20656));
    Odrv4 I__3224 (
            .O(N__20656),
            .I(\b2v_inst11.N_366 ));
    InMux I__3223 (
            .O(N__20653),
            .I(N__20650));
    LocalMux I__3222 (
            .O(N__20650),
            .I(N__20647));
    Odrv4 I__3221 (
            .O(N__20647),
            .I(\b2v_inst200.count_3_13 ));
    InMux I__3220 (
            .O(N__20644),
            .I(N__20640));
    InMux I__3219 (
            .O(N__20643),
            .I(N__20637));
    LocalMux I__3218 (
            .O(N__20640),
            .I(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ));
    LocalMux I__3217 (
            .O(N__20637),
            .I(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ));
    InMux I__3216 (
            .O(N__20632),
            .I(N__20629));
    LocalMux I__3215 (
            .O(N__20629),
            .I(\b2v_inst200.countZ0Z_13 ));
    CascadeMux I__3214 (
            .O(N__20626),
            .I(\b2v_inst200.countZ0Z_13_cascade_ ));
    InMux I__3213 (
            .O(N__20623),
            .I(N__20619));
    InMux I__3212 (
            .O(N__20622),
            .I(N__20616));
    LocalMux I__3211 (
            .O(N__20619),
            .I(\b2v_inst200.countZ0Z_0 ));
    LocalMux I__3210 (
            .O(N__20616),
            .I(\b2v_inst200.countZ0Z_0 ));
    InMux I__3209 (
            .O(N__20611),
            .I(N__20607));
    InMux I__3208 (
            .O(N__20610),
            .I(N__20604));
    LocalMux I__3207 (
            .O(N__20607),
            .I(N__20601));
    LocalMux I__3206 (
            .O(N__20604),
            .I(N__20598));
    Span4Mux_h I__3205 (
            .O(N__20601),
            .I(N__20593));
    Span4Mux_s1_v I__3204 (
            .O(N__20598),
            .I(N__20593));
    Odrv4 I__3203 (
            .O(N__20593),
            .I(\b2v_inst200.countZ0Z_7 ));
    InMux I__3202 (
            .O(N__20590),
            .I(N__20586));
    InMux I__3201 (
            .O(N__20589),
            .I(N__20583));
    LocalMux I__3200 (
            .O(N__20586),
            .I(N__20578));
    LocalMux I__3199 (
            .O(N__20583),
            .I(N__20578));
    Span4Mux_s1_v I__3198 (
            .O(N__20578),
            .I(N__20575));
    Odrv4 I__3197 (
            .O(N__20575),
            .I(\b2v_inst200.countZ0Z_5 ));
    CascadeMux I__3196 (
            .O(N__20572),
            .I(\b2v_inst200.un25_clk_100khz_10_cascade_ ));
    InMux I__3195 (
            .O(N__20569),
            .I(N__20566));
    LocalMux I__3194 (
            .O(N__20566),
            .I(\b2v_inst200.un25_clk_100khz_3 ));
    InMux I__3193 (
            .O(N__20563),
            .I(N__20559));
    InMux I__3192 (
            .O(N__20562),
            .I(N__20556));
    LocalMux I__3191 (
            .O(N__20559),
            .I(\b2v_inst200.countZ0Z_15 ));
    LocalMux I__3190 (
            .O(N__20556),
            .I(\b2v_inst200.countZ0Z_15 ));
    InMux I__3189 (
            .O(N__20551),
            .I(N__20545));
    InMux I__3188 (
            .O(N__20550),
            .I(N__20545));
    LocalMux I__3187 (
            .O(N__20545),
            .I(\b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ));
    InMux I__3186 (
            .O(N__20542),
            .I(N__20539));
    LocalMux I__3185 (
            .O(N__20539),
            .I(\b2v_inst200.count_3_15 ));
    InMux I__3184 (
            .O(N__20536),
            .I(N__20530));
    InMux I__3183 (
            .O(N__20535),
            .I(N__20530));
    LocalMux I__3182 (
            .O(N__20530),
            .I(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ));
    InMux I__3181 (
            .O(N__20527),
            .I(N__20524));
    LocalMux I__3180 (
            .O(N__20524),
            .I(\b2v_inst200.count_3_14 ));
    InMux I__3179 (
            .O(N__20521),
            .I(N__20517));
    InMux I__3178 (
            .O(N__20520),
            .I(N__20514));
    LocalMux I__3177 (
            .O(N__20517),
            .I(\b2v_inst200.countZ0Z_14 ));
    LocalMux I__3176 (
            .O(N__20514),
            .I(\b2v_inst200.countZ0Z_14 ));
    InMux I__3175 (
            .O(N__20509),
            .I(N__20506));
    LocalMux I__3174 (
            .O(N__20506),
            .I(N__20503));
    Span4Mux_v I__3173 (
            .O(N__20503),
            .I(N__20500));
    Odrv4 I__3172 (
            .O(N__20500),
            .I(\b2v_inst200.count_0_16 ));
    InMux I__3171 (
            .O(N__20497),
            .I(N__20493));
    CascadeMux I__3170 (
            .O(N__20496),
            .I(N__20490));
    LocalMux I__3169 (
            .O(N__20493),
            .I(N__20487));
    InMux I__3168 (
            .O(N__20490),
            .I(N__20484));
    Odrv4 I__3167 (
            .O(N__20487),
            .I(\b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79 ));
    LocalMux I__3166 (
            .O(N__20484),
            .I(\b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79 ));
    InMux I__3165 (
            .O(N__20479),
            .I(N__20476));
    LocalMux I__3164 (
            .O(N__20476),
            .I(\b2v_inst200.countZ0Z_6 ));
    CascadeMux I__3163 (
            .O(N__20473),
            .I(\b2v_inst200.countZ0Z_6_cascade_ ));
    InMux I__3162 (
            .O(N__20470),
            .I(N__20466));
    InMux I__3161 (
            .O(N__20469),
            .I(N__20463));
    LocalMux I__3160 (
            .O(N__20466),
            .I(\b2v_inst200.countZ0Z_8 ));
    LocalMux I__3159 (
            .O(N__20463),
            .I(\b2v_inst200.countZ0Z_8 ));
    InMux I__3158 (
            .O(N__20458),
            .I(N__20452));
    InMux I__3157 (
            .O(N__20457),
            .I(N__20452));
    LocalMux I__3156 (
            .O(N__20452),
            .I(\b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ));
    CascadeMux I__3155 (
            .O(N__20449),
            .I(N__20446));
    InMux I__3154 (
            .O(N__20446),
            .I(N__20443));
    LocalMux I__3153 (
            .O(N__20443),
            .I(\b2v_inst200.count_3_6 ));
    InMux I__3152 (
            .O(N__20440),
            .I(N__20434));
    InMux I__3151 (
            .O(N__20439),
            .I(N__20434));
    LocalMux I__3150 (
            .O(N__20434),
            .I(\b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0 ));
    InMux I__3149 (
            .O(N__20431),
            .I(N__20428));
    LocalMux I__3148 (
            .O(N__20428),
            .I(\b2v_inst200.count_3_8 ));
    InMux I__3147 (
            .O(N__20425),
            .I(N__20422));
    LocalMux I__3146 (
            .O(N__20422),
            .I(\b2v_inst200.count_1_0 ));
    CascadeMux I__3145 (
            .O(N__20419),
            .I(\b2v_inst200.countZ0Z_0_cascade_ ));
    InMux I__3144 (
            .O(N__20416),
            .I(N__20413));
    LocalMux I__3143 (
            .O(N__20413),
            .I(\b2v_inst200.count_3_0 ));
    InMux I__3142 (
            .O(N__20410),
            .I(N__20406));
    InMux I__3141 (
            .O(N__20409),
            .I(N__20403));
    LocalMux I__3140 (
            .O(N__20406),
            .I(N__20400));
    LocalMux I__3139 (
            .O(N__20403),
            .I(N__20397));
    Odrv12 I__3138 (
            .O(N__20400),
            .I(\b2v_inst200.countZ0Z_12 ));
    Odrv4 I__3137 (
            .O(N__20397),
            .I(\b2v_inst200.countZ0Z_12 ));
    InMux I__3136 (
            .O(N__20392),
            .I(N__20389));
    LocalMux I__3135 (
            .O(N__20389),
            .I(N__20385));
    InMux I__3134 (
            .O(N__20388),
            .I(N__20382));
    Span4Mux_h I__3133 (
            .O(N__20385),
            .I(N__20379));
    LocalMux I__3132 (
            .O(N__20382),
            .I(\b2v_inst20.counterZ0Z_7 ));
    Odrv4 I__3131 (
            .O(N__20379),
            .I(\b2v_inst20.counterZ0Z_7 ));
    InMux I__3130 (
            .O(N__20374),
            .I(N__20371));
    LocalMux I__3129 (
            .O(N__20371),
            .I(N__20367));
    InMux I__3128 (
            .O(N__20370),
            .I(N__20363));
    Span4Mux_v I__3127 (
            .O(N__20367),
            .I(N__20360));
    InMux I__3126 (
            .O(N__20366),
            .I(N__20357));
    LocalMux I__3125 (
            .O(N__20363),
            .I(\b2v_inst20.counterZ0Z_5 ));
    Odrv4 I__3124 (
            .O(N__20360),
            .I(\b2v_inst20.counterZ0Z_5 ));
    LocalMux I__3123 (
            .O(N__20357),
            .I(\b2v_inst20.counterZ0Z_5 ));
    InMux I__3122 (
            .O(N__20350),
            .I(N__20347));
    LocalMux I__3121 (
            .O(N__20347),
            .I(N__20343));
    CascadeMux I__3120 (
            .O(N__20346),
            .I(N__20339));
    Span4Mux_h I__3119 (
            .O(N__20343),
            .I(N__20336));
    InMux I__3118 (
            .O(N__20342),
            .I(N__20331));
    InMux I__3117 (
            .O(N__20339),
            .I(N__20331));
    Odrv4 I__3116 (
            .O(N__20336),
            .I(\b2v_inst20.counterZ0Z_6 ));
    LocalMux I__3115 (
            .O(N__20331),
            .I(\b2v_inst20.counterZ0Z_6 ));
    InMux I__3114 (
            .O(N__20326),
            .I(N__20323));
    LocalMux I__3113 (
            .O(N__20323),
            .I(N__20319));
    InMux I__3112 (
            .O(N__20322),
            .I(N__20315));
    Span4Mux_s3_h I__3111 (
            .O(N__20319),
            .I(N__20312));
    InMux I__3110 (
            .O(N__20318),
            .I(N__20309));
    LocalMux I__3109 (
            .O(N__20315),
            .I(\b2v_inst20.counterZ0Z_1 ));
    Odrv4 I__3108 (
            .O(N__20312),
            .I(\b2v_inst20.counterZ0Z_1 ));
    LocalMux I__3107 (
            .O(N__20309),
            .I(\b2v_inst20.counterZ0Z_1 ));
    InMux I__3106 (
            .O(N__20302),
            .I(N__20299));
    LocalMux I__3105 (
            .O(N__20299),
            .I(N__20296));
    Odrv4 I__3104 (
            .O(N__20296),
            .I(\b2v_inst20.un4_counter_1_and ));
    InMux I__3103 (
            .O(N__20293),
            .I(N__20290));
    LocalMux I__3102 (
            .O(N__20290),
            .I(N__20284));
    InMux I__3101 (
            .O(N__20289),
            .I(N__20281));
    InMux I__3100 (
            .O(N__20288),
            .I(N__20278));
    CascadeMux I__3099 (
            .O(N__20287),
            .I(N__20273));
    Span4Mux_v I__3098 (
            .O(N__20284),
            .I(N__20270));
    LocalMux I__3097 (
            .O(N__20281),
            .I(N__20267));
    LocalMux I__3096 (
            .O(N__20278),
            .I(N__20264));
    InMux I__3095 (
            .O(N__20277),
            .I(N__20261));
    CascadeMux I__3094 (
            .O(N__20276),
            .I(N__20256));
    InMux I__3093 (
            .O(N__20273),
            .I(N__20253));
    Span4Mux_h I__3092 (
            .O(N__20270),
            .I(N__20248));
    Span4Mux_h I__3091 (
            .O(N__20267),
            .I(N__20248));
    Span12Mux_s7_h I__3090 (
            .O(N__20264),
            .I(N__20243));
    LocalMux I__3089 (
            .O(N__20261),
            .I(N__20243));
    InMux I__3088 (
            .O(N__20260),
            .I(N__20236));
    InMux I__3087 (
            .O(N__20259),
            .I(N__20236));
    InMux I__3086 (
            .O(N__20256),
            .I(N__20236));
    LocalMux I__3085 (
            .O(N__20253),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    Odrv4 I__3084 (
            .O(N__20248),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    Odrv12 I__3083 (
            .O(N__20243),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    LocalMux I__3082 (
            .O(N__20236),
            .I(SYNTHESIZED_WIRE_1keep_3_fast));
    IoInMux I__3081 (
            .O(N__20227),
            .I(N__20224));
    LocalMux I__3080 (
            .O(N__20224),
            .I(N__20221));
    Span12Mux_s4_h I__3079 (
            .O(N__20221),
            .I(N__20218));
    Odrv12 I__3078 (
            .O(N__20218),
            .I(HDA_SDO_ATP_c));
    InMux I__3077 (
            .O(N__20215),
            .I(N__20212));
    LocalMux I__3076 (
            .O(N__20212),
            .I(\b2v_inst200.N_205 ));
    CascadeMux I__3075 (
            .O(N__20209),
            .I(\b2v_inst200.N_205_cascade_ ));
    CascadeMux I__3074 (
            .O(N__20206),
            .I(G_2734_cascade_));
    InMux I__3073 (
            .O(N__20203),
            .I(N__20197));
    InMux I__3072 (
            .O(N__20202),
            .I(N__20197));
    LocalMux I__3071 (
            .O(N__20197),
            .I(\b2v_inst200.curr_stateZ0Z_2 ));
    CascadeMux I__3070 (
            .O(N__20194),
            .I(\b2v_inst200.curr_stateZ0Z_2_cascade_ ));
    CascadeMux I__3069 (
            .O(N__20191),
            .I(N__20188));
    InMux I__3068 (
            .O(N__20188),
            .I(N__20185));
    LocalMux I__3067 (
            .O(N__20185),
            .I(\b2v_inst200.HDA_SDO_ATP_0 ));
    InMux I__3066 (
            .O(N__20182),
            .I(N__20179));
    LocalMux I__3065 (
            .O(N__20179),
            .I(G_2734));
    InMux I__3064 (
            .O(N__20176),
            .I(N__20173));
    LocalMux I__3063 (
            .O(N__20173),
            .I(\b2v_inst200.curr_state_0_2 ));
    CascadeMux I__3062 (
            .O(N__20170),
            .I(N_73_mux_i_i_a7_4_0_cascade_));
    CascadeMux I__3061 (
            .O(N__20167),
            .I(N__20164));
    InMux I__3060 (
            .O(N__20164),
            .I(N__20161));
    LocalMux I__3059 (
            .O(N__20161),
            .I(\b2v_inst11.N_73_mux_i_i_1 ));
    InMux I__3058 (
            .O(N__20158),
            .I(N__20154));
    InMux I__3057 (
            .O(N__20157),
            .I(N__20151));
    LocalMux I__3056 (
            .O(N__20154),
            .I(\b2v_inst11.N_73_mux_i_i_2 ));
    LocalMux I__3055 (
            .O(N__20151),
            .I(\b2v_inst11.N_73_mux_i_i_2 ));
    InMux I__3054 (
            .O(N__20146),
            .I(N__20142));
    InMux I__3053 (
            .O(N__20145),
            .I(N__20139));
    LocalMux I__3052 (
            .O(N__20142),
            .I(N__20134));
    LocalMux I__3051 (
            .O(N__20139),
            .I(N__20134));
    Span4Mux_v I__3050 (
            .O(N__20134),
            .I(N__20131));
    Odrv4 I__3049 (
            .O(N__20131),
            .I(N_15));
    CascadeMux I__3048 (
            .O(N__20128),
            .I(\b2v_inst11.N_73_mux_i_i_1_cascade_ ));
    InMux I__3047 (
            .O(N__20125),
            .I(N__20113));
    InMux I__3046 (
            .O(N__20124),
            .I(N__20113));
    InMux I__3045 (
            .O(N__20123),
            .I(N__20113));
    InMux I__3044 (
            .O(N__20122),
            .I(N__20113));
    LocalMux I__3043 (
            .O(N__20113),
            .I(\b2v_inst11.dutycycle_0_5 ));
    InMux I__3042 (
            .O(N__20110),
            .I(N__20107));
    LocalMux I__3041 (
            .O(N__20107),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx ));
    CascadeMux I__3040 (
            .O(N__20104),
            .I(RSMRSTn_fast_RNIGMH81_cascade_));
    CascadeMux I__3039 (
            .O(N__20101),
            .I(N__20098));
    InMux I__3038 (
            .O(N__20098),
            .I(N__20095));
    LocalMux I__3037 (
            .O(N__20095),
            .I(N__20091));
    InMux I__3036 (
            .O(N__20094),
            .I(N__20088));
    Odrv12 I__3035 (
            .O(N__20091),
            .I(N_7_2));
    LocalMux I__3034 (
            .O(N__20088),
            .I(N_7_2));
    InMux I__3033 (
            .O(N__20083),
            .I(N__20078));
    InMux I__3032 (
            .O(N__20082),
            .I(N__20073));
    InMux I__3031 (
            .O(N__20081),
            .I(N__20073));
    LocalMux I__3030 (
            .O(N__20078),
            .I(N__20070));
    LocalMux I__3029 (
            .O(N__20073),
            .I(N_10_0));
    Odrv4 I__3028 (
            .O(N__20070),
            .I(N_10_0));
    InMux I__3027 (
            .O(N__20065),
            .I(N__20062));
    LocalMux I__3026 (
            .O(N__20062),
            .I(\b2v_inst20.tmp_1_rep1_RNI07FZ0Z73 ));
    InMux I__3025 (
            .O(N__20059),
            .I(N__20056));
    LocalMux I__3024 (
            .O(N__20056),
            .I(N__20053));
    Span4Mux_h I__3023 (
            .O(N__20053),
            .I(N__20050));
    Span4Mux_h I__3022 (
            .O(N__20050),
            .I(N__20047));
    Odrv4 I__3021 (
            .O(N__20047),
            .I(\b2v_inst20.counter_1_cry_5_THRU_CO ));
    CascadeMux I__3020 (
            .O(N__20044),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_5_cascade_ ));
    CascadeMux I__3019 (
            .O(N__20041),
            .I(N__20035));
    InMux I__3018 (
            .O(N__20040),
            .I(N__20028));
    InMux I__3017 (
            .O(N__20039),
            .I(N__20028));
    InMux I__3016 (
            .O(N__20038),
            .I(N__20028));
    InMux I__3015 (
            .O(N__20035),
            .I(N__20025));
    LocalMux I__3014 (
            .O(N__20028),
            .I(N__20022));
    LocalMux I__3013 (
            .O(N__20025),
            .I(N__20016));
    Span4Mux_h I__3012 (
            .O(N__20022),
            .I(N__20016));
    InMux I__3011 (
            .O(N__20021),
            .I(N__20013));
    Odrv4 I__3010 (
            .O(N__20016),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_1 ));
    LocalMux I__3009 (
            .O(N__20013),
            .I(\b2v_inst11.dutycycle_RNI_3Z0Z_1 ));
    CascadeMux I__3008 (
            .O(N__20008),
            .I(\b2v_inst11.N_73_mux_i_i_o7_1_cascade_ ));
    InMux I__3007 (
            .O(N__20005),
            .I(N__20002));
    LocalMux I__3006 (
            .O(N__20002),
            .I(\b2v_inst11.dutycycle_RNIUNGA5Z0Z_5 ));
    InMux I__3005 (
            .O(N__19999),
            .I(N__19996));
    LocalMux I__3004 (
            .O(N__19996),
            .I(\b2v_inst11.N_73_mux_i_i_0 ));
    CascadeMux I__3003 (
            .O(N__19993),
            .I(\b2v_inst11.N_73_mux_i_i_a7_1_cascade_ ));
    InMux I__3002 (
            .O(N__19990),
            .I(N__19983));
    InMux I__3001 (
            .O(N__19989),
            .I(N__19983));
    InMux I__3000 (
            .O(N__19988),
            .I(N__19980));
    LocalMux I__2999 (
            .O(N__19983),
            .I(N__19977));
    LocalMux I__2998 (
            .O(N__19980),
            .I(N__19972));
    Span4Mux_h I__2997 (
            .O(N__19977),
            .I(N__19972));
    Span4Mux_v I__2996 (
            .O(N__19972),
            .I(N__19969));
    Odrv4 I__2995 (
            .O(N__19969),
            .I(g0_0_0));
    InMux I__2994 (
            .O(N__19966),
            .I(N__19959));
    InMux I__2993 (
            .O(N__19965),
            .I(N__19959));
    InMux I__2992 (
            .O(N__19964),
            .I(N__19956));
    LocalMux I__2991 (
            .O(N__19959),
            .I(N_5_0));
    LocalMux I__2990 (
            .O(N__19956),
            .I(N_5_0));
    InMux I__2989 (
            .O(N__19951),
            .I(N__19948));
    LocalMux I__2988 (
            .O(N__19948),
            .I(N__19944));
    InMux I__2987 (
            .O(N__19947),
            .I(N__19941));
    Span4Mux_h I__2986 (
            .O(N__19944),
            .I(N__19936));
    LocalMux I__2985 (
            .O(N__19941),
            .I(N__19936));
    Odrv4 I__2984 (
            .O(N__19936),
            .I(b2v_inst11_un1_dutycycle_172_m3_amcf1));
    CascadeMux I__2983 (
            .O(N__19933),
            .I(N_73_mux_i_i_a7_4_0_1_cascade_));
    CascadeMux I__2982 (
            .O(N__19930),
            .I(\b2v_inst5.N_2897_i_cascade_ ));
    InMux I__2981 (
            .O(N__19927),
            .I(N__19924));
    LocalMux I__2980 (
            .O(N__19924),
            .I(\b2v_inst5.curr_state_0_0 ));
    CascadeMux I__2979 (
            .O(N__19921),
            .I(\b2v_inst5.m4_0_cascade_ ));
    CascadeMux I__2978 (
            .O(N__19918),
            .I(\b2v_inst11.g2_0_1_cascade_ ));
    CascadeMux I__2977 (
            .O(N__19915),
            .I(dutycycle_RNISSAOS1_0_5_cascade_));
    InMux I__2976 (
            .O(N__19912),
            .I(N__19909));
    LocalMux I__2975 (
            .O(N__19909),
            .I(\b2v_inst11.N_301 ));
    CascadeMux I__2974 (
            .O(N__19906),
            .I(\b2v_inst11.N_382_cascade_ ));
    CascadeMux I__2973 (
            .O(N__19903),
            .I(\b2v_inst11.g0_2_0_cascade_ ));
    CascadeMux I__2972 (
            .O(N__19900),
            .I(N__19897));
    InMux I__2971 (
            .O(N__19897),
            .I(N__19893));
    InMux I__2970 (
            .O(N__19896),
            .I(N__19890));
    LocalMux I__2969 (
            .O(N__19893),
            .I(N__19885));
    LocalMux I__2968 (
            .O(N__19890),
            .I(N__19885));
    Span4Mux_h I__2967 (
            .O(N__19885),
            .I(N__19882));
    Odrv4 I__2966 (
            .O(N__19882),
            .I(\b2v_inst11.N_430 ));
    InMux I__2965 (
            .O(N__19879),
            .I(N__19876));
    LocalMux I__2964 (
            .O(N__19876),
            .I(\b2v_inst11.func_state_RNIRF2E4Z0Z_0 ));
    IoInMux I__2963 (
            .O(N__19873),
            .I(N__19870));
    LocalMux I__2962 (
            .O(N__19870),
            .I(N__19867));
    IoSpan4Mux I__2961 (
            .O(N__19867),
            .I(N__19864));
    Span4Mux_s2_h I__2960 (
            .O(N__19864),
            .I(N__19861));
    Odrv4 I__2959 (
            .O(N__19861),
            .I(VCCST_EN_i_0_i));
    CascadeMux I__2958 (
            .O(N__19858),
            .I(N__19855));
    InMux I__2957 (
            .O(N__19855),
            .I(N__19852));
    LocalMux I__2956 (
            .O(N__19852),
            .I(\b2v_inst11.un1_clk_100khz_2_i_o3_sx ));
    InMux I__2955 (
            .O(N__19849),
            .I(N__19844));
    CascadeMux I__2954 (
            .O(N__19848),
            .I(N__19836));
    CascadeMux I__2953 (
            .O(N__19847),
            .I(N__19833));
    LocalMux I__2952 (
            .O(N__19844),
            .I(N__19830));
    InMux I__2951 (
            .O(N__19843),
            .I(N__19827));
    InMux I__2950 (
            .O(N__19842),
            .I(N__19822));
    InMux I__2949 (
            .O(N__19841),
            .I(N__19822));
    CascadeMux I__2948 (
            .O(N__19840),
            .I(N__19819));
    InMux I__2947 (
            .O(N__19839),
            .I(N__19816));
    InMux I__2946 (
            .O(N__19836),
            .I(N__19808));
    InMux I__2945 (
            .O(N__19833),
            .I(N__19808));
    Span4Mux_s2_h I__2944 (
            .O(N__19830),
            .I(N__19803));
    LocalMux I__2943 (
            .O(N__19827),
            .I(N__19803));
    LocalMux I__2942 (
            .O(N__19822),
            .I(N__19800));
    InMux I__2941 (
            .O(N__19819),
            .I(N__19797));
    LocalMux I__2940 (
            .O(N__19816),
            .I(N__19794));
    InMux I__2939 (
            .O(N__19815),
            .I(N__19787));
    InMux I__2938 (
            .O(N__19814),
            .I(N__19787));
    InMux I__2937 (
            .O(N__19813),
            .I(N__19787));
    LocalMux I__2936 (
            .O(N__19808),
            .I(N__19784));
    Span4Mux_v I__2935 (
            .O(N__19803),
            .I(N__19781));
    Span4Mux_s3_h I__2934 (
            .O(N__19800),
            .I(N__19778));
    LocalMux I__2933 (
            .O(N__19797),
            .I(N__19775));
    Odrv12 I__2932 (
            .O(N__19794),
            .I(\b2v_inst11.func_state ));
    LocalMux I__2931 (
            .O(N__19787),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__2930 (
            .O(N__19784),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__2929 (
            .O(N__19781),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__2928 (
            .O(N__19778),
            .I(\b2v_inst11.func_state ));
    Odrv4 I__2927 (
            .O(N__19775),
            .I(\b2v_inst11.func_state ));
    InMux I__2926 (
            .O(N__19762),
            .I(N__19757));
    InMux I__2925 (
            .O(N__19761),
            .I(N__19751));
    InMux I__2924 (
            .O(N__19760),
            .I(N__19751));
    LocalMux I__2923 (
            .O(N__19757),
            .I(N__19748));
    InMux I__2922 (
            .O(N__19756),
            .I(N__19745));
    LocalMux I__2921 (
            .O(N__19751),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    Odrv4 I__2920 (
            .O(N__19748),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    LocalMux I__2919 (
            .O(N__19745),
            .I(\b2v_inst11.func_state_RNI_0Z0Z_0 ));
    InMux I__2918 (
            .O(N__19738),
            .I(N__19735));
    LocalMux I__2917 (
            .O(N__19735),
            .I(\b2v_inst11.N_305 ));
    InMux I__2916 (
            .O(N__19732),
            .I(N__19729));
    LocalMux I__2915 (
            .O(N__19729),
            .I(N__19723));
    InMux I__2914 (
            .O(N__19728),
            .I(N__19720));
    InMux I__2913 (
            .O(N__19727),
            .I(N__19715));
    InMux I__2912 (
            .O(N__19726),
            .I(N__19715));
    Odrv4 I__2911 (
            .O(N__19723),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_6 ));
    LocalMux I__2910 (
            .O(N__19720),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_6 ));
    LocalMux I__2909 (
            .O(N__19715),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_6 ));
    CascadeMux I__2908 (
            .O(N__19708),
            .I(\b2v_inst11.dutycycle_RNIZ0Z_6_cascade_ ));
    CascadeMux I__2907 (
            .O(N__19705),
            .I(\b2v_inst11.i2_mux_cascade_ ));
    CascadeMux I__2906 (
            .O(N__19702),
            .I(\b2v_inst11.N_307_cascade_ ));
    InMux I__2905 (
            .O(N__19699),
            .I(N__19696));
    LocalMux I__2904 (
            .O(N__19696),
            .I(\b2v_inst11.N_234_N ));
    InMux I__2903 (
            .O(N__19693),
            .I(N__19690));
    LocalMux I__2902 (
            .O(N__19690),
            .I(N__19687));
    Odrv4 I__2901 (
            .O(N__19687),
            .I(\b2v_inst11.N_308 ));
    CascadeMux I__2900 (
            .O(N__19684),
            .I(\b2v_inst11.N_234_N_cascade_ ));
    CascadeMux I__2899 (
            .O(N__19681),
            .I(\b2v_inst11.func_state_RNI9R6T4Z0Z_1_cascade_ ));
    InMux I__2898 (
            .O(N__19678),
            .I(N__19675));
    LocalMux I__2897 (
            .O(N__19675),
            .I(\b2v_inst11.func_state_RNI9R6T4Z0Z_1 ));
    CascadeMux I__2896 (
            .O(N__19672),
            .I(N__19669));
    InMux I__2895 (
            .O(N__19669),
            .I(N__19663));
    InMux I__2894 (
            .O(N__19668),
            .I(N__19663));
    LocalMux I__2893 (
            .O(N__19663),
            .I(\b2v_inst11.dutycycleZ1Z_11 ));
    InMux I__2892 (
            .O(N__19660),
            .I(N__19657));
    LocalMux I__2891 (
            .O(N__19657),
            .I(N__19654));
    Odrv4 I__2890 (
            .O(N__19654),
            .I(\b2v_inst11.N_159 ));
    InMux I__2889 (
            .O(N__19651),
            .I(N__19648));
    LocalMux I__2888 (
            .O(N__19648),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ));
    CascadeMux I__2887 (
            .O(N__19645),
            .I(\b2v_inst11.N_155_N_cascade_ ));
    CascadeMux I__2886 (
            .O(N__19642),
            .I(\b2v_inst11.dutycycle_en_11_cascade_ ));
    InMux I__2885 (
            .O(N__19639),
            .I(N__19636));
    LocalMux I__2884 (
            .O(N__19636),
            .I(\b2v_inst11.g2_0 ));
    CascadeMux I__2883 (
            .O(N__19633),
            .I(\b2v_inst11.dutycycle_eena_8_cascade_ ));
    InMux I__2882 (
            .O(N__19630),
            .I(N__19627));
    LocalMux I__2881 (
            .O(N__19627),
            .I(\b2v_inst11.dutycycle_rst_7 ));
    InMux I__2880 (
            .O(N__19624),
            .I(N__19618));
    InMux I__2879 (
            .O(N__19623),
            .I(N__19618));
    LocalMux I__2878 (
            .O(N__19618),
            .I(\b2v_inst11.dutycycle_0_3 ));
    CascadeMux I__2877 (
            .O(N__19615),
            .I(\b2v_inst11.dutycycle_rst_7_cascade_ ));
    InMux I__2876 (
            .O(N__19612),
            .I(N__19609));
    LocalMux I__2875 (
            .O(N__19609),
            .I(\b2v_inst11.dutycycle_eena_8 ));
    CascadeMux I__2874 (
            .O(N__19606),
            .I(\b2v_inst11.dutycycleZ0Z_3_cascade_ ));
    InMux I__2873 (
            .O(N__19603),
            .I(N__19600));
    LocalMux I__2872 (
            .O(N__19600),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_0_d_0 ));
    InMux I__2871 (
            .O(N__19597),
            .I(N__19594));
    LocalMux I__2870 (
            .O(N__19594),
            .I(N__19591));
    Odrv4 I__2869 (
            .O(N__19591),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_0_ccf1 ));
    CascadeMux I__2868 (
            .O(N__19588),
            .I(N__19585));
    InMux I__2867 (
            .O(N__19585),
            .I(N__19582));
    LocalMux I__2866 (
            .O(N__19582),
            .I(\b2v_inst11.un1_clk_100khz_43_and_i_0_c ));
    InMux I__2865 (
            .O(N__19579),
            .I(N__19573));
    InMux I__2864 (
            .O(N__19578),
            .I(N__19573));
    LocalMux I__2863 (
            .O(N__19573),
            .I(N__19570));
    Odrv4 I__2862 (
            .O(N__19570),
            .I(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ));
    InMux I__2861 (
            .O(N__19567),
            .I(N__19564));
    LocalMux I__2860 (
            .O(N__19564),
            .I(N__19560));
    InMux I__2859 (
            .O(N__19563),
            .I(N__19557));
    Span4Mux_v I__2858 (
            .O(N__19560),
            .I(N__19554));
    LocalMux I__2857 (
            .O(N__19557),
            .I(\b2v_inst11.count_off_1_6 ));
    Odrv4 I__2856 (
            .O(N__19554),
            .I(\b2v_inst11.count_off_1_6 ));
    InMux I__2855 (
            .O(N__19549),
            .I(N__19543));
    InMux I__2854 (
            .O(N__19548),
            .I(N__19543));
    LocalMux I__2853 (
            .O(N__19543),
            .I(N__19540));
    Odrv4 I__2852 (
            .O(N__19540),
            .I(\b2v_inst11.count_offZ0Z_7 ));
    CascadeMux I__2851 (
            .O(N__19537),
            .I(N__19527));
    CEMux I__2850 (
            .O(N__19536),
            .I(N__19522));
    InMux I__2849 (
            .O(N__19535),
            .I(N__19510));
    InMux I__2848 (
            .O(N__19534),
            .I(N__19510));
    InMux I__2847 (
            .O(N__19533),
            .I(N__19503));
    InMux I__2846 (
            .O(N__19532),
            .I(N__19503));
    InMux I__2845 (
            .O(N__19531),
            .I(N__19503));
    InMux I__2844 (
            .O(N__19530),
            .I(N__19496));
    InMux I__2843 (
            .O(N__19527),
            .I(N__19496));
    CEMux I__2842 (
            .O(N__19526),
            .I(N__19496));
    CEMux I__2841 (
            .O(N__19525),
            .I(N__19491));
    LocalMux I__2840 (
            .O(N__19522),
            .I(N__19481));
    CEMux I__2839 (
            .O(N__19521),
            .I(N__19476));
    InMux I__2838 (
            .O(N__19520),
            .I(N__19476));
    InMux I__2837 (
            .O(N__19519),
            .I(N__19465));
    InMux I__2836 (
            .O(N__19518),
            .I(N__19465));
    CEMux I__2835 (
            .O(N__19517),
            .I(N__19465));
    InMux I__2834 (
            .O(N__19516),
            .I(N__19465));
    InMux I__2833 (
            .O(N__19515),
            .I(N__19465));
    LocalMux I__2832 (
            .O(N__19510),
            .I(N__19462));
    LocalMux I__2831 (
            .O(N__19503),
            .I(N__19459));
    LocalMux I__2830 (
            .O(N__19496),
            .I(N__19455));
    InMux I__2829 (
            .O(N__19495),
            .I(N__19450));
    InMux I__2828 (
            .O(N__19494),
            .I(N__19450));
    LocalMux I__2827 (
            .O(N__19491),
            .I(N__19447));
    InMux I__2826 (
            .O(N__19490),
            .I(N__19438));
    InMux I__2825 (
            .O(N__19489),
            .I(N__19438));
    InMux I__2824 (
            .O(N__19488),
            .I(N__19438));
    InMux I__2823 (
            .O(N__19487),
            .I(N__19438));
    CascadeMux I__2822 (
            .O(N__19486),
            .I(N__19435));
    CascadeMux I__2821 (
            .O(N__19485),
            .I(N__19432));
    CEMux I__2820 (
            .O(N__19484),
            .I(N__19428));
    Span4Mux_s3_v I__2819 (
            .O(N__19481),
            .I(N__19421));
    LocalMux I__2818 (
            .O(N__19476),
            .I(N__19421));
    LocalMux I__2817 (
            .O(N__19465),
            .I(N__19421));
    Span4Mux_h I__2816 (
            .O(N__19462),
            .I(N__19416));
    Span4Mux_h I__2815 (
            .O(N__19459),
            .I(N__19416));
    InMux I__2814 (
            .O(N__19458),
            .I(N__19413));
    Span4Mux_v I__2813 (
            .O(N__19455),
            .I(N__19410));
    LocalMux I__2812 (
            .O(N__19450),
            .I(N__19407));
    Span4Mux_s3_v I__2811 (
            .O(N__19447),
            .I(N__19402));
    LocalMux I__2810 (
            .O(N__19438),
            .I(N__19402));
    InMux I__2809 (
            .O(N__19435),
            .I(N__19395));
    InMux I__2808 (
            .O(N__19432),
            .I(N__19395));
    InMux I__2807 (
            .O(N__19431),
            .I(N__19395));
    LocalMux I__2806 (
            .O(N__19428),
            .I(N__19392));
    Span4Mux_v I__2805 (
            .O(N__19421),
            .I(N__19389));
    Span4Mux_v I__2804 (
            .O(N__19416),
            .I(N__19384));
    LocalMux I__2803 (
            .O(N__19413),
            .I(N__19384));
    Span4Mux_h I__2802 (
            .O(N__19410),
            .I(N__19379));
    Span4Mux_h I__2801 (
            .O(N__19407),
            .I(N__19379));
    Span4Mux_h I__2800 (
            .O(N__19402),
            .I(N__19374));
    LocalMux I__2799 (
            .O(N__19395),
            .I(N__19374));
    Odrv12 I__2798 (
            .O(N__19392),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2797 (
            .O(N__19389),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2796 (
            .O(N__19384),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2795 (
            .O(N__19379),
            .I(\b2v_inst11.count_off_enZ0 ));
    Odrv4 I__2794 (
            .O(N__19374),
            .I(\b2v_inst11.count_off_enZ0 ));
    InMux I__2793 (
            .O(N__19363),
            .I(N__19357));
    InMux I__2792 (
            .O(N__19362),
            .I(N__19357));
    LocalMux I__2791 (
            .O(N__19357),
            .I(N__19354));
    Odrv4 I__2790 (
            .O(N__19354),
            .I(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ));
    CascadeMux I__2789 (
            .O(N__19351),
            .I(N__19344));
    InMux I__2788 (
            .O(N__19350),
            .I(N__19310));
    InMux I__2787 (
            .O(N__19349),
            .I(N__19310));
    InMux I__2786 (
            .O(N__19348),
            .I(N__19310));
    InMux I__2785 (
            .O(N__19347),
            .I(N__19305));
    InMux I__2784 (
            .O(N__19344),
            .I(N__19305));
    InMux I__2783 (
            .O(N__19343),
            .I(N__19302));
    InMux I__2782 (
            .O(N__19342),
            .I(N__19293));
    InMux I__2781 (
            .O(N__19341),
            .I(N__19293));
    InMux I__2780 (
            .O(N__19340),
            .I(N__19293));
    InMux I__2779 (
            .O(N__19339),
            .I(N__19293));
    InMux I__2778 (
            .O(N__19338),
            .I(N__19286));
    InMux I__2777 (
            .O(N__19337),
            .I(N__19286));
    InMux I__2776 (
            .O(N__19336),
            .I(N__19286));
    InMux I__2775 (
            .O(N__19335),
            .I(N__19273));
    InMux I__2774 (
            .O(N__19334),
            .I(N__19273));
    InMux I__2773 (
            .O(N__19333),
            .I(N__19273));
    InMux I__2772 (
            .O(N__19332),
            .I(N__19273));
    InMux I__2771 (
            .O(N__19331),
            .I(N__19273));
    InMux I__2770 (
            .O(N__19330),
            .I(N__19273));
    InMux I__2769 (
            .O(N__19329),
            .I(N__19260));
    InMux I__2768 (
            .O(N__19328),
            .I(N__19260));
    InMux I__2767 (
            .O(N__19327),
            .I(N__19260));
    InMux I__2766 (
            .O(N__19326),
            .I(N__19260));
    InMux I__2765 (
            .O(N__19325),
            .I(N__19260));
    InMux I__2764 (
            .O(N__19324),
            .I(N__19260));
    InMux I__2763 (
            .O(N__19323),
            .I(N__19245));
    InMux I__2762 (
            .O(N__19322),
            .I(N__19245));
    InMux I__2761 (
            .O(N__19321),
            .I(N__19245));
    InMux I__2760 (
            .O(N__19320),
            .I(N__19245));
    InMux I__2759 (
            .O(N__19319),
            .I(N__19245));
    InMux I__2758 (
            .O(N__19318),
            .I(N__19245));
    InMux I__2757 (
            .O(N__19317),
            .I(N__19245));
    LocalMux I__2756 (
            .O(N__19310),
            .I(N__19240));
    LocalMux I__2755 (
            .O(N__19305),
            .I(N__19240));
    LocalMux I__2754 (
            .O(N__19302),
            .I(N__19229));
    LocalMux I__2753 (
            .O(N__19293),
            .I(N__19229));
    LocalMux I__2752 (
            .O(N__19286),
            .I(N__19229));
    LocalMux I__2751 (
            .O(N__19273),
            .I(N__19229));
    LocalMux I__2750 (
            .O(N__19260),
            .I(N__19229));
    LocalMux I__2749 (
            .O(N__19245),
            .I(N__19224));
    Span4Mux_h I__2748 (
            .O(N__19240),
            .I(N__19224));
    Span4Mux_v I__2747 (
            .O(N__19229),
            .I(N__19221));
    Odrv4 I__2746 (
            .O(N__19224),
            .I(\b2v_inst11.N_125 ));
    Odrv4 I__2745 (
            .O(N__19221),
            .I(\b2v_inst11.N_125 ));
    InMux I__2744 (
            .O(N__19216),
            .I(N__19212));
    InMux I__2743 (
            .O(N__19215),
            .I(N__19209));
    LocalMux I__2742 (
            .O(N__19212),
            .I(N__19206));
    LocalMux I__2741 (
            .O(N__19209),
            .I(N__19203));
    Span4Mux_s2_v I__2740 (
            .O(N__19206),
            .I(N__19198));
    Span4Mux_s2_v I__2739 (
            .O(N__19203),
            .I(N__19198));
    Odrv4 I__2738 (
            .O(N__19198),
            .I(\b2v_inst11.count_off_1_7 ));
    CascadeMux I__2737 (
            .O(N__19195),
            .I(N__19192));
    InMux I__2736 (
            .O(N__19192),
            .I(N__19189));
    LocalMux I__2735 (
            .O(N__19189),
            .I(\b2v_inst11.g0_3_0 ));
    InMux I__2734 (
            .O(N__19186),
            .I(N__19182));
    InMux I__2733 (
            .O(N__19185),
            .I(N__19179));
    LocalMux I__2732 (
            .O(N__19182),
            .I(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ));
    LocalMux I__2731 (
            .O(N__19179),
            .I(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ));
    InMux I__2730 (
            .O(N__19174),
            .I(N__19168));
    InMux I__2729 (
            .O(N__19173),
            .I(N__19168));
    LocalMux I__2728 (
            .O(N__19168),
            .I(\b2v_inst11.count_offZ0Z_2 ));
    InMux I__2727 (
            .O(N__19165),
            .I(N__19161));
    InMux I__2726 (
            .O(N__19164),
            .I(N__19158));
    LocalMux I__2725 (
            .O(N__19161),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    LocalMux I__2724 (
            .O(N__19158),
            .I(\b2v_inst11.count_offZ0Z_5 ));
    CascadeMux I__2723 (
            .O(N__19153),
            .I(N__19150));
    InMux I__2722 (
            .O(N__19150),
            .I(N__19146));
    InMux I__2721 (
            .O(N__19149),
            .I(N__19142));
    LocalMux I__2720 (
            .O(N__19146),
            .I(N__19139));
    InMux I__2719 (
            .O(N__19145),
            .I(N__19136));
    LocalMux I__2718 (
            .O(N__19142),
            .I(N__19133));
    Span4Mux_h I__2717 (
            .O(N__19139),
            .I(N__19126));
    LocalMux I__2716 (
            .O(N__19136),
            .I(N__19126));
    Span4Mux_v I__2715 (
            .O(N__19133),
            .I(N__19126));
    Odrv4 I__2714 (
            .O(N__19126),
            .I(\b2v_inst11.count_offZ0Z_1 ));
    InMux I__2713 (
            .O(N__19123),
            .I(N__19120));
    LocalMux I__2712 (
            .O(N__19120),
            .I(\b2v_inst11.un34_clk_100khz_0 ));
    InMux I__2711 (
            .O(N__19117),
            .I(N__19114));
    LocalMux I__2710 (
            .O(N__19114),
            .I(\b2v_inst11.un34_clk_100khz_2 ));
    CascadeMux I__2709 (
            .O(N__19111),
            .I(\b2v_inst11.un34_clk_100khz_1_cascade_ ));
    InMux I__2708 (
            .O(N__19108),
            .I(N__19105));
    LocalMux I__2707 (
            .O(N__19105),
            .I(N__19102));
    Odrv4 I__2706 (
            .O(N__19102),
            .I(\b2v_inst11.un34_clk_100khz_3 ));
    InMux I__2705 (
            .O(N__19099),
            .I(N__19096));
    LocalMux I__2704 (
            .O(N__19096),
            .I(\b2v_inst11.un34_clk_100khz_12 ));
    CascadeMux I__2703 (
            .O(N__19093),
            .I(N__19089));
    InMux I__2702 (
            .O(N__19092),
            .I(N__19084));
    InMux I__2701 (
            .O(N__19089),
            .I(N__19084));
    LocalMux I__2700 (
            .O(N__19084),
            .I(\b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ));
    CascadeMux I__2699 (
            .O(N__19081),
            .I(N__19078));
    InMux I__2698 (
            .O(N__19078),
            .I(N__19075));
    LocalMux I__2697 (
            .O(N__19075),
            .I(\b2v_inst11.count_off_0_5 ));
    InMux I__2696 (
            .O(N__19072),
            .I(N__19069));
    LocalMux I__2695 (
            .O(N__19069),
            .I(N__19066));
    Span4Mux_s2_h I__2694 (
            .O(N__19066),
            .I(N__19062));
    InMux I__2693 (
            .O(N__19065),
            .I(N__19059));
    Span4Mux_v I__2692 (
            .O(N__19062),
            .I(N__19056));
    LocalMux I__2691 (
            .O(N__19059),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    Odrv4 I__2690 (
            .O(N__19056),
            .I(\b2v_inst11.count_offZ0Z_6 ));
    InMux I__2689 (
            .O(N__19051),
            .I(N__19045));
    InMux I__2688 (
            .O(N__19050),
            .I(N__19045));
    LocalMux I__2687 (
            .O(N__19045),
            .I(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ));
    InMux I__2686 (
            .O(N__19042),
            .I(N__19039));
    LocalMux I__2685 (
            .O(N__19039),
            .I(\b2v_inst11.count_off_1_9 ));
    InMux I__2684 (
            .O(N__19036),
            .I(N__19032));
    InMux I__2683 (
            .O(N__19035),
            .I(N__19029));
    LocalMux I__2682 (
            .O(N__19032),
            .I(\b2v_inst11.count_offZ0Z_9 ));
    LocalMux I__2681 (
            .O(N__19029),
            .I(\b2v_inst11.count_offZ0Z_9 ));
    CascadeMux I__2680 (
            .O(N__19024),
            .I(\b2v_inst11.count_off_1_9_cascade_ ));
    InMux I__2679 (
            .O(N__19021),
            .I(N__19018));
    LocalMux I__2678 (
            .O(N__19018),
            .I(\b2v_inst11.un3_count_off_1_axb_9 ));
    CascadeMux I__2677 (
            .O(N__19015),
            .I(\b2v_inst11.count_off_1_3_cascade_ ));
    InMux I__2676 (
            .O(N__19012),
            .I(N__19009));
    LocalMux I__2675 (
            .O(N__19009),
            .I(\b2v_inst11.un3_count_off_1_axb_3 ));
    InMux I__2674 (
            .O(N__19006),
            .I(N__19003));
    LocalMux I__2673 (
            .O(N__19003),
            .I(\b2v_inst11.count_offZ0Z_4 ));
    InMux I__2672 (
            .O(N__19000),
            .I(N__18997));
    LocalMux I__2671 (
            .O(N__18997),
            .I(\b2v_inst11.count_off_1_3 ));
    CascadeMux I__2670 (
            .O(N__18994),
            .I(\b2v_inst11.count_offZ0Z_4_cascade_ ));
    InMux I__2669 (
            .O(N__18991),
            .I(N__18985));
    InMux I__2668 (
            .O(N__18990),
            .I(N__18985));
    LocalMux I__2667 (
            .O(N__18985),
            .I(\b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ));
    InMux I__2666 (
            .O(N__18982),
            .I(N__18976));
    InMux I__2665 (
            .O(N__18981),
            .I(N__18976));
    LocalMux I__2664 (
            .O(N__18976),
            .I(\b2v_inst11.count_offZ0Z_3 ));
    CascadeMux I__2663 (
            .O(N__18973),
            .I(N__18970));
    InMux I__2662 (
            .O(N__18970),
            .I(N__18964));
    InMux I__2661 (
            .O(N__18969),
            .I(N__18964));
    LocalMux I__2660 (
            .O(N__18964),
            .I(\b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ));
    CascadeMux I__2659 (
            .O(N__18961),
            .I(N__18958));
    InMux I__2658 (
            .O(N__18958),
            .I(N__18955));
    LocalMux I__2657 (
            .O(N__18955),
            .I(\b2v_inst11.count_off_0_4 ));
    InMux I__2656 (
            .O(N__18952),
            .I(N__18949));
    LocalMux I__2655 (
            .O(N__18949),
            .I(\b2v_inst11.count_off_0_14 ));
    CascadeMux I__2654 (
            .O(N__18946),
            .I(N__18943));
    InMux I__2653 (
            .O(N__18943),
            .I(N__18937));
    InMux I__2652 (
            .O(N__18942),
            .I(N__18937));
    LocalMux I__2651 (
            .O(N__18937),
            .I(\b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ));
    InMux I__2650 (
            .O(N__18934),
            .I(N__18930));
    InMux I__2649 (
            .O(N__18933),
            .I(N__18927));
    LocalMux I__2648 (
            .O(N__18930),
            .I(\b2v_inst11.count_offZ0Z_14 ));
    LocalMux I__2647 (
            .O(N__18927),
            .I(\b2v_inst11.count_offZ0Z_14 ));
    InMux I__2646 (
            .O(N__18922),
            .I(N__18916));
    InMux I__2645 (
            .O(N__18921),
            .I(N__18916));
    LocalMux I__2644 (
            .O(N__18916),
            .I(\b2v_inst11.count_off_1_2 ));
    InMux I__2643 (
            .O(N__18913),
            .I(N__18910));
    LocalMux I__2642 (
            .O(N__18910),
            .I(\b2v_inst11.un3_count_off_1_axb_2 ));
    InMux I__2641 (
            .O(N__18907),
            .I(\b2v_inst200.un2_count_1_cry_10 ));
    InMux I__2640 (
            .O(N__18904),
            .I(N__18900));
    InMux I__2639 (
            .O(N__18903),
            .I(N__18897));
    LocalMux I__2638 (
            .O(N__18900),
            .I(N__18894));
    LocalMux I__2637 (
            .O(N__18897),
            .I(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ));
    Odrv4 I__2636 (
            .O(N__18894),
            .I(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ));
    InMux I__2635 (
            .O(N__18889),
            .I(\b2v_inst200.un2_count_1_cry_11 ));
    InMux I__2634 (
            .O(N__18886),
            .I(\b2v_inst200.un2_count_1_cry_12 ));
    InMux I__2633 (
            .O(N__18883),
            .I(\b2v_inst200.un2_count_1_cry_13 ));
    InMux I__2632 (
            .O(N__18880),
            .I(\b2v_inst200.un2_count_1_cry_14 ));
    InMux I__2631 (
            .O(N__18877),
            .I(bfn_5_3_0_));
    InMux I__2630 (
            .O(N__18874),
            .I(\b2v_inst200.un2_count_1_cry_16 ));
    InMux I__2629 (
            .O(N__18871),
            .I(N__18868));
    LocalMux I__2628 (
            .O(N__18868),
            .I(\b2v_inst200.count_0_17 ));
    InMux I__2627 (
            .O(N__18865),
            .I(N__18861));
    InMux I__2626 (
            .O(N__18864),
            .I(N__18858));
    LocalMux I__2625 (
            .O(N__18861),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    LocalMux I__2624 (
            .O(N__18858),
            .I(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ));
    InMux I__2623 (
            .O(N__18853),
            .I(N__18849));
    InMux I__2622 (
            .O(N__18852),
            .I(N__18846));
    LocalMux I__2621 (
            .O(N__18849),
            .I(\b2v_inst200.countZ0Z_3 ));
    LocalMux I__2620 (
            .O(N__18846),
            .I(\b2v_inst200.countZ0Z_3 ));
    InMux I__2619 (
            .O(N__18841),
            .I(N__18835));
    InMux I__2618 (
            .O(N__18840),
            .I(N__18835));
    LocalMux I__2617 (
            .O(N__18835),
            .I(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ));
    InMux I__2616 (
            .O(N__18832),
            .I(\b2v_inst200.un2_count_1_cry_2 ));
    InMux I__2615 (
            .O(N__18829),
            .I(N__18825));
    InMux I__2614 (
            .O(N__18828),
            .I(N__18822));
    LocalMux I__2613 (
            .O(N__18825),
            .I(\b2v_inst200.countZ0Z_4 ));
    LocalMux I__2612 (
            .O(N__18822),
            .I(\b2v_inst200.countZ0Z_4 ));
    InMux I__2611 (
            .O(N__18817),
            .I(N__18813));
    InMux I__2610 (
            .O(N__18816),
            .I(N__18810));
    LocalMux I__2609 (
            .O(N__18813),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    LocalMux I__2608 (
            .O(N__18810),
            .I(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ));
    InMux I__2607 (
            .O(N__18805),
            .I(\b2v_inst200.un2_count_1_cry_3 ));
    InMux I__2606 (
            .O(N__18802),
            .I(N__18799));
    LocalMux I__2605 (
            .O(N__18799),
            .I(N__18795));
    InMux I__2604 (
            .O(N__18798),
            .I(N__18792));
    Span4Mux_v I__2603 (
            .O(N__18795),
            .I(N__18789));
    LocalMux I__2602 (
            .O(N__18792),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    Odrv4 I__2601 (
            .O(N__18789),
            .I(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ));
    InMux I__2600 (
            .O(N__18784),
            .I(\b2v_inst200.un2_count_1_cry_4 ));
    InMux I__2599 (
            .O(N__18781),
            .I(\b2v_inst200.un2_count_1_cry_5_cZ0 ));
    InMux I__2598 (
            .O(N__18778),
            .I(N__18775));
    LocalMux I__2597 (
            .O(N__18775),
            .I(N__18771));
    InMux I__2596 (
            .O(N__18774),
            .I(N__18768));
    Span4Mux_h I__2595 (
            .O(N__18771),
            .I(N__18765));
    LocalMux I__2594 (
            .O(N__18768),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    Odrv4 I__2593 (
            .O(N__18765),
            .I(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ));
    InMux I__2592 (
            .O(N__18760),
            .I(\b2v_inst200.un2_count_1_cry_6 ));
    InMux I__2591 (
            .O(N__18757),
            .I(bfn_5_2_0_));
    InMux I__2590 (
            .O(N__18754),
            .I(\b2v_inst200.un2_count_1_cry_8 ));
    InMux I__2589 (
            .O(N__18751),
            .I(\b2v_inst200.un2_count_1_cry_9 ));
    CascadeMux I__2588 (
            .O(N__18748),
            .I(N__18745));
    InMux I__2587 (
            .O(N__18745),
            .I(N__18742));
    LocalMux I__2586 (
            .O(N__18742),
            .I(N__18737));
    InMux I__2585 (
            .O(N__18741),
            .I(N__18731));
    InMux I__2584 (
            .O(N__18740),
            .I(N__18731));
    Span4Mux_s3_h I__2583 (
            .O(N__18737),
            .I(N__18728));
    InMux I__2582 (
            .O(N__18736),
            .I(N__18725));
    LocalMux I__2581 (
            .O(N__18731),
            .I(\b2v_inst20.counterZ0Z_0 ));
    Odrv4 I__2580 (
            .O(N__18728),
            .I(\b2v_inst20.counterZ0Z_0 ));
    LocalMux I__2579 (
            .O(N__18725),
            .I(\b2v_inst20.counterZ0Z_0 ));
    CascadeMux I__2578 (
            .O(N__18718),
            .I(N__18714));
    InMux I__2577 (
            .O(N__18717),
            .I(N__18709));
    InMux I__2576 (
            .O(N__18714),
            .I(N__18709));
    LocalMux I__2575 (
            .O(N__18709),
            .I(N__18706));
    Span4Mux_s2_h I__2574 (
            .O(N__18706),
            .I(N__18703));
    Span4Mux_v I__2573 (
            .O(N__18703),
            .I(N__18700));
    Span4Mux_v I__2572 (
            .O(N__18700),
            .I(N__18696));
    InMux I__2571 (
            .O(N__18699),
            .I(N__18693));
    Odrv4 I__2570 (
            .O(N__18696),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    LocalMux I__2569 (
            .O(N__18693),
            .I(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    InMux I__2568 (
            .O(N__18688),
            .I(N__18685));
    LocalMux I__2567 (
            .O(N__18685),
            .I(N__18682));
    Span4Mux_h I__2566 (
            .O(N__18682),
            .I(N__18679));
    Odrv4 I__2565 (
            .O(N__18679),
            .I(\b2v_inst20.counter_1_cry_3_THRU_CO ));
    InMux I__2564 (
            .O(N__18676),
            .I(N__18673));
    LocalMux I__2563 (
            .O(N__18673),
            .I(N__18669));
    InMux I__2562 (
            .O(N__18672),
            .I(N__18665));
    Span4Mux_v I__2561 (
            .O(N__18669),
            .I(N__18662));
    InMux I__2560 (
            .O(N__18668),
            .I(N__18659));
    LocalMux I__2559 (
            .O(N__18665),
            .I(\b2v_inst20.counterZ0Z_4 ));
    Odrv4 I__2558 (
            .O(N__18662),
            .I(\b2v_inst20.counterZ0Z_4 ));
    LocalMux I__2557 (
            .O(N__18659),
            .I(\b2v_inst20.counterZ0Z_4 ));
    InMux I__2556 (
            .O(N__18652),
            .I(N__18649));
    LocalMux I__2555 (
            .O(N__18649),
            .I(N__18646));
    Span4Mux_h I__2554 (
            .O(N__18646),
            .I(N__18643));
    Odrv4 I__2553 (
            .O(N__18643),
            .I(\b2v_inst20.counter_1_cry_4_THRU_CO ));
    IoInMux I__2552 (
            .O(N__18640),
            .I(N__18637));
    LocalMux I__2551 (
            .O(N__18637),
            .I(N__18632));
    IoInMux I__2550 (
            .O(N__18636),
            .I(N__18629));
    IoInMux I__2549 (
            .O(N__18635),
            .I(N__18626));
    IoSpan4Mux I__2548 (
            .O(N__18632),
            .I(N__18621));
    LocalMux I__2547 (
            .O(N__18629),
            .I(N__18621));
    LocalMux I__2546 (
            .O(N__18626),
            .I(N__18618));
    IoSpan4Mux I__2545 (
            .O(N__18621),
            .I(N__18615));
    Span12Mux_s0_v I__2544 (
            .O(N__18618),
            .I(N__18612));
    Odrv4 I__2543 (
            .O(N__18615),
            .I(delayed_vccin_vccinaux_ok_RNI8L1J7_0));
    Odrv12 I__2542 (
            .O(N__18612),
            .I(delayed_vccin_vccinaux_ok_RNI8L1J7_0));
    InMux I__2541 (
            .O(N__18607),
            .I(N__18604));
    LocalMux I__2540 (
            .O(N__18604),
            .I(N__18601));
    Span4Mux_s3_v I__2539 (
            .O(N__18601),
            .I(N__18598));
    Odrv4 I__2538 (
            .O(N__18598),
            .I(\b2v_inst20.counter_1_cry_1_THRU_CO ));
    InMux I__2537 (
            .O(N__18595),
            .I(N__18592));
    LocalMux I__2536 (
            .O(N__18592),
            .I(N__18588));
    InMux I__2535 (
            .O(N__18591),
            .I(N__18584));
    Span4Mux_s3_h I__2534 (
            .O(N__18588),
            .I(N__18581));
    InMux I__2533 (
            .O(N__18587),
            .I(N__18578));
    LocalMux I__2532 (
            .O(N__18584),
            .I(\b2v_inst20.counterZ0Z_2 ));
    Odrv4 I__2531 (
            .O(N__18581),
            .I(\b2v_inst20.counterZ0Z_2 ));
    LocalMux I__2530 (
            .O(N__18578),
            .I(\b2v_inst20.counterZ0Z_2 ));
    CascadeMux I__2529 (
            .O(N__18571),
            .I(N__18568));
    InMux I__2528 (
            .O(N__18568),
            .I(N__18564));
    InMux I__2527 (
            .O(N__18567),
            .I(N__18561));
    LocalMux I__2526 (
            .O(N__18564),
            .I(\b2v_inst200.countZ0Z_1 ));
    LocalMux I__2525 (
            .O(N__18561),
            .I(\b2v_inst200.countZ0Z_1 ));
    InMux I__2524 (
            .O(N__18556),
            .I(N__18550));
    InMux I__2523 (
            .O(N__18555),
            .I(N__18550));
    LocalMux I__2522 (
            .O(N__18550),
            .I(\b2v_inst200.count_RNIC03N_5Z0Z_0 ));
    InMux I__2521 (
            .O(N__18547),
            .I(\b2v_inst200.un2_count_1_cry_1_cy ));
    InMux I__2520 (
            .O(N__18544),
            .I(N__18540));
    InMux I__2519 (
            .O(N__18543),
            .I(N__18537));
    LocalMux I__2518 (
            .O(N__18540),
            .I(\b2v_inst200.countZ0Z_2 ));
    LocalMux I__2517 (
            .O(N__18537),
            .I(\b2v_inst200.countZ0Z_2 ));
    InMux I__2516 (
            .O(N__18532),
            .I(N__18526));
    InMux I__2515 (
            .O(N__18531),
            .I(N__18526));
    LocalMux I__2514 (
            .O(N__18526),
            .I(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ));
    InMux I__2513 (
            .O(N__18523),
            .I(\b2v_inst200.un2_count_1_cry_1 ));
    InMux I__2512 (
            .O(N__18520),
            .I(N__18517));
    LocalMux I__2511 (
            .O(N__18517),
            .I(N__18514));
    Odrv4 I__2510 (
            .O(N__18514),
            .I(\b2v_inst20.un4_counter_0_and ));
    CascadeMux I__2509 (
            .O(N__18511),
            .I(\b2v_inst11.N_381_cascade_ ));
    InMux I__2508 (
            .O(N__18508),
            .I(N__18505));
    LocalMux I__2507 (
            .O(N__18505),
            .I(N__18502));
    Odrv12 I__2506 (
            .O(N__18502),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ));
    CascadeMux I__2505 (
            .O(N__18499),
            .I(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ));
    InMux I__2504 (
            .O(N__18496),
            .I(N__18493));
    LocalMux I__2503 (
            .O(N__18493),
            .I(N__18490));
    Span12Mux_s3_h I__2502 (
            .O(N__18490),
            .I(N__18487));
    Odrv12 I__2501 (
            .O(N__18487),
            .I(\b2v_inst11.N_381_0 ));
    InMux I__2500 (
            .O(N__18484),
            .I(N__18481));
    LocalMux I__2499 (
            .O(N__18481),
            .I(N__18478));
    Span4Mux_s2_v I__2498 (
            .O(N__18478),
            .I(N__18475));
    Span4Mux_v I__2497 (
            .O(N__18475),
            .I(N__18472));
    Span4Mux_v I__2496 (
            .O(N__18472),
            .I(N__18469));
    Odrv4 I__2495 (
            .O(N__18469),
            .I(N_15_i_0_a4_0_1));
    InMux I__2494 (
            .O(N__18466),
            .I(N__18463));
    LocalMux I__2493 (
            .O(N__18463),
            .I(N__18460));
    Span4Mux_s3_v I__2492 (
            .O(N__18460),
            .I(N__18457));
    Odrv4 I__2491 (
            .O(N__18457),
            .I(\b2v_inst20.counter_1_cry_2_THRU_CO ));
    InMux I__2490 (
            .O(N__18454),
            .I(N__18451));
    LocalMux I__2489 (
            .O(N__18451),
            .I(N__18447));
    CascadeMux I__2488 (
            .O(N__18450),
            .I(N__18443));
    Span4Mux_s3_h I__2487 (
            .O(N__18447),
            .I(N__18440));
    InMux I__2486 (
            .O(N__18446),
            .I(N__18435));
    InMux I__2485 (
            .O(N__18443),
            .I(N__18435));
    Odrv4 I__2484 (
            .O(N__18440),
            .I(\b2v_inst20.counterZ0Z_3 ));
    LocalMux I__2483 (
            .O(N__18435),
            .I(\b2v_inst20.counterZ0Z_3 ));
    InMux I__2482 (
            .O(N__18430),
            .I(N__18425));
    CascadeMux I__2481 (
            .O(N__18429),
            .I(N__18422));
    InMux I__2480 (
            .O(N__18428),
            .I(N__18419));
    LocalMux I__2479 (
            .O(N__18425),
            .I(N__18416));
    InMux I__2478 (
            .O(N__18422),
            .I(N__18413));
    LocalMux I__2477 (
            .O(N__18419),
            .I(N__18410));
    Span4Mux_s3_h I__2476 (
            .O(N__18416),
            .I(N__18407));
    LocalMux I__2475 (
            .O(N__18413),
            .I(N__18404));
    Span4Mux_s3_h I__2474 (
            .O(N__18410),
            .I(N__18401));
    Span4Mux_v I__2473 (
            .O(N__18407),
            .I(N__18396));
    Span4Mux_s3_h I__2472 (
            .O(N__18404),
            .I(N__18396));
    Odrv4 I__2471 (
            .O(N__18401),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    Odrv4 I__2470 (
            .O(N__18396),
            .I(\b2v_inst11.count_clkZ0Z_8 ));
    InMux I__2469 (
            .O(N__18391),
            .I(N__18388));
    LocalMux I__2468 (
            .O(N__18388),
            .I(N__18385));
    Span4Mux_v I__2467 (
            .O(N__18385),
            .I(N__18381));
    InMux I__2466 (
            .O(N__18384),
            .I(N__18378));
    Odrv4 I__2465 (
            .O(N__18381),
            .I(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ));
    LocalMux I__2464 (
            .O(N__18378),
            .I(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ));
    InMux I__2463 (
            .O(N__18373),
            .I(N__18370));
    LocalMux I__2462 (
            .O(N__18370),
            .I(N__18367));
    Span4Mux_h I__2461 (
            .O(N__18367),
            .I(N__18364));
    Odrv4 I__2460 (
            .O(N__18364),
            .I(\b2v_inst11.count_clk_0_2 ));
    InMux I__2459 (
            .O(N__18361),
            .I(N__18357));
    InMux I__2458 (
            .O(N__18360),
            .I(N__18353));
    LocalMux I__2457 (
            .O(N__18357),
            .I(N__18350));
    InMux I__2456 (
            .O(N__18356),
            .I(N__18347));
    LocalMux I__2455 (
            .O(N__18353),
            .I(N__18344));
    Span4Mux_h I__2454 (
            .O(N__18350),
            .I(N__18341));
    LocalMux I__2453 (
            .O(N__18347),
            .I(N__18338));
    Span4Mux_s3_h I__2452 (
            .O(N__18344),
            .I(N__18335));
    Span4Mux_v I__2451 (
            .O(N__18341),
            .I(N__18332));
    Span4Mux_s3_h I__2450 (
            .O(N__18338),
            .I(N__18329));
    Odrv4 I__2449 (
            .O(N__18335),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    Odrv4 I__2448 (
            .O(N__18332),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    Odrv4 I__2447 (
            .O(N__18329),
            .I(\b2v_inst11.count_clkZ0Z_2 ));
    CascadeMux I__2446 (
            .O(N__18322),
            .I(N__18317));
    InMux I__2445 (
            .O(N__18321),
            .I(N__18313));
    InMux I__2444 (
            .O(N__18320),
            .I(N__18308));
    InMux I__2443 (
            .O(N__18317),
            .I(N__18308));
    InMux I__2442 (
            .O(N__18316),
            .I(N__18305));
    LocalMux I__2441 (
            .O(N__18313),
            .I(N__18302));
    LocalMux I__2440 (
            .O(N__18308),
            .I(N__18299));
    LocalMux I__2439 (
            .O(N__18305),
            .I(N__18296));
    Span4Mux_s3_h I__2438 (
            .O(N__18302),
            .I(N__18293));
    Span4Mux_s3_h I__2437 (
            .O(N__18299),
            .I(N__18288));
    Span4Mux_s3_h I__2436 (
            .O(N__18296),
            .I(N__18288));
    Odrv4 I__2435 (
            .O(N__18293),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    Odrv4 I__2434 (
            .O(N__18288),
            .I(\b2v_inst11.count_clkZ0Z_5 ));
    InMux I__2433 (
            .O(N__18283),
            .I(N__18280));
    LocalMux I__2432 (
            .O(N__18280),
            .I(N__18276));
    InMux I__2431 (
            .O(N__18279),
            .I(N__18273));
    Odrv4 I__2430 (
            .O(N__18276),
            .I(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ));
    LocalMux I__2429 (
            .O(N__18273),
            .I(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ));
    InMux I__2428 (
            .O(N__18268),
            .I(N__18265));
    LocalMux I__2427 (
            .O(N__18265),
            .I(N__18262));
    Odrv4 I__2426 (
            .O(N__18262),
            .I(\b2v_inst11.count_clk_0_9 ));
    InMux I__2425 (
            .O(N__18259),
            .I(N__18249));
    InMux I__2424 (
            .O(N__18258),
            .I(N__18249));
    InMux I__2423 (
            .O(N__18257),
            .I(N__18249));
    InMux I__2422 (
            .O(N__18256),
            .I(N__18246));
    LocalMux I__2421 (
            .O(N__18249),
            .I(N__18243));
    LocalMux I__2420 (
            .O(N__18246),
            .I(N__18240));
    Span4Mux_s3_h I__2419 (
            .O(N__18243),
            .I(N__18237));
    Odrv4 I__2418 (
            .O(N__18240),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    Odrv4 I__2417 (
            .O(N__18237),
            .I(\b2v_inst11.count_clkZ0Z_9 ));
    InMux I__2416 (
            .O(N__18232),
            .I(N__18228));
    InMux I__2415 (
            .O(N__18231),
            .I(N__18225));
    LocalMux I__2414 (
            .O(N__18228),
            .I(N__18220));
    LocalMux I__2413 (
            .O(N__18225),
            .I(N__18220));
    Span4Mux_v I__2412 (
            .O(N__18220),
            .I(N__18217));
    Odrv4 I__2411 (
            .O(N__18217),
            .I(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ));
    InMux I__2410 (
            .O(N__18214),
            .I(N__18211));
    LocalMux I__2409 (
            .O(N__18211),
            .I(\b2v_inst11.count_clk_0_3 ));
    InMux I__2408 (
            .O(N__18208),
            .I(N__18204));
    InMux I__2407 (
            .O(N__18207),
            .I(N__18201));
    LocalMux I__2406 (
            .O(N__18204),
            .I(N__18198));
    LocalMux I__2405 (
            .O(N__18201),
            .I(N__18195));
    Span4Mux_v I__2404 (
            .O(N__18198),
            .I(N__18192));
    Span4Mux_h I__2403 (
            .O(N__18195),
            .I(N__18189));
    Odrv4 I__2402 (
            .O(N__18192),
            .I(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ));
    Odrv4 I__2401 (
            .O(N__18189),
            .I(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ));
    InMux I__2400 (
            .O(N__18184),
            .I(N__18181));
    LocalMux I__2399 (
            .O(N__18181),
            .I(\b2v_inst11.count_clk_0_5 ));
    InMux I__2398 (
            .O(N__18178),
            .I(N__18174));
    InMux I__2397 (
            .O(N__18177),
            .I(N__18171));
    LocalMux I__2396 (
            .O(N__18174),
            .I(N__18168));
    LocalMux I__2395 (
            .O(N__18171),
            .I(N__18165));
    Span4Mux_v I__2394 (
            .O(N__18168),
            .I(N__18162));
    Span4Mux_h I__2393 (
            .O(N__18165),
            .I(N__18159));
    Odrv4 I__2392 (
            .O(N__18162),
            .I(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ));
    Odrv4 I__2391 (
            .O(N__18159),
            .I(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ));
    InMux I__2390 (
            .O(N__18154),
            .I(N__18151));
    LocalMux I__2389 (
            .O(N__18151),
            .I(\b2v_inst11.count_clk_0_6 ));
    InMux I__2388 (
            .O(N__18148),
            .I(N__18144));
    InMux I__2387 (
            .O(N__18147),
            .I(N__18141));
    LocalMux I__2386 (
            .O(N__18144),
            .I(N__18138));
    LocalMux I__2385 (
            .O(N__18141),
            .I(N__18135));
    Span4Mux_v I__2384 (
            .O(N__18138),
            .I(N__18132));
    Span4Mux_h I__2383 (
            .O(N__18135),
            .I(N__18129));
    Odrv4 I__2382 (
            .O(N__18132),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ));
    Odrv4 I__2381 (
            .O(N__18129),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ));
    InMux I__2380 (
            .O(N__18124),
            .I(N__18121));
    LocalMux I__2379 (
            .O(N__18121),
            .I(\b2v_inst11.count_clk_0_8 ));
    CEMux I__2378 (
            .O(N__18118),
            .I(N__18115));
    LocalMux I__2377 (
            .O(N__18115),
            .I(N__18108));
    CascadeMux I__2376 (
            .O(N__18114),
            .I(N__18103));
    CascadeMux I__2375 (
            .O(N__18113),
            .I(N__18099));
    CascadeMux I__2374 (
            .O(N__18112),
            .I(N__18096));
    CEMux I__2373 (
            .O(N__18111),
            .I(N__18092));
    Span4Mux_v I__2372 (
            .O(N__18108),
            .I(N__18088));
    CEMux I__2371 (
            .O(N__18107),
            .I(N__18085));
    InMux I__2370 (
            .O(N__18106),
            .I(N__18069));
    InMux I__2369 (
            .O(N__18103),
            .I(N__18069));
    InMux I__2368 (
            .O(N__18102),
            .I(N__18069));
    InMux I__2367 (
            .O(N__18099),
            .I(N__18069));
    InMux I__2366 (
            .O(N__18096),
            .I(N__18069));
    InMux I__2365 (
            .O(N__18095),
            .I(N__18069));
    LocalMux I__2364 (
            .O(N__18092),
            .I(N__18065));
    CEMux I__2363 (
            .O(N__18091),
            .I(N__18062));
    Span4Mux_h I__2362 (
            .O(N__18088),
            .I(N__18057));
    LocalMux I__2361 (
            .O(N__18085),
            .I(N__18057));
    CascadeMux I__2360 (
            .O(N__18084),
            .I(N__18051));
    InMux I__2359 (
            .O(N__18083),
            .I(N__18043));
    CEMux I__2358 (
            .O(N__18082),
            .I(N__18043));
    LocalMux I__2357 (
            .O(N__18069),
            .I(N__18040));
    CascadeMux I__2356 (
            .O(N__18068),
            .I(N__18037));
    Span4Mux_v I__2355 (
            .O(N__18065),
            .I(N__18034));
    LocalMux I__2354 (
            .O(N__18062),
            .I(N__18031));
    Span4Mux_s1_h I__2353 (
            .O(N__18057),
            .I(N__18028));
    InMux I__2352 (
            .O(N__18056),
            .I(N__18021));
    InMux I__2351 (
            .O(N__18055),
            .I(N__18021));
    InMux I__2350 (
            .O(N__18054),
            .I(N__18021));
    InMux I__2349 (
            .O(N__18051),
            .I(N__18018));
    InMux I__2348 (
            .O(N__18050),
            .I(N__18011));
    InMux I__2347 (
            .O(N__18049),
            .I(N__18011));
    InMux I__2346 (
            .O(N__18048),
            .I(N__18011));
    LocalMux I__2345 (
            .O(N__18043),
            .I(N__18006));
    Span4Mux_h I__2344 (
            .O(N__18040),
            .I(N__18006));
    InMux I__2343 (
            .O(N__18037),
            .I(N__18003));
    Odrv4 I__2342 (
            .O(N__18034),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__2341 (
            .O(N__18031),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__2340 (
            .O(N__18028),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2339 (
            .O(N__18021),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2338 (
            .O(N__18018),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2337 (
            .O(N__18011),
            .I(\b2v_inst11.count_clk_en ));
    Odrv4 I__2336 (
            .O(N__18006),
            .I(\b2v_inst11.count_clk_en ));
    LocalMux I__2335 (
            .O(N__18003),
            .I(\b2v_inst11.count_clk_en ));
    CascadeMux I__2334 (
            .O(N__17986),
            .I(N__17983));
    InMux I__2333 (
            .O(N__17983),
            .I(N__17980));
    LocalMux I__2332 (
            .O(N__17980),
            .I(N__17977));
    Span4Mux_v I__2331 (
            .O(N__17977),
            .I(N__17974));
    Odrv4 I__2330 (
            .O(N__17974),
            .I(func_state_RNIVS8U1_4_1));
    CascadeMux I__2329 (
            .O(N__17971),
            .I(N__17968));
    InMux I__2328 (
            .O(N__17968),
            .I(N__17962));
    InMux I__2327 (
            .O(N__17967),
            .I(N__17962));
    LocalMux I__2326 (
            .O(N__17962),
            .I(\b2v_inst11.func_stateZ0Z_1 ));
    InMux I__2325 (
            .O(N__17959),
            .I(N__17956));
    LocalMux I__2324 (
            .O(N__17956),
            .I(N__17952));
    CascadeMux I__2323 (
            .O(N__17955),
            .I(N__17949));
    Span4Mux_s3_h I__2322 (
            .O(N__17952),
            .I(N__17943));
    InMux I__2321 (
            .O(N__17949),
            .I(N__17938));
    InMux I__2320 (
            .O(N__17948),
            .I(N__17938));
    InMux I__2319 (
            .O(N__17947),
            .I(N__17933));
    InMux I__2318 (
            .O(N__17946),
            .I(N__17933));
    Odrv4 I__2317 (
            .O(N__17943),
            .I(\b2v_inst11.count_clk_enZ0Z_0 ));
    LocalMux I__2316 (
            .O(N__17938),
            .I(\b2v_inst11.count_clk_enZ0Z_0 ));
    LocalMux I__2315 (
            .O(N__17933),
            .I(\b2v_inst11.count_clk_enZ0Z_0 ));
    CascadeMux I__2314 (
            .O(N__17926),
            .I(VCCST_EN_i_0_o3_0_cascade_));
    InMux I__2313 (
            .O(N__17923),
            .I(N__17917));
    InMux I__2312 (
            .O(N__17922),
            .I(N__17917));
    LocalMux I__2311 (
            .O(N__17917),
            .I(\b2v_inst11.func_state_1_m2_1 ));
    CascadeMux I__2310 (
            .O(N__17914),
            .I(func_state_RNI6BE8E_0_1_cascade_));
    InMux I__2309 (
            .O(N__17911),
            .I(N__17908));
    LocalMux I__2308 (
            .O(N__17908),
            .I(\b2v_inst11.count_0_7 ));
    InMux I__2307 (
            .O(N__17905),
            .I(N__17900));
    InMux I__2306 (
            .O(N__17904),
            .I(N__17897));
    InMux I__2305 (
            .O(N__17903),
            .I(N__17894));
    LocalMux I__2304 (
            .O(N__17900),
            .I(N__17891));
    LocalMux I__2303 (
            .O(N__17897),
            .I(N__17886));
    LocalMux I__2302 (
            .O(N__17894),
            .I(N__17886));
    Span4Mux_h I__2301 (
            .O(N__17891),
            .I(N__17883));
    Span4Mux_s3_h I__2300 (
            .O(N__17886),
            .I(N__17880));
    Odrv4 I__2299 (
            .O(N__17883),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    Odrv4 I__2298 (
            .O(N__17880),
            .I(\b2v_inst11.count_clkZ0Z_3 ));
    InMux I__2297 (
            .O(N__17875),
            .I(N__17871));
    InMux I__2296 (
            .O(N__17874),
            .I(N__17867));
    LocalMux I__2295 (
            .O(N__17871),
            .I(N__17864));
    InMux I__2294 (
            .O(N__17870),
            .I(N__17861));
    LocalMux I__2293 (
            .O(N__17867),
            .I(N__17856));
    Span4Mux_s2_h I__2292 (
            .O(N__17864),
            .I(N__17856));
    LocalMux I__2291 (
            .O(N__17861),
            .I(N__17853));
    Span4Mux_v I__2290 (
            .O(N__17856),
            .I(N__17850));
    Span4Mux_s3_h I__2289 (
            .O(N__17853),
            .I(N__17847));
    Odrv4 I__2288 (
            .O(N__17850),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    Odrv4 I__2287 (
            .O(N__17847),
            .I(\b2v_inst11.count_clkZ0Z_6 ));
    InMux I__2286 (
            .O(N__17842),
            .I(N__17838));
    InMux I__2285 (
            .O(N__17841),
            .I(N__17835));
    LocalMux I__2284 (
            .O(N__17838),
            .I(N__17831));
    LocalMux I__2283 (
            .O(N__17835),
            .I(N__17828));
    InMux I__2282 (
            .O(N__17834),
            .I(N__17825));
    Span4Mux_h I__2281 (
            .O(N__17831),
            .I(N__17822));
    Span12Mux_s7_v I__2280 (
            .O(N__17828),
            .I(N__17819));
    LocalMux I__2279 (
            .O(N__17825),
            .I(N__17816));
    Odrv4 I__2278 (
            .O(N__17822),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    Odrv12 I__2277 (
            .O(N__17819),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    Odrv12 I__2276 (
            .O(N__17816),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1 ));
    CascadeMux I__2275 (
            .O(N__17809),
            .I(\b2v_inst11.func_state_1_m2_am_1_1_cascade_ ));
    InMux I__2274 (
            .O(N__17806),
            .I(N__17803));
    LocalMux I__2273 (
            .O(N__17803),
            .I(N__17800));
    Span4Mux_h I__2272 (
            .O(N__17800),
            .I(N__17794));
    InMux I__2271 (
            .O(N__17799),
            .I(N__17787));
    InMux I__2270 (
            .O(N__17798),
            .I(N__17787));
    InMux I__2269 (
            .O(N__17797),
            .I(N__17787));
    Odrv4 I__2268 (
            .O(N__17794),
            .I(\b2v_inst11.count_off_RNIZ0Z_9 ));
    LocalMux I__2267 (
            .O(N__17787),
            .I(\b2v_inst11.count_off_RNIZ0Z_9 ));
    CascadeMux I__2266 (
            .O(N__17782),
            .I(\b2v_inst11.func_state_RNIR5S85Z0Z_1_cascade_ ));
    CascadeMux I__2265 (
            .O(N__17779),
            .I(\b2v_inst11.func_state_cascade_ ));
    CascadeMux I__2264 (
            .O(N__17776),
            .I(N__17772));
    InMux I__2263 (
            .O(N__17775),
            .I(N__17767));
    InMux I__2262 (
            .O(N__17772),
            .I(N__17767));
    LocalMux I__2261 (
            .O(N__17767),
            .I(\b2v_inst11.func_stateZ0Z_0 ));
    InMux I__2260 (
            .O(N__17764),
            .I(N__17758));
    InMux I__2259 (
            .O(N__17763),
            .I(N__17758));
    LocalMux I__2258 (
            .O(N__17758),
            .I(N__17755));
    Odrv12 I__2257 (
            .O(N__17755),
            .I(\b2v_inst11.N_160_i ));
    CascadeMux I__2256 (
            .O(N__17752),
            .I(N__17747));
    CascadeMux I__2255 (
            .O(N__17751),
            .I(N__17742));
    InMux I__2254 (
            .O(N__17750),
            .I(N__17737));
    InMux I__2253 (
            .O(N__17747),
            .I(N__17731));
    InMux I__2252 (
            .O(N__17746),
            .I(N__17731));
    InMux I__2251 (
            .O(N__17745),
            .I(N__17728));
    InMux I__2250 (
            .O(N__17742),
            .I(N__17720));
    InMux I__2249 (
            .O(N__17741),
            .I(N__17720));
    InMux I__2248 (
            .O(N__17740),
            .I(N__17720));
    LocalMux I__2247 (
            .O(N__17737),
            .I(N__17717));
    InMux I__2246 (
            .O(N__17736),
            .I(N__17714));
    LocalMux I__2245 (
            .O(N__17731),
            .I(N__17711));
    LocalMux I__2244 (
            .O(N__17728),
            .I(N__17708));
    InMux I__2243 (
            .O(N__17727),
            .I(N__17705));
    LocalMux I__2242 (
            .O(N__17720),
            .I(N__17702));
    Span12Mux_s10_v I__2241 (
            .O(N__17717),
            .I(N__17699));
    LocalMux I__2240 (
            .O(N__17714),
            .I(N__17696));
    Span4Mux_s3_h I__2239 (
            .O(N__17711),
            .I(N__17693));
    Span4Mux_s3_h I__2238 (
            .O(N__17708),
            .I(N__17690));
    LocalMux I__2237 (
            .O(N__17705),
            .I(N__17685));
    Span4Mux_s3_h I__2236 (
            .O(N__17702),
            .I(N__17685));
    Odrv12 I__2235 (
            .O(N__17699),
            .I(\b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ));
    Odrv12 I__2234 (
            .O(N__17696),
            .I(\b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ));
    Odrv4 I__2233 (
            .O(N__17693),
            .I(\b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ));
    Odrv4 I__2232 (
            .O(N__17690),
            .I(\b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ));
    Odrv4 I__2231 (
            .O(N__17685),
            .I(\b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ));
    InMux I__2230 (
            .O(N__17674),
            .I(N__17671));
    LocalMux I__2229 (
            .O(N__17671),
            .I(N__17668));
    Odrv4 I__2228 (
            .O(N__17668),
            .I(\b2v_inst11.func_state_1_m0_0_1_0 ));
    CascadeMux I__2227 (
            .O(N__17665),
            .I(\b2v_inst11.func_state_1_m2_1_0_cascade_ ));
    CascadeMux I__2226 (
            .O(N__17662),
            .I(N__17658));
    InMux I__2225 (
            .O(N__17661),
            .I(N__17650));
    InMux I__2224 (
            .O(N__17658),
            .I(N__17650));
    InMux I__2223 (
            .O(N__17657),
            .I(N__17650));
    LocalMux I__2222 (
            .O(N__17650),
            .I(\b2v_inst11.N_76 ));
    InMux I__2221 (
            .O(N__17647),
            .I(N__17641));
    InMux I__2220 (
            .O(N__17646),
            .I(N__17641));
    LocalMux I__2219 (
            .O(N__17641),
            .I(\b2v_inst11.func_state_1_m2_0 ));
    CascadeMux I__2218 (
            .O(N__17638),
            .I(\b2v_inst11.func_state_RNI_2Z0Z_1_cascade_ ));
    InMux I__2217 (
            .O(N__17635),
            .I(N__17632));
    LocalMux I__2216 (
            .O(N__17632),
            .I(N__17629));
    Span4Mux_v I__2215 (
            .O(N__17629),
            .I(N__17626));
    Odrv4 I__2214 (
            .O(N__17626),
            .I(\b2v_inst11.N_337 ));
    CascadeMux I__2213 (
            .O(N__17623),
            .I(\b2v_inst11.func_state_1_m2s2_i_0_cascade_ ));
    InMux I__2212 (
            .O(N__17620),
            .I(N__17617));
    LocalMux I__2211 (
            .O(N__17617),
            .I(N__17614));
    Span4Mux_h I__2210 (
            .O(N__17614),
            .I(N__17611));
    Odrv4 I__2209 (
            .O(N__17611),
            .I(\b2v_inst11.N_338 ));
    CascadeMux I__2208 (
            .O(N__17608),
            .I(\b2v_inst11.dutycycle_RNI_5Z0Z_6_cascade_ ));
    InMux I__2207 (
            .O(N__17605),
            .I(N__17602));
    LocalMux I__2206 (
            .O(N__17602),
            .I(N__17599));
    Odrv4 I__2205 (
            .O(N__17599),
            .I(\b2v_inst11.N_231_N ));
    CascadeMux I__2204 (
            .O(N__17596),
            .I(\b2v_inst11.N_306_cascade_ ));
    CascadeMux I__2203 (
            .O(N__17593),
            .I(\b2v_inst11.N_354_cascade_ ));
    InMux I__2202 (
            .O(N__17590),
            .I(N__17587));
    LocalMux I__2201 (
            .O(N__17587),
            .I(N__17584));
    Odrv4 I__2200 (
            .O(N__17584),
            .I(b2v_inst11_g0_i_m2_i_a6_3_2));
    CascadeMux I__2199 (
            .O(N__17581),
            .I(\b2v_inst11.N_159_cascade_ ));
    CascadeMux I__2198 (
            .O(N__17578),
            .I(\b2v_inst11.func_state_1_m0_0_1_1_0_cascade_ ));
    InMux I__2197 (
            .O(N__17575),
            .I(N__17572));
    LocalMux I__2196 (
            .O(N__17572),
            .I(N__17569));
    Span4Mux_h I__2195 (
            .O(N__17569),
            .I(N__17566));
    Odrv4 I__2194 (
            .O(N__17566),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_313_N ));
    CascadeMux I__2193 (
            .O(N__17563),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_sx_cascade_ ));
    InMux I__2192 (
            .O(N__17560),
            .I(N__17557));
    LocalMux I__2191 (
            .O(N__17557),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1 ));
    InMux I__2190 (
            .O(N__17554),
            .I(N__17549));
    InMux I__2189 (
            .O(N__17553),
            .I(N__17544));
    InMux I__2188 (
            .O(N__17552),
            .I(N__17544));
    LocalMux I__2187 (
            .O(N__17549),
            .I(\b2v_inst11.dutycycleZ1Z_7 ));
    LocalMux I__2186 (
            .O(N__17544),
            .I(\b2v_inst11.dutycycleZ1Z_7 ));
    InMux I__2185 (
            .O(N__17539),
            .I(N__17535));
    InMux I__2184 (
            .O(N__17538),
            .I(N__17532));
    LocalMux I__2183 (
            .O(N__17535),
            .I(N__17527));
    LocalMux I__2182 (
            .O(N__17532),
            .I(N__17527));
    Odrv4 I__2181 (
            .O(N__17527),
            .I(\b2v_inst11.dutycycle_RNI24DD8Z0Z_7 ));
    CascadeMux I__2180 (
            .O(N__17524),
            .I(\b2v_inst11.dutycycle_RNIVGS13Z0Z_7_cascade_ ));
    CascadeMux I__2179 (
            .O(N__17521),
            .I(\b2v_inst11.N_160_i_cascade_ ));
    InMux I__2178 (
            .O(N__17518),
            .I(N__17515));
    LocalMux I__2177 (
            .O(N__17515),
            .I(N__17512));
    Odrv4 I__2176 (
            .O(N__17512),
            .I(\b2v_inst11.g1_0_sx ));
    CascadeMux I__2175 (
            .O(N__17509),
            .I(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_0_cascade_ ));
    InMux I__2174 (
            .O(N__17506),
            .I(N__17503));
    LocalMux I__2173 (
            .O(N__17503),
            .I(N__17500));
    Span4Mux_v I__2172 (
            .O(N__17500),
            .I(N__17497));
    Odrv4 I__2171 (
            .O(N__17497),
            .I(\b2v_inst11.func_state_RNI608H1_0Z0Z_1 ));
    InMux I__2170 (
            .O(N__17494),
            .I(N__17488));
    InMux I__2169 (
            .O(N__17493),
            .I(N__17488));
    LocalMux I__2168 (
            .O(N__17488),
            .I(N__17485));
    Odrv4 I__2167 (
            .O(N__17485),
            .I(\b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ));
    CascadeMux I__2166 (
            .O(N__17482),
            .I(N__17479));
    InMux I__2165 (
            .O(N__17479),
            .I(N__17476));
    LocalMux I__2164 (
            .O(N__17476),
            .I(\b2v_inst11.count_off_0_12 ));
    InMux I__2163 (
            .O(N__17473),
            .I(N__17469));
    InMux I__2162 (
            .O(N__17472),
            .I(N__17466));
    LocalMux I__2161 (
            .O(N__17469),
            .I(\b2v_inst11.count_offZ0Z_12 ));
    LocalMux I__2160 (
            .O(N__17466),
            .I(\b2v_inst11.count_offZ0Z_12 ));
    CascadeMux I__2159 (
            .O(N__17461),
            .I(N__17458));
    InMux I__2158 (
            .O(N__17458),
            .I(N__17455));
    LocalMux I__2157 (
            .O(N__17455),
            .I(N__17451));
    InMux I__2156 (
            .O(N__17454),
            .I(N__17448));
    Span4Mux_h I__2155 (
            .O(N__17451),
            .I(N__17445));
    LocalMux I__2154 (
            .O(N__17448),
            .I(N__17442));
    Odrv4 I__2153 (
            .O(N__17445),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    Odrv4 I__2152 (
            .O(N__17442),
            .I(\b2v_inst11.count_offZ0Z_10 ));
    InMux I__2151 (
            .O(N__17437),
            .I(N__17434));
    LocalMux I__2150 (
            .O(N__17434),
            .I(\b2v_inst11.un34_clk_100khz_5 ));
    CascadeMux I__2149 (
            .O(N__17431),
            .I(\b2v_inst11.un34_clk_100khz_4_cascade_ ));
    InMux I__2148 (
            .O(N__17428),
            .I(N__17425));
    LocalMux I__2147 (
            .O(N__17425),
            .I(N__17422));
    Odrv4 I__2146 (
            .O(N__17422),
            .I(\b2v_inst11.un34_clk_100khz_11 ));
    InMux I__2145 (
            .O(N__17419),
            .I(N__17413));
    InMux I__2144 (
            .O(N__17418),
            .I(N__17413));
    LocalMux I__2143 (
            .O(N__17413),
            .I(\b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ));
    InMux I__2142 (
            .O(N__17410),
            .I(N__17404));
    InMux I__2141 (
            .O(N__17409),
            .I(N__17404));
    LocalMux I__2140 (
            .O(N__17404),
            .I(\b2v_inst11.count_offZ0Z_11 ));
    CascadeMux I__2139 (
            .O(N__17401),
            .I(\b2v_inst11.g4_cascade_ ));
    CascadeMux I__2138 (
            .O(N__17398),
            .I(\b2v_inst11.g0_17_N_3L3_1_cascade_ ));
    InMux I__2137 (
            .O(N__17395),
            .I(N__17392));
    LocalMux I__2136 (
            .O(N__17392),
            .I(\b2v_inst11.dutycycle_RNIVGS13Z0Z_7 ));
    InMux I__2135 (
            .O(N__17389),
            .I(\b2v_inst11.un3_count_off_1_cry_11 ));
    InMux I__2134 (
            .O(N__17386),
            .I(N__17383));
    LocalMux I__2133 (
            .O(N__17383),
            .I(N__17380));
    Odrv4 I__2132 (
            .O(N__17380),
            .I(\b2v_inst11.count_offZ0Z_13 ));
    CascadeMux I__2131 (
            .O(N__17377),
            .I(N__17374));
    InMux I__2130 (
            .O(N__17374),
            .I(N__17370));
    InMux I__2129 (
            .O(N__17373),
            .I(N__17367));
    LocalMux I__2128 (
            .O(N__17370),
            .I(N__17364));
    LocalMux I__2127 (
            .O(N__17367),
            .I(N__17361));
    Odrv12 I__2126 (
            .O(N__17364),
            .I(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ));
    Odrv4 I__2125 (
            .O(N__17361),
            .I(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ));
    InMux I__2124 (
            .O(N__17356),
            .I(\b2v_inst11.un3_count_off_1_cry_12 ));
    InMux I__2123 (
            .O(N__17353),
            .I(\b2v_inst11.un3_count_off_1_cry_13 ));
    InMux I__2122 (
            .O(N__17350),
            .I(N__17347));
    LocalMux I__2121 (
            .O(N__17347),
            .I(N__17343));
    InMux I__2120 (
            .O(N__17346),
            .I(N__17340));
    Odrv4 I__2119 (
            .O(N__17343),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    LocalMux I__2118 (
            .O(N__17340),
            .I(\b2v_inst11.count_offZ0Z_15 ));
    InMux I__2117 (
            .O(N__17335),
            .I(\b2v_inst11.un3_count_off_1_cry_14 ));
    CascadeMux I__2116 (
            .O(N__17332),
            .I(N__17329));
    InMux I__2115 (
            .O(N__17329),
            .I(N__17323));
    InMux I__2114 (
            .O(N__17328),
            .I(N__17323));
    LocalMux I__2113 (
            .O(N__17323),
            .I(N__17320));
    Odrv4 I__2112 (
            .O(N__17320),
            .I(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ));
    InMux I__2111 (
            .O(N__17317),
            .I(N__17314));
    LocalMux I__2110 (
            .O(N__17314),
            .I(\b2v_inst11.un3_count_off_1_axb_11 ));
    InMux I__2109 (
            .O(N__17311),
            .I(N__17308));
    LocalMux I__2108 (
            .O(N__17308),
            .I(\b2v_inst11.count_off_1_11 ));
    CascadeMux I__2107 (
            .O(N__17305),
            .I(\b2v_inst11.count_off_1_11_cascade_ ));
    InMux I__2106 (
            .O(N__17302),
            .I(\b2v_inst11.un3_count_off_1_cry_3 ));
    InMux I__2105 (
            .O(N__17299),
            .I(\b2v_inst11.un3_count_off_1_cry_4 ));
    InMux I__2104 (
            .O(N__17296),
            .I(N__17293));
    LocalMux I__2103 (
            .O(N__17293),
            .I(N__17290));
    Span4Mux_h I__2102 (
            .O(N__17290),
            .I(N__17287));
    Span4Mux_v I__2101 (
            .O(N__17287),
            .I(N__17284));
    Odrv4 I__2100 (
            .O(N__17284),
            .I(\b2v_inst11.un3_count_off_1_axb_6 ));
    InMux I__2099 (
            .O(N__17281),
            .I(\b2v_inst11.un3_count_off_1_cry_5 ));
    CascadeMux I__2098 (
            .O(N__17278),
            .I(N__17275));
    InMux I__2097 (
            .O(N__17275),
            .I(N__17272));
    LocalMux I__2096 (
            .O(N__17272),
            .I(\b2v_inst11.un3_count_off_1_axb_7 ));
    InMux I__2095 (
            .O(N__17269),
            .I(\b2v_inst11.un3_count_off_1_cry_6 ));
    InMux I__2094 (
            .O(N__17266),
            .I(N__17263));
    LocalMux I__2093 (
            .O(N__17263),
            .I(\b2v_inst11.count_offZ0Z_8 ));
    CascadeMux I__2092 (
            .O(N__17260),
            .I(N__17257));
    InMux I__2091 (
            .O(N__17257),
            .I(N__17251));
    InMux I__2090 (
            .O(N__17256),
            .I(N__17251));
    LocalMux I__2089 (
            .O(N__17251),
            .I(\b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ));
    InMux I__2088 (
            .O(N__17248),
            .I(\b2v_inst11.un3_count_off_1_cry_7 ));
    InMux I__2087 (
            .O(N__17245),
            .I(bfn_4_5_0_));
    InMux I__2086 (
            .O(N__17242),
            .I(N__17238));
    InMux I__2085 (
            .O(N__17241),
            .I(N__17235));
    LocalMux I__2084 (
            .O(N__17238),
            .I(N__17230));
    LocalMux I__2083 (
            .O(N__17235),
            .I(N__17230));
    Odrv4 I__2082 (
            .O(N__17230),
            .I(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ));
    InMux I__2081 (
            .O(N__17227),
            .I(\b2v_inst11.un3_count_off_1_cry_9 ));
    InMux I__2080 (
            .O(N__17224),
            .I(\b2v_inst11.un3_count_off_1_cry_10 ));
    InMux I__2079 (
            .O(N__17221),
            .I(N__17218));
    LocalMux I__2078 (
            .O(N__17218),
            .I(\b2v_inst11.count_off_0_15 ));
    InMux I__2077 (
            .O(N__17215),
            .I(N__17212));
    LocalMux I__2076 (
            .O(N__17212),
            .I(N__17209));
    Span4Mux_h I__2075 (
            .O(N__17209),
            .I(N__17206));
    Odrv4 I__2074 (
            .O(N__17206),
            .I(\b2v_inst11.count_off_0_13 ));
    CascadeMux I__2073 (
            .O(N__17203),
            .I(\b2v_inst11.count_offZ0Z_13_cascade_ ));
    InMux I__2072 (
            .O(N__17200),
            .I(N__17197));
    LocalMux I__2071 (
            .O(N__17197),
            .I(\b2v_inst11.count_off_0_8 ));
    CascadeMux I__2070 (
            .O(N__17194),
            .I(\b2v_inst11.count_offZ0Z_8_cascade_ ));
    InMux I__2069 (
            .O(N__17191),
            .I(N__17187));
    CascadeMux I__2068 (
            .O(N__17190),
            .I(N__17184));
    LocalMux I__2067 (
            .O(N__17187),
            .I(N__17181));
    InMux I__2066 (
            .O(N__17184),
            .I(N__17178));
    Span4Mux_v I__2065 (
            .O(N__17181),
            .I(N__17175));
    LocalMux I__2064 (
            .O(N__17178),
            .I(N__17172));
    Span4Mux_v I__2063 (
            .O(N__17175),
            .I(N__17165));
    Span4Mux_v I__2062 (
            .O(N__17172),
            .I(N__17165));
    InMux I__2061 (
            .O(N__17171),
            .I(N__17160));
    InMux I__2060 (
            .O(N__17170),
            .I(N__17160));
    Odrv4 I__2059 (
            .O(N__17165),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    LocalMux I__2058 (
            .O(N__17160),
            .I(\b2v_inst11.count_offZ0Z_0 ));
    InMux I__2057 (
            .O(N__17155),
            .I(\b2v_inst11.un3_count_off_1_cry_1 ));
    InMux I__2056 (
            .O(N__17152),
            .I(\b2v_inst11.un3_count_off_1_cry_2 ));
    InMux I__2055 (
            .O(N__17149),
            .I(N__17146));
    LocalMux I__2054 (
            .O(N__17146),
            .I(\b2v_inst200.count_3_3 ));
    InMux I__2053 (
            .O(N__17143),
            .I(N__17140));
    LocalMux I__2052 (
            .O(N__17140),
            .I(N__17137));
    Odrv12 I__2051 (
            .O(N__17137),
            .I(\b2v_inst200.count_3_12 ));
    InMux I__2050 (
            .O(N__17134),
            .I(N__17131));
    LocalMux I__2049 (
            .O(N__17131),
            .I(\b2v_inst200.count_3_4 ));
    InMux I__2048 (
            .O(N__17128),
            .I(N__17125));
    LocalMux I__2047 (
            .O(N__17125),
            .I(N__17122));
    Odrv12 I__2046 (
            .O(N__17122),
            .I(\b2v_inst200.count_3_5 ));
    InMux I__2045 (
            .O(N__17119),
            .I(N__17116));
    LocalMux I__2044 (
            .O(N__17116),
            .I(N__17113));
    Odrv4 I__2043 (
            .O(N__17113),
            .I(\b2v_inst200.count_3_7 ));
    InMux I__2042 (
            .O(N__17110),
            .I(bfn_2_16_0_));
    InMux I__2041 (
            .O(N__17107),
            .I(N__17103));
    InMux I__2040 (
            .O(N__17106),
            .I(N__17100));
    LocalMux I__2039 (
            .O(N__17103),
            .I(\b2v_inst20.counterZ0Z_31 ));
    LocalMux I__2038 (
            .O(N__17100),
            .I(\b2v_inst20.counterZ0Z_31 ));
    InMux I__2037 (
            .O(N__17095),
            .I(N__17091));
    InMux I__2036 (
            .O(N__17094),
            .I(N__17088));
    LocalMux I__2035 (
            .O(N__17091),
            .I(\b2v_inst20.counterZ0Z_29 ));
    LocalMux I__2034 (
            .O(N__17088),
            .I(\b2v_inst20.counterZ0Z_29 ));
    CascadeMux I__2033 (
            .O(N__17083),
            .I(N__17079));
    InMux I__2032 (
            .O(N__17082),
            .I(N__17076));
    InMux I__2031 (
            .O(N__17079),
            .I(N__17073));
    LocalMux I__2030 (
            .O(N__17076),
            .I(\b2v_inst20.counterZ0Z_30 ));
    LocalMux I__2029 (
            .O(N__17073),
            .I(\b2v_inst20.counterZ0Z_30 ));
    InMux I__2028 (
            .O(N__17068),
            .I(N__17064));
    InMux I__2027 (
            .O(N__17067),
            .I(N__17061));
    LocalMux I__2026 (
            .O(N__17064),
            .I(\b2v_inst20.counterZ0Z_28 ));
    LocalMux I__2025 (
            .O(N__17061),
            .I(\b2v_inst20.counterZ0Z_28 ));
    InMux I__2024 (
            .O(N__17056),
            .I(N__17053));
    LocalMux I__2023 (
            .O(N__17053),
            .I(\b2v_inst20.un4_counter_7_and ));
    InMux I__2022 (
            .O(N__17050),
            .I(N__17046));
    InMux I__2021 (
            .O(N__17049),
            .I(N__17043));
    LocalMux I__2020 (
            .O(N__17046),
            .I(\b2v_inst20.counterZ0Z_27 ));
    LocalMux I__2019 (
            .O(N__17043),
            .I(\b2v_inst20.counterZ0Z_27 ));
    InMux I__2018 (
            .O(N__17038),
            .I(N__17034));
    InMux I__2017 (
            .O(N__17037),
            .I(N__17031));
    LocalMux I__2016 (
            .O(N__17034),
            .I(\b2v_inst20.counterZ0Z_25 ));
    LocalMux I__2015 (
            .O(N__17031),
            .I(\b2v_inst20.counterZ0Z_25 ));
    CascadeMux I__2014 (
            .O(N__17026),
            .I(N__17022));
    InMux I__2013 (
            .O(N__17025),
            .I(N__17019));
    InMux I__2012 (
            .O(N__17022),
            .I(N__17016));
    LocalMux I__2011 (
            .O(N__17019),
            .I(\b2v_inst20.counterZ0Z_26 ));
    LocalMux I__2010 (
            .O(N__17016),
            .I(\b2v_inst20.counterZ0Z_26 ));
    InMux I__2009 (
            .O(N__17011),
            .I(N__17007));
    InMux I__2008 (
            .O(N__17010),
            .I(N__17004));
    LocalMux I__2007 (
            .O(N__17007),
            .I(\b2v_inst20.counterZ0Z_24 ));
    LocalMux I__2006 (
            .O(N__17004),
            .I(\b2v_inst20.counterZ0Z_24 ));
    InMux I__2005 (
            .O(N__16999),
            .I(N__16996));
    LocalMux I__2004 (
            .O(N__16996),
            .I(\b2v_inst20.un4_counter_6_and ));
    InMux I__2003 (
            .O(N__16993),
            .I(N__16990));
    LocalMux I__2002 (
            .O(N__16990),
            .I(\b2v_inst200.count_3_1 ));
    InMux I__2001 (
            .O(N__16987),
            .I(N__16984));
    LocalMux I__2000 (
            .O(N__16984),
            .I(\b2v_inst200.count_3_2 ));
    InMux I__1999 (
            .O(N__16981),
            .I(N__16978));
    LocalMux I__1998 (
            .O(N__16978),
            .I(N__16975));
    IoSpan4Mux I__1997 (
            .O(N__16975),
            .I(N__16972));
    IoSpan4Mux I__1996 (
            .O(N__16972),
            .I(N__16969));
    Odrv4 I__1995 (
            .O(N__16969),
            .I(VPP_OK_c));
    IoInMux I__1994 (
            .O(N__16966),
            .I(N__16963));
    LocalMux I__1993 (
            .O(N__16963),
            .I(N__16960));
    Odrv12 I__1992 (
            .O(N__16960),
            .I(VDDQ_EN_c));
    CascadeMux I__1991 (
            .O(N__16957),
            .I(N__16954));
    InMux I__1990 (
            .O(N__16954),
            .I(N__16951));
    LocalMux I__1989 (
            .O(N__16951),
            .I(\b2v_inst20.un4_counter_2_and ));
    CascadeMux I__1988 (
            .O(N__16948),
            .I(N__16945));
    InMux I__1987 (
            .O(N__16945),
            .I(N__16942));
    LocalMux I__1986 (
            .O(N__16942),
            .I(\b2v_inst20.un4_counter_3_and ));
    InMux I__1985 (
            .O(N__16939),
            .I(N__16936));
    LocalMux I__1984 (
            .O(N__16936),
            .I(\b2v_inst20.un4_counter_4_and ));
    InMux I__1983 (
            .O(N__16933),
            .I(N__16930));
    LocalMux I__1982 (
            .O(N__16930),
            .I(\b2v_inst20.un4_counter_5_and ));
    InMux I__1981 (
            .O(N__16927),
            .I(N__16923));
    InMux I__1980 (
            .O(N__16926),
            .I(N__16920));
    LocalMux I__1979 (
            .O(N__16923),
            .I(N__16917));
    LocalMux I__1978 (
            .O(N__16920),
            .I(N__16914));
    Span4Mux_s1_h I__1977 (
            .O(N__16917),
            .I(N__16911));
    Odrv4 I__1976 (
            .O(N__16914),
            .I(\b2v_inst11.count_clk_1_14 ));
    Odrv4 I__1975 (
            .O(N__16911),
            .I(\b2v_inst11.count_clk_1_14 ));
    InMux I__1974 (
            .O(N__16906),
            .I(\b2v_inst11.un1_count_clk_2_cry_13 ));
    InMux I__1973 (
            .O(N__16903),
            .I(N__16900));
    LocalMux I__1972 (
            .O(N__16900),
            .I(N__16896));
    InMux I__1971 (
            .O(N__16899),
            .I(N__16893));
    Odrv4 I__1970 (
            .O(N__16896),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    LocalMux I__1969 (
            .O(N__16893),
            .I(\b2v_inst11.count_clkZ0Z_15 ));
    CascadeMux I__1968 (
            .O(N__16888),
            .I(N__16881));
    InMux I__1967 (
            .O(N__16887),
            .I(N__16862));
    InMux I__1966 (
            .O(N__16886),
            .I(N__16859));
    InMux I__1965 (
            .O(N__16885),
            .I(N__16852));
    InMux I__1964 (
            .O(N__16884),
            .I(N__16852));
    InMux I__1963 (
            .O(N__16881),
            .I(N__16852));
    InMux I__1962 (
            .O(N__16880),
            .I(N__16845));
    InMux I__1961 (
            .O(N__16879),
            .I(N__16845));
    InMux I__1960 (
            .O(N__16878),
            .I(N__16845));
    InMux I__1959 (
            .O(N__16877),
            .I(N__16838));
    InMux I__1958 (
            .O(N__16876),
            .I(N__16838));
    InMux I__1957 (
            .O(N__16875),
            .I(N__16838));
    InMux I__1956 (
            .O(N__16874),
            .I(N__16831));
    InMux I__1955 (
            .O(N__16873),
            .I(N__16831));
    InMux I__1954 (
            .O(N__16872),
            .I(N__16831));
    InMux I__1953 (
            .O(N__16871),
            .I(N__16816));
    InMux I__1952 (
            .O(N__16870),
            .I(N__16816));
    InMux I__1951 (
            .O(N__16869),
            .I(N__16816));
    InMux I__1950 (
            .O(N__16868),
            .I(N__16816));
    InMux I__1949 (
            .O(N__16867),
            .I(N__16816));
    InMux I__1948 (
            .O(N__16866),
            .I(N__16816));
    InMux I__1947 (
            .O(N__16865),
            .I(N__16816));
    LocalMux I__1946 (
            .O(N__16862),
            .I(N__16809));
    LocalMux I__1945 (
            .O(N__16859),
            .I(N__16809));
    LocalMux I__1944 (
            .O(N__16852),
            .I(N__16809));
    LocalMux I__1943 (
            .O(N__16845),
            .I(\b2v_inst11.func_state_RNICGI84_0_0 ));
    LocalMux I__1942 (
            .O(N__16838),
            .I(\b2v_inst11.func_state_RNICGI84_0_0 ));
    LocalMux I__1941 (
            .O(N__16831),
            .I(\b2v_inst11.func_state_RNICGI84_0_0 ));
    LocalMux I__1940 (
            .O(N__16816),
            .I(\b2v_inst11.func_state_RNICGI84_0_0 ));
    Odrv4 I__1939 (
            .O(N__16809),
            .I(\b2v_inst11.func_state_RNICGI84_0_0 ));
    InMux I__1938 (
            .O(N__16798),
            .I(\b2v_inst11.un1_count_clk_2_cry_14 ));
    CascadeMux I__1937 (
            .O(N__16795),
            .I(N__16791));
    InMux I__1936 (
            .O(N__16794),
            .I(N__16786));
    InMux I__1935 (
            .O(N__16791),
            .I(N__16786));
    LocalMux I__1934 (
            .O(N__16786),
            .I(N__16783));
    Odrv4 I__1933 (
            .O(N__16783),
            .I(\b2v_inst11.count_clk_1_15 ));
    InMux I__1932 (
            .O(N__16780),
            .I(N__16776));
    InMux I__1931 (
            .O(N__16779),
            .I(N__16773));
    LocalMux I__1930 (
            .O(N__16776),
            .I(\b2v_inst20.counterZ0Z_11 ));
    LocalMux I__1929 (
            .O(N__16773),
            .I(\b2v_inst20.counterZ0Z_11 ));
    InMux I__1928 (
            .O(N__16768),
            .I(N__16764));
    InMux I__1927 (
            .O(N__16767),
            .I(N__16761));
    LocalMux I__1926 (
            .O(N__16764),
            .I(\b2v_inst20.counterZ0Z_9 ));
    LocalMux I__1925 (
            .O(N__16761),
            .I(\b2v_inst20.counterZ0Z_9 ));
    CascadeMux I__1924 (
            .O(N__16756),
            .I(N__16752));
    InMux I__1923 (
            .O(N__16755),
            .I(N__16749));
    InMux I__1922 (
            .O(N__16752),
            .I(N__16746));
    LocalMux I__1921 (
            .O(N__16749),
            .I(\b2v_inst20.counterZ0Z_10 ));
    LocalMux I__1920 (
            .O(N__16746),
            .I(\b2v_inst20.counterZ0Z_10 ));
    InMux I__1919 (
            .O(N__16741),
            .I(N__16737));
    InMux I__1918 (
            .O(N__16740),
            .I(N__16734));
    LocalMux I__1917 (
            .O(N__16737),
            .I(\b2v_inst20.counterZ0Z_8 ));
    LocalMux I__1916 (
            .O(N__16734),
            .I(\b2v_inst20.counterZ0Z_8 ));
    InMux I__1915 (
            .O(N__16729),
            .I(N__16725));
    InMux I__1914 (
            .O(N__16728),
            .I(N__16722));
    LocalMux I__1913 (
            .O(N__16725),
            .I(\b2v_inst20.counterZ0Z_15 ));
    LocalMux I__1912 (
            .O(N__16722),
            .I(\b2v_inst20.counterZ0Z_15 ));
    InMux I__1911 (
            .O(N__16717),
            .I(N__16713));
    InMux I__1910 (
            .O(N__16716),
            .I(N__16710));
    LocalMux I__1909 (
            .O(N__16713),
            .I(\b2v_inst20.counterZ0Z_14 ));
    LocalMux I__1908 (
            .O(N__16710),
            .I(\b2v_inst20.counterZ0Z_14 ));
    CascadeMux I__1907 (
            .O(N__16705),
            .I(N__16701));
    InMux I__1906 (
            .O(N__16704),
            .I(N__16698));
    InMux I__1905 (
            .O(N__16701),
            .I(N__16695));
    LocalMux I__1904 (
            .O(N__16698),
            .I(\b2v_inst20.counterZ0Z_13 ));
    LocalMux I__1903 (
            .O(N__16695),
            .I(\b2v_inst20.counterZ0Z_13 ));
    InMux I__1902 (
            .O(N__16690),
            .I(N__16686));
    InMux I__1901 (
            .O(N__16689),
            .I(N__16683));
    LocalMux I__1900 (
            .O(N__16686),
            .I(\b2v_inst20.counterZ0Z_12 ));
    LocalMux I__1899 (
            .O(N__16683),
            .I(\b2v_inst20.counterZ0Z_12 ));
    InMux I__1898 (
            .O(N__16678),
            .I(N__16674));
    InMux I__1897 (
            .O(N__16677),
            .I(N__16671));
    LocalMux I__1896 (
            .O(N__16674),
            .I(\b2v_inst20.counterZ0Z_19 ));
    LocalMux I__1895 (
            .O(N__16671),
            .I(\b2v_inst20.counterZ0Z_19 ));
    InMux I__1894 (
            .O(N__16666),
            .I(N__16662));
    InMux I__1893 (
            .O(N__16665),
            .I(N__16659));
    LocalMux I__1892 (
            .O(N__16662),
            .I(\b2v_inst20.counterZ0Z_17 ));
    LocalMux I__1891 (
            .O(N__16659),
            .I(\b2v_inst20.counterZ0Z_17 ));
    CascadeMux I__1890 (
            .O(N__16654),
            .I(N__16650));
    InMux I__1889 (
            .O(N__16653),
            .I(N__16647));
    InMux I__1888 (
            .O(N__16650),
            .I(N__16644));
    LocalMux I__1887 (
            .O(N__16647),
            .I(\b2v_inst20.counterZ0Z_18 ));
    LocalMux I__1886 (
            .O(N__16644),
            .I(\b2v_inst20.counterZ0Z_18 ));
    InMux I__1885 (
            .O(N__16639),
            .I(N__16635));
    InMux I__1884 (
            .O(N__16638),
            .I(N__16632));
    LocalMux I__1883 (
            .O(N__16635),
            .I(\b2v_inst20.counterZ0Z_16 ));
    LocalMux I__1882 (
            .O(N__16632),
            .I(\b2v_inst20.counterZ0Z_16 ));
    InMux I__1881 (
            .O(N__16627),
            .I(N__16623));
    InMux I__1880 (
            .O(N__16626),
            .I(N__16620));
    LocalMux I__1879 (
            .O(N__16623),
            .I(\b2v_inst20.counterZ0Z_23 ));
    LocalMux I__1878 (
            .O(N__16620),
            .I(\b2v_inst20.counterZ0Z_23 ));
    InMux I__1877 (
            .O(N__16615),
            .I(N__16611));
    InMux I__1876 (
            .O(N__16614),
            .I(N__16608));
    LocalMux I__1875 (
            .O(N__16611),
            .I(\b2v_inst20.counterZ0Z_21 ));
    LocalMux I__1874 (
            .O(N__16608),
            .I(\b2v_inst20.counterZ0Z_21 ));
    CascadeMux I__1873 (
            .O(N__16603),
            .I(N__16599));
    InMux I__1872 (
            .O(N__16602),
            .I(N__16596));
    InMux I__1871 (
            .O(N__16599),
            .I(N__16593));
    LocalMux I__1870 (
            .O(N__16596),
            .I(\b2v_inst20.counterZ0Z_22 ));
    LocalMux I__1869 (
            .O(N__16593),
            .I(\b2v_inst20.counterZ0Z_22 ));
    InMux I__1868 (
            .O(N__16588),
            .I(N__16584));
    InMux I__1867 (
            .O(N__16587),
            .I(N__16581));
    LocalMux I__1866 (
            .O(N__16584),
            .I(\b2v_inst20.counterZ0Z_20 ));
    LocalMux I__1865 (
            .O(N__16581),
            .I(\b2v_inst20.counterZ0Z_20 ));
    InMux I__1864 (
            .O(N__16576),
            .I(\b2v_inst11.un1_count_clk_2_cry_5 ));
    InMux I__1863 (
            .O(N__16573),
            .I(N__16569));
    InMux I__1862 (
            .O(N__16572),
            .I(N__16563));
    LocalMux I__1861 (
            .O(N__16569),
            .I(N__16560));
    InMux I__1860 (
            .O(N__16568),
            .I(N__16555));
    InMux I__1859 (
            .O(N__16567),
            .I(N__16555));
    InMux I__1858 (
            .O(N__16566),
            .I(N__16552));
    LocalMux I__1857 (
            .O(N__16563),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    Odrv12 I__1856 (
            .O(N__16560),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    LocalMux I__1855 (
            .O(N__16555),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    LocalMux I__1854 (
            .O(N__16552),
            .I(\b2v_inst11.count_clkZ0Z_7 ));
    InMux I__1853 (
            .O(N__16543),
            .I(N__16537));
    InMux I__1852 (
            .O(N__16542),
            .I(N__16537));
    LocalMux I__1851 (
            .O(N__16537),
            .I(N__16534));
    Odrv4 I__1850 (
            .O(N__16534),
            .I(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ));
    InMux I__1849 (
            .O(N__16531),
            .I(\b2v_inst11.un1_count_clk_2_cry_6 ));
    InMux I__1848 (
            .O(N__16528),
            .I(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__1847 (
            .O(N__16525),
            .I(bfn_2_13_0_));
    InMux I__1846 (
            .O(N__16522),
            .I(N__16519));
    LocalMux I__1845 (
            .O(N__16519),
            .I(\b2v_inst11.count_clkZ0Z_10 ));
    CascadeMux I__1844 (
            .O(N__16516),
            .I(N__16513));
    InMux I__1843 (
            .O(N__16513),
            .I(N__16507));
    InMux I__1842 (
            .O(N__16512),
            .I(N__16507));
    LocalMux I__1841 (
            .O(N__16507),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ));
    InMux I__1840 (
            .O(N__16504),
            .I(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ));
    InMux I__1839 (
            .O(N__16501),
            .I(N__16497));
    InMux I__1838 (
            .O(N__16500),
            .I(N__16494));
    LocalMux I__1837 (
            .O(N__16497),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    LocalMux I__1836 (
            .O(N__16494),
            .I(\b2v_inst11.count_clkZ0Z_11 ));
    CascadeMux I__1835 (
            .O(N__16489),
            .I(N__16486));
    InMux I__1834 (
            .O(N__16486),
            .I(N__16480));
    InMux I__1833 (
            .O(N__16485),
            .I(N__16480));
    LocalMux I__1832 (
            .O(N__16480),
            .I(\b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0 ));
    InMux I__1831 (
            .O(N__16477),
            .I(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ));
    InMux I__1830 (
            .O(N__16474),
            .I(N__16470));
    InMux I__1829 (
            .O(N__16473),
            .I(N__16467));
    LocalMux I__1828 (
            .O(N__16470),
            .I(\b2v_inst11.count_clkZ0Z_12 ));
    LocalMux I__1827 (
            .O(N__16467),
            .I(\b2v_inst11.count_clkZ0Z_12 ));
    InMux I__1826 (
            .O(N__16462),
            .I(N__16456));
    InMux I__1825 (
            .O(N__16461),
            .I(N__16456));
    LocalMux I__1824 (
            .O(N__16456),
            .I(\b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0 ));
    InMux I__1823 (
            .O(N__16453),
            .I(\b2v_inst11.un1_count_clk_2_cry_11 ));
    InMux I__1822 (
            .O(N__16450),
            .I(N__16446));
    CascadeMux I__1821 (
            .O(N__16449),
            .I(N__16442));
    LocalMux I__1820 (
            .O(N__16446),
            .I(N__16439));
    InMux I__1819 (
            .O(N__16445),
            .I(N__16434));
    InMux I__1818 (
            .O(N__16442),
            .I(N__16434));
    Odrv4 I__1817 (
            .O(N__16439),
            .I(\b2v_inst11.count_clkZ0Z_13 ));
    LocalMux I__1816 (
            .O(N__16434),
            .I(\b2v_inst11.count_clkZ0Z_13 ));
    InMux I__1815 (
            .O(N__16429),
            .I(N__16423));
    InMux I__1814 (
            .O(N__16428),
            .I(N__16423));
    LocalMux I__1813 (
            .O(N__16423),
            .I(N__16420));
    Span4Mux_s1_h I__1812 (
            .O(N__16420),
            .I(N__16417));
    Odrv4 I__1811 (
            .O(N__16417),
            .I(\b2v_inst11.count_clk_1_13 ));
    InMux I__1810 (
            .O(N__16414),
            .I(\b2v_inst11.un1_count_clk_2_cry_12 ));
    InMux I__1809 (
            .O(N__16411),
            .I(N__16408));
    LocalMux I__1808 (
            .O(N__16408),
            .I(N__16403));
    InMux I__1807 (
            .O(N__16407),
            .I(N__16398));
    InMux I__1806 (
            .O(N__16406),
            .I(N__16398));
    Odrv4 I__1805 (
            .O(N__16403),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    LocalMux I__1804 (
            .O(N__16398),
            .I(\b2v_inst11.count_clkZ0Z_14 ));
    InMux I__1803 (
            .O(N__16393),
            .I(N__16390));
    LocalMux I__1802 (
            .O(N__16390),
            .I(\b2v_inst11.count_clk_0_14 ));
    InMux I__1801 (
            .O(N__16387),
            .I(N__16384));
    LocalMux I__1800 (
            .O(N__16384),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_2 ));
    InMux I__1799 (
            .O(N__16381),
            .I(N__16378));
    LocalMux I__1798 (
            .O(N__16378),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_3 ));
    InMux I__1797 (
            .O(N__16375),
            .I(N__16371));
    InMux I__1796 (
            .O(N__16374),
            .I(N__16365));
    LocalMux I__1795 (
            .O(N__16371),
            .I(N__16362));
    InMux I__1794 (
            .O(N__16370),
            .I(N__16359));
    InMux I__1793 (
            .O(N__16369),
            .I(N__16356));
    InMux I__1792 (
            .O(N__16368),
            .I(N__16353));
    LocalMux I__1791 (
            .O(N__16365),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    Odrv4 I__1790 (
            .O(N__16362),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    LocalMux I__1789 (
            .O(N__16359),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    LocalMux I__1788 (
            .O(N__16356),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    LocalMux I__1787 (
            .O(N__16353),
            .I(\b2v_inst11.count_clkZ0Z_1 ));
    CascadeMux I__1786 (
            .O(N__16342),
            .I(N__16338));
    InMux I__1785 (
            .O(N__16341),
            .I(N__16331));
    InMux I__1784 (
            .O(N__16338),
            .I(N__16327));
    InMux I__1783 (
            .O(N__16337),
            .I(N__16324));
    InMux I__1782 (
            .O(N__16336),
            .I(N__16317));
    InMux I__1781 (
            .O(N__16335),
            .I(N__16317));
    InMux I__1780 (
            .O(N__16334),
            .I(N__16317));
    LocalMux I__1779 (
            .O(N__16331),
            .I(N__16314));
    InMux I__1778 (
            .O(N__16330),
            .I(N__16311));
    LocalMux I__1777 (
            .O(N__16327),
            .I(N__16308));
    LocalMux I__1776 (
            .O(N__16324),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    LocalMux I__1775 (
            .O(N__16317),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    Odrv4 I__1774 (
            .O(N__16314),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    LocalMux I__1773 (
            .O(N__16311),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    Odrv4 I__1772 (
            .O(N__16308),
            .I(\b2v_inst11.count_clkZ0Z_0 ));
    InMux I__1771 (
            .O(N__16297),
            .I(\b2v_inst11.un1_count_clk_2_cry_1 ));
    InMux I__1770 (
            .O(N__16294),
            .I(\b2v_inst11.un1_count_clk_2_cry_2 ));
    InMux I__1769 (
            .O(N__16291),
            .I(N__16288));
    LocalMux I__1768 (
            .O(N__16288),
            .I(N__16283));
    InMux I__1767 (
            .O(N__16287),
            .I(N__16278));
    InMux I__1766 (
            .O(N__16286),
            .I(N__16278));
    Odrv4 I__1765 (
            .O(N__16283),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    LocalMux I__1764 (
            .O(N__16278),
            .I(\b2v_inst11.count_clkZ0Z_4 ));
    InMux I__1763 (
            .O(N__16273),
            .I(N__16270));
    LocalMux I__1762 (
            .O(N__16270),
            .I(N__16267));
    Span4Mux_v I__1761 (
            .O(N__16267),
            .I(N__16263));
    InMux I__1760 (
            .O(N__16266),
            .I(N__16260));
    Span4Mux_v I__1759 (
            .O(N__16263),
            .I(N__16255));
    LocalMux I__1758 (
            .O(N__16260),
            .I(N__16255));
    Odrv4 I__1757 (
            .O(N__16255),
            .I(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ));
    InMux I__1756 (
            .O(N__16252),
            .I(\b2v_inst11.un1_count_clk_2_cry_3 ));
    InMux I__1755 (
            .O(N__16249),
            .I(\b2v_inst11.un1_count_clk_2_cry_4 ));
    InMux I__1754 (
            .O(N__16246),
            .I(N__16243));
    LocalMux I__1753 (
            .O(N__16243),
            .I(\b2v_inst11.count_clk_0_0 ));
    InMux I__1752 (
            .O(N__16240),
            .I(N__16237));
    LocalMux I__1751 (
            .O(N__16237),
            .I(\b2v_inst11.count_clk_0_7 ));
    CascadeMux I__1750 (
            .O(N__16234),
            .I(\b2v_inst11.N_168_cascade_ ));
    CascadeMux I__1749 (
            .O(N__16231),
            .I(\b2v_inst11.func_state_RNICGI84_0_0_cascade_ ));
    InMux I__1748 (
            .O(N__16228),
            .I(N__16225));
    LocalMux I__1747 (
            .O(N__16225),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_0 ));
    CascadeMux I__1746 (
            .O(N__16222),
            .I(N__16219));
    InMux I__1745 (
            .O(N__16219),
            .I(N__16216));
    LocalMux I__1744 (
            .O(N__16216),
            .I(\b2v_inst11.func_state_RNIVS8U1_0Z0Z_0 ));
    InMux I__1743 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__1742 (
            .O(N__16210),
            .I(N__16207));
    Odrv4 I__1741 (
            .O(N__16207),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1 ));
    InMux I__1740 (
            .O(N__16204),
            .I(N__16201));
    LocalMux I__1739 (
            .O(N__16201),
            .I(N__16198));
    Odrv12 I__1738 (
            .O(N__16198),
            .I(\b2v_inst11.N_340 ));
    InMux I__1737 (
            .O(N__16195),
            .I(N__16192));
    LocalMux I__1736 (
            .O(N__16192),
            .I(\b2v_inst11.func_state_1_ss0_i_0_o3_1 ));
    InMux I__1735 (
            .O(N__16189),
            .I(N__16184));
    InMux I__1734 (
            .O(N__16188),
            .I(N__16179));
    InMux I__1733 (
            .O(N__16187),
            .I(N__16179));
    LocalMux I__1732 (
            .O(N__16184),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    LocalMux I__1731 (
            .O(N__16179),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_1 ));
    InMux I__1730 (
            .O(N__16174),
            .I(N__16171));
    LocalMux I__1729 (
            .O(N__16171),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz ));
    CascadeMux I__1728 (
            .O(N__16168),
            .I(\b2v_inst11.count_off_RNIZ0Z_9_cascade_ ));
    CascadeMux I__1727 (
            .O(N__16165),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_1_cascade_ ));
    InMux I__1726 (
            .O(N__16162),
            .I(N__16159));
    LocalMux I__1725 (
            .O(N__16159),
            .I(\b2v_inst11.un1_func_state25_4_i_a3_0_1 ));
    CascadeMux I__1724 (
            .O(N__16156),
            .I(\b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ));
    CascadeMux I__1723 (
            .O(N__16153),
            .I(\b2v_inst11.count_clkZ0Z_1_cascade_ ));
    InMux I__1722 (
            .O(N__16150),
            .I(N__16147));
    LocalMux I__1721 (
            .O(N__16147),
            .I(\b2v_inst11.count_clk_0_1 ));
    CascadeMux I__1720 (
            .O(N__16144),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_ ));
    CascadeMux I__1719 (
            .O(N__16141),
            .I(N__16138));
    InMux I__1718 (
            .O(N__16138),
            .I(N__16135));
    LocalMux I__1717 (
            .O(N__16135),
            .I(N__16131));
    InMux I__1716 (
            .O(N__16134),
            .I(N__16128));
    Odrv4 I__1715 (
            .O(N__16131),
            .I(\b2v_inst11.count_clk_RNIVS8U1Z0Z_13 ));
    LocalMux I__1714 (
            .O(N__16128),
            .I(\b2v_inst11.count_clk_RNIVS8U1Z0Z_13 ));
    InMux I__1713 (
            .O(N__16123),
            .I(N__16120));
    LocalMux I__1712 (
            .O(N__16120),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_329_N ));
    CascadeMux I__1711 (
            .O(N__16117),
            .I(\b2v_inst11.un1_func_state25_6_0_1_cascade_ ));
    InMux I__1710 (
            .O(N__16114),
            .I(N__16110));
    InMux I__1709 (
            .O(N__16113),
            .I(N__16107));
    LocalMux I__1708 (
            .O(N__16110),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_0 ));
    LocalMux I__1707 (
            .O(N__16107),
            .I(\b2v_inst11.func_state_RNI_1Z0Z_0 ));
    InMux I__1706 (
            .O(N__16102),
            .I(N__16099));
    LocalMux I__1705 (
            .O(N__16099),
            .I(N__16096));
    Span4Mux_s1_h I__1704 (
            .O(N__16096),
            .I(N__16093));
    Odrv4 I__1703 (
            .O(N__16093),
            .I(N_236_0));
    InMux I__1702 (
            .O(N__16090),
            .I(N__16087));
    LocalMux I__1701 (
            .O(N__16087),
            .I(\b2v_inst11.g1_0_0_1 ));
    InMux I__1700 (
            .O(N__16084),
            .I(N__16081));
    LocalMux I__1699 (
            .O(N__16081),
            .I(\b2v_inst11.un1_func_state25_6_0_o_N_331_N ));
    InMux I__1698 (
            .O(N__16078),
            .I(N__16075));
    LocalMux I__1697 (
            .O(N__16075),
            .I(N__16072));
    Odrv4 I__1696 (
            .O(N__16072),
            .I(\b2v_inst11.count_clk_en_1 ));
    CascadeMux I__1695 (
            .O(N__16069),
            .I(N__16066));
    InMux I__1694 (
            .O(N__16066),
            .I(N__16063));
    LocalMux I__1693 (
            .O(N__16063),
            .I(\b2v_inst11.N_328 ));
    CascadeMux I__1692 (
            .O(N__16060),
            .I(\b2v_inst16.N_268_cascade_ ));
    InMux I__1691 (
            .O(N__16057),
            .I(N__16046));
    InMux I__1690 (
            .O(N__16056),
            .I(N__16046));
    InMux I__1689 (
            .O(N__16055),
            .I(N__16046));
    CascadeMux I__1688 (
            .O(N__16054),
            .I(N__16040));
    CascadeMux I__1687 (
            .O(N__16053),
            .I(N__16031));
    LocalMux I__1686 (
            .O(N__16046),
            .I(N__16020));
    InMux I__1685 (
            .O(N__16045),
            .I(N__16009));
    InMux I__1684 (
            .O(N__16044),
            .I(N__16009));
    InMux I__1683 (
            .O(N__16043),
            .I(N__16009));
    InMux I__1682 (
            .O(N__16040),
            .I(N__16009));
    InMux I__1681 (
            .O(N__16039),
            .I(N__16009));
    InMux I__1680 (
            .O(N__16038),
            .I(N__16004));
    InMux I__1679 (
            .O(N__16037),
            .I(N__16004));
    InMux I__1678 (
            .O(N__16036),
            .I(N__15999));
    InMux I__1677 (
            .O(N__16035),
            .I(N__15999));
    InMux I__1676 (
            .O(N__16034),
            .I(N__15992));
    InMux I__1675 (
            .O(N__16031),
            .I(N__15992));
    InMux I__1674 (
            .O(N__16030),
            .I(N__15992));
    InMux I__1673 (
            .O(N__16029),
            .I(N__15985));
    InMux I__1672 (
            .O(N__16028),
            .I(N__15985));
    InMux I__1671 (
            .O(N__16027),
            .I(N__15985));
    InMux I__1670 (
            .O(N__16026),
            .I(N__15977));
    InMux I__1669 (
            .O(N__16025),
            .I(N__15977));
    InMux I__1668 (
            .O(N__16024),
            .I(N__15970));
    InMux I__1667 (
            .O(N__16023),
            .I(N__15970));
    Span4Mux_v I__1666 (
            .O(N__16020),
            .I(N__15965));
    LocalMux I__1665 (
            .O(N__16009),
            .I(N__15965));
    LocalMux I__1664 (
            .O(N__16004),
            .I(N__15956));
    LocalMux I__1663 (
            .O(N__15999),
            .I(N__15956));
    LocalMux I__1662 (
            .O(N__15992),
            .I(N__15956));
    LocalMux I__1661 (
            .O(N__15985),
            .I(N__15956));
    InMux I__1660 (
            .O(N__15984),
            .I(N__15949));
    InMux I__1659 (
            .O(N__15983),
            .I(N__15949));
    InMux I__1658 (
            .O(N__15982),
            .I(N__15949));
    LocalMux I__1657 (
            .O(N__15977),
            .I(N__15946));
    InMux I__1656 (
            .O(N__15976),
            .I(N__15941));
    InMux I__1655 (
            .O(N__15975),
            .I(N__15941));
    LocalMux I__1654 (
            .O(N__15970),
            .I(N__15932));
    Span4Mux_s2_v I__1653 (
            .O(N__15965),
            .I(N__15932));
    Span4Mux_s2_v I__1652 (
            .O(N__15956),
            .I(N__15932));
    LocalMux I__1651 (
            .O(N__15949),
            .I(N__15932));
    Odrv12 I__1650 (
            .O(N__15946),
            .I(\b2v_inst16.N_26 ));
    LocalMux I__1649 (
            .O(N__15941),
            .I(\b2v_inst16.N_26 ));
    Odrv4 I__1648 (
            .O(N__15932),
            .I(\b2v_inst16.N_26 ));
    CascadeMux I__1647 (
            .O(N__15925),
            .I(\b2v_inst11.un1_func_state25_6_0_a3_0_0_cascade_ ));
    CascadeMux I__1646 (
            .O(N__15922),
            .I(\b2v_inst11.func_state_RNINPGR_2Z0Z_1_cascade_ ));
    InMux I__1645 (
            .O(N__15919),
            .I(N__15916));
    LocalMux I__1644 (
            .O(N__15916),
            .I(\b2v_inst11.g0_20_1 ));
    InMux I__1643 (
            .O(N__15913),
            .I(N__15910));
    LocalMux I__1642 (
            .O(N__15910),
            .I(\b2v_inst11.count_off_0_10 ));
    InMux I__1641 (
            .O(N__15907),
            .I(N__15904));
    LocalMux I__1640 (
            .O(N__15904),
            .I(\b2v_inst16.N_1440 ));
    CascadeMux I__1639 (
            .O(N__15901),
            .I(\b2v_inst16.curr_state_RNI3B692Z0Z_0_cascade_ ));
    CascadeMux I__1638 (
            .O(N__15898),
            .I(N__15891));
    InMux I__1637 (
            .O(N__15897),
            .I(N__15878));
    InMux I__1636 (
            .O(N__15896),
            .I(N__15873));
    InMux I__1635 (
            .O(N__15895),
            .I(N__15873));
    InMux I__1634 (
            .O(N__15894),
            .I(N__15870));
    InMux I__1633 (
            .O(N__15891),
            .I(N__15859));
    InMux I__1632 (
            .O(N__15890),
            .I(N__15859));
    InMux I__1631 (
            .O(N__15889),
            .I(N__15859));
    InMux I__1630 (
            .O(N__15888),
            .I(N__15859));
    InMux I__1629 (
            .O(N__15887),
            .I(N__15859));
    InMux I__1628 (
            .O(N__15886),
            .I(N__15856));
    InMux I__1627 (
            .O(N__15885),
            .I(N__15845));
    InMux I__1626 (
            .O(N__15884),
            .I(N__15845));
    InMux I__1625 (
            .O(N__15883),
            .I(N__15845));
    InMux I__1624 (
            .O(N__15882),
            .I(N__15845));
    InMux I__1623 (
            .O(N__15881),
            .I(N__15845));
    LocalMux I__1622 (
            .O(N__15878),
            .I(N__15838));
    LocalMux I__1621 (
            .O(N__15873),
            .I(N__15838));
    LocalMux I__1620 (
            .O(N__15870),
            .I(N__15838));
    LocalMux I__1619 (
            .O(N__15859),
            .I(\b2v_inst16.N_416 ));
    LocalMux I__1618 (
            .O(N__15856),
            .I(\b2v_inst16.N_416 ));
    LocalMux I__1617 (
            .O(N__15845),
            .I(\b2v_inst16.N_416 ));
    Odrv12 I__1616 (
            .O(N__15838),
            .I(\b2v_inst16.N_416 ));
    CascadeMux I__1615 (
            .O(N__15829),
            .I(\b2v_inst16.curr_state_7_0_1_cascade_ ));
    InMux I__1614 (
            .O(N__15826),
            .I(N__15823));
    LocalMux I__1613 (
            .O(N__15823),
            .I(\b2v_inst16.curr_state_2_1 ));
    CascadeMux I__1612 (
            .O(N__15820),
            .I(\b2v_inst16.curr_stateZ0Z_1_cascade_ ));
    InMux I__1611 (
            .O(N__15817),
            .I(N__15814));
    LocalMux I__1610 (
            .O(N__15814),
            .I(\b2v_inst16.curr_state_2_0 ));
    CascadeMux I__1609 (
            .O(N__15811),
            .I(N__15804));
    InMux I__1608 (
            .O(N__15810),
            .I(N__15795));
    InMux I__1607 (
            .O(N__15809),
            .I(N__15795));
    InMux I__1606 (
            .O(N__15808),
            .I(N__15795));
    InMux I__1605 (
            .O(N__15807),
            .I(N__15790));
    InMux I__1604 (
            .O(N__15804),
            .I(N__15790));
    InMux I__1603 (
            .O(N__15803),
            .I(N__15785));
    InMux I__1602 (
            .O(N__15802),
            .I(N__15785));
    LocalMux I__1601 (
            .O(N__15795),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    LocalMux I__1600 (
            .O(N__15790),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    LocalMux I__1599 (
            .O(N__15785),
            .I(\b2v_inst16.curr_stateZ0Z_1 ));
    CascadeMux I__1598 (
            .O(N__15778),
            .I(N__15774));
    InMux I__1597 (
            .O(N__15777),
            .I(N__15769));
    InMux I__1596 (
            .O(N__15774),
            .I(N__15762));
    InMux I__1595 (
            .O(N__15773),
            .I(N__15762));
    InMux I__1594 (
            .O(N__15772),
            .I(N__15762));
    LocalMux I__1593 (
            .O(N__15769),
            .I(\b2v_inst16.curr_state_RNI3B692Z0Z_0 ));
    LocalMux I__1592 (
            .O(N__15762),
            .I(\b2v_inst16.curr_state_RNI3B692Z0Z_0 ));
    InMux I__1591 (
            .O(N__15757),
            .I(N__15754));
    LocalMux I__1590 (
            .O(N__15754),
            .I(\b2v_inst16.N_268 ));
    InMux I__1589 (
            .O(N__15751),
            .I(N__15748));
    LocalMux I__1588 (
            .O(N__15748),
            .I(N__15745));
    Odrv4 I__1587 (
            .O(N__15745),
            .I(\b2v_inst16.count_4_i_a3_8_0 ));
    InMux I__1586 (
            .O(N__15742),
            .I(N__15739));
    LocalMux I__1585 (
            .O(N__15739),
            .I(\b2v_inst16.count_4_i_a3_10_0 ));
    CascadeMux I__1584 (
            .O(N__15736),
            .I(\b2v_inst16.count_4_i_a3_7_0_cascade_ ));
    InMux I__1583 (
            .O(N__15733),
            .I(N__15730));
    LocalMux I__1582 (
            .O(N__15730),
            .I(\b2v_inst16.count_4_i_a3_9_0 ));
    InMux I__1581 (
            .O(N__15727),
            .I(N__15721));
    InMux I__1580 (
            .O(N__15726),
            .I(N__15721));
    LocalMux I__1579 (
            .O(N__15721),
            .I(N__15718));
    Span4Mux_s0_v I__1578 (
            .O(N__15718),
            .I(N__15715));
    Odrv4 I__1577 (
            .O(N__15715),
            .I(\b2v_inst16.N_414 ));
    InMux I__1576 (
            .O(N__15712),
            .I(N__15702));
    InMux I__1575 (
            .O(N__15711),
            .I(N__15702));
    InMux I__1574 (
            .O(N__15710),
            .I(N__15702));
    CascadeMux I__1573 (
            .O(N__15709),
            .I(N__15699));
    LocalMux I__1572 (
            .O(N__15702),
            .I(N__15695));
    InMux I__1571 (
            .O(N__15699),
            .I(N__15692));
    InMux I__1570 (
            .O(N__15698),
            .I(N__15689));
    Span4Mux_v I__1569 (
            .O(N__15695),
            .I(N__15684));
    LocalMux I__1568 (
            .O(N__15692),
            .I(N__15684));
    LocalMux I__1567 (
            .O(N__15689),
            .I(\b2v_inst16.countZ0Z_0 ));
    Odrv4 I__1566 (
            .O(N__15684),
            .I(\b2v_inst16.countZ0Z_0 ));
    CascadeMux I__1565 (
            .O(N__15679),
            .I(\b2v_inst16.N_414_cascade_ ));
    InMux I__1564 (
            .O(N__15676),
            .I(N__15673));
    LocalMux I__1563 (
            .O(N__15673),
            .I(N__15670));
    Odrv12 I__1562 (
            .O(N__15670),
            .I(\b2v_inst16.count_4_0 ));
    CascadeMux I__1561 (
            .O(N__15667),
            .I(\b2v_inst11.count_offZ0Z_0_cascade_ ));
    InMux I__1560 (
            .O(N__15664),
            .I(N__15661));
    LocalMux I__1559 (
            .O(N__15661),
            .I(\b2v_inst11.count_off_RNIZ0Z_1 ));
    CascadeMux I__1558 (
            .O(N__15658),
            .I(\b2v_inst11.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__1557 (
            .O(N__15655),
            .I(N__15652));
    LocalMux I__1556 (
            .O(N__15652),
            .I(\b2v_inst11.count_off_0_1 ));
    CascadeMux I__1555 (
            .O(N__15649),
            .I(N__15646));
    InMux I__1554 (
            .O(N__15646),
            .I(N__15643));
    LocalMux I__1553 (
            .O(N__15643),
            .I(\b2v_inst11.count_off_0_0 ));
    CascadeMux I__1552 (
            .O(N__15640),
            .I(\b2v_inst16.count_rst_9_cascade_ ));
    CascadeMux I__1551 (
            .O(N__15637),
            .I(N__15634));
    InMux I__1550 (
            .O(N__15634),
            .I(N__15627));
    InMux I__1549 (
            .O(N__15633),
            .I(N__15627));
    InMux I__1548 (
            .O(N__15632),
            .I(N__15624));
    LocalMux I__1547 (
            .O(N__15627),
            .I(\b2v_inst16.countZ0Z_4 ));
    LocalMux I__1546 (
            .O(N__15624),
            .I(\b2v_inst16.countZ0Z_4 ));
    InMux I__1545 (
            .O(N__15619),
            .I(N__15613));
    InMux I__1544 (
            .O(N__15618),
            .I(N__15613));
    LocalMux I__1543 (
            .O(N__15613),
            .I(\b2v_inst16.un4_count_1_cry_3_THRU_CO ));
    CascadeMux I__1542 (
            .O(N__15610),
            .I(\b2v_inst16.countZ0Z_4_cascade_ ));
    InMux I__1541 (
            .O(N__15607),
            .I(N__15604));
    LocalMux I__1540 (
            .O(N__15604),
            .I(\b2v_inst16.count_4_4 ));
    InMux I__1539 (
            .O(N__15601),
            .I(N__15595));
    InMux I__1538 (
            .O(N__15600),
            .I(N__15595));
    LocalMux I__1537 (
            .O(N__15595),
            .I(\b2v_inst16.count_rst_2 ));
    InMux I__1536 (
            .O(N__15592),
            .I(N__15589));
    LocalMux I__1535 (
            .O(N__15589),
            .I(\b2v_inst16.count_4_13 ));
    CascadeMux I__1534 (
            .O(N__15586),
            .I(\b2v_inst16.un4_count_1_axb_1_cascade_ ));
    InMux I__1533 (
            .O(N__15583),
            .I(N__15579));
    InMux I__1532 (
            .O(N__15582),
            .I(N__15576));
    LocalMux I__1531 (
            .O(N__15579),
            .I(\b2v_inst16.un4_count_1_axb_1 ));
    LocalMux I__1530 (
            .O(N__15576),
            .I(\b2v_inst16.un4_count_1_axb_1 ));
    InMux I__1529 (
            .O(N__15571),
            .I(N__15568));
    LocalMux I__1528 (
            .O(N__15568),
            .I(N__15565));
    Span4Mux_s2_h I__1527 (
            .O(N__15565),
            .I(N__15561));
    InMux I__1526 (
            .O(N__15564),
            .I(N__15558));
    Odrv4 I__1525 (
            .O(N__15561),
            .I(\b2v_inst16.countZ0Z_6 ));
    LocalMux I__1524 (
            .O(N__15558),
            .I(\b2v_inst16.countZ0Z_6 ));
    InMux I__1523 (
            .O(N__15553),
            .I(N__15549));
    InMux I__1522 (
            .O(N__15552),
            .I(N__15546));
    LocalMux I__1521 (
            .O(N__15549),
            .I(\b2v_inst16.countZ0Z_12 ));
    LocalMux I__1520 (
            .O(N__15546),
            .I(\b2v_inst16.countZ0Z_12 ));
    CascadeMux I__1519 (
            .O(N__15541),
            .I(N__15537));
    CascadeMux I__1518 (
            .O(N__15540),
            .I(N__15534));
    InMux I__1517 (
            .O(N__15537),
            .I(N__15531));
    InMux I__1516 (
            .O(N__15534),
            .I(N__15528));
    LocalMux I__1515 (
            .O(N__15531),
            .I(N__15523));
    LocalMux I__1514 (
            .O(N__15528),
            .I(N__15523));
    Odrv4 I__1513 (
            .O(N__15523),
            .I(\b2v_inst16.countZ0Z_10 ));
    InMux I__1512 (
            .O(N__15520),
            .I(N__15516));
    InMux I__1511 (
            .O(N__15519),
            .I(N__15513));
    LocalMux I__1510 (
            .O(N__15516),
            .I(N__15510));
    LocalMux I__1509 (
            .O(N__15513),
            .I(N__15507));
    Odrv4 I__1508 (
            .O(N__15510),
            .I(\b2v_inst16.countZ0Z_2 ));
    Odrv12 I__1507 (
            .O(N__15507),
            .I(\b2v_inst16.countZ0Z_2 ));
    InMux I__1506 (
            .O(N__15502),
            .I(N__15498));
    InMux I__1505 (
            .O(N__15501),
            .I(N__15495));
    LocalMux I__1504 (
            .O(N__15498),
            .I(\b2v_inst16.count_4_1 ));
    LocalMux I__1503 (
            .O(N__15495),
            .I(\b2v_inst16.count_4_1 ));
    InMux I__1502 (
            .O(N__15490),
            .I(N__15484));
    InMux I__1501 (
            .O(N__15489),
            .I(N__15484));
    LocalMux I__1500 (
            .O(N__15484),
            .I(\b2v_inst16.count_rst_6 ));
    InMux I__1499 (
            .O(N__15481),
            .I(N__15478));
    LocalMux I__1498 (
            .O(N__15478),
            .I(N__15474));
    InMux I__1497 (
            .O(N__15477),
            .I(N__15471));
    Span12Mux_s1_h I__1496 (
            .O(N__15474),
            .I(N__15466));
    LocalMux I__1495 (
            .O(N__15471),
            .I(N__15466));
    Odrv12 I__1494 (
            .O(N__15466),
            .I(\b2v_inst16.countZ0Z_15 ));
    CascadeMux I__1493 (
            .O(N__15463),
            .I(\b2v_inst16.countZ0Z_1_cascade_ ));
    InMux I__1492 (
            .O(N__15460),
            .I(N__15457));
    LocalMux I__1491 (
            .O(N__15457),
            .I(N__15453));
    InMux I__1490 (
            .O(N__15456),
            .I(N__15449));
    Span4Mux_v I__1489 (
            .O(N__15453),
            .I(N__15446));
    InMux I__1488 (
            .O(N__15452),
            .I(N__15443));
    LocalMux I__1487 (
            .O(N__15449),
            .I(N__15440));
    Odrv4 I__1486 (
            .O(N__15446),
            .I(\b2v_inst16.countZ0Z_11 ));
    LocalMux I__1485 (
            .O(N__15443),
            .I(\b2v_inst16.countZ0Z_11 ));
    Odrv12 I__1484 (
            .O(N__15440),
            .I(\b2v_inst16.countZ0Z_11 ));
    InMux I__1483 (
            .O(N__15433),
            .I(N__15427));
    InMux I__1482 (
            .O(N__15432),
            .I(N__15427));
    LocalMux I__1481 (
            .O(N__15427),
            .I(N__15424));
    Span4Mux_s1_v I__1480 (
            .O(N__15424),
            .I(N__15421));
    Odrv4 I__1479 (
            .O(N__15421),
            .I(\b2v_inst16.count_rst_4 ));
    InMux I__1478 (
            .O(N__15418),
            .I(N__15415));
    LocalMux I__1477 (
            .O(N__15415),
            .I(\b2v_inst16.count_4_15 ));
    InMux I__1476 (
            .O(N__15412),
            .I(N__15409));
    LocalMux I__1475 (
            .O(N__15409),
            .I(\b2v_inst16.count_4_14 ));
    InMux I__1474 (
            .O(N__15406),
            .I(N__15400));
    InMux I__1473 (
            .O(N__15405),
            .I(N__15400));
    LocalMux I__1472 (
            .O(N__15400),
            .I(\b2v_inst16.count_rst_3 ));
    InMux I__1471 (
            .O(N__15397),
            .I(N__15394));
    LocalMux I__1470 (
            .O(N__15394),
            .I(\b2v_inst16.countZ0Z_14 ));
    CascadeMux I__1469 (
            .O(N__15391),
            .I(N__15386));
    InMux I__1468 (
            .O(N__15390),
            .I(N__15383));
    InMux I__1467 (
            .O(N__15389),
            .I(N__15380));
    InMux I__1466 (
            .O(N__15386),
            .I(N__15377));
    LocalMux I__1465 (
            .O(N__15383),
            .I(N__15374));
    LocalMux I__1464 (
            .O(N__15380),
            .I(N__15371));
    LocalMux I__1463 (
            .O(N__15377),
            .I(\b2v_inst16.countZ0Z_3 ));
    Odrv4 I__1462 (
            .O(N__15374),
            .I(\b2v_inst16.countZ0Z_3 ));
    Odrv4 I__1461 (
            .O(N__15371),
            .I(\b2v_inst16.countZ0Z_3 ));
    CascadeMux I__1460 (
            .O(N__15364),
            .I(\b2v_inst16.countZ0Z_14_cascade_ ));
    InMux I__1459 (
            .O(N__15361),
            .I(N__15357));
    InMux I__1458 (
            .O(N__15360),
            .I(N__15354));
    LocalMux I__1457 (
            .O(N__15357),
            .I(\b2v_inst16.countZ0Z_13 ));
    LocalMux I__1456 (
            .O(N__15354),
            .I(\b2v_inst16.countZ0Z_13 ));
    InMux I__1455 (
            .O(N__15349),
            .I(N__15345));
    InMux I__1454 (
            .O(N__15348),
            .I(N__15341));
    LocalMux I__1453 (
            .O(N__15345),
            .I(N__15338));
    InMux I__1452 (
            .O(N__15344),
            .I(N__15335));
    LocalMux I__1451 (
            .O(N__15341),
            .I(N__15332));
    Odrv4 I__1450 (
            .O(N__15338),
            .I(\b2v_inst16.countZ0Z_8 ));
    LocalMux I__1449 (
            .O(N__15335),
            .I(\b2v_inst16.countZ0Z_8 ));
    Odrv4 I__1448 (
            .O(N__15332),
            .I(\b2v_inst16.countZ0Z_8 ));
    CascadeMux I__1447 (
            .O(N__15325),
            .I(\b2v_inst16.N_416_cascade_ ));
    InMux I__1446 (
            .O(N__15322),
            .I(N__15318));
    InMux I__1445 (
            .O(N__15321),
            .I(N__15315));
    LocalMux I__1444 (
            .O(N__15318),
            .I(N__15310));
    LocalMux I__1443 (
            .O(N__15315),
            .I(N__15310));
    Odrv4 I__1442 (
            .O(N__15310),
            .I(\b2v_inst16.un4_count_1_cry_7_THRU_CO ));
    InMux I__1441 (
            .O(N__15307),
            .I(N__15304));
    LocalMux I__1440 (
            .O(N__15304),
            .I(\b2v_inst16.count_rst_13 ));
    InMux I__1439 (
            .O(N__15301),
            .I(N__15298));
    LocalMux I__1438 (
            .O(N__15298),
            .I(\b2v_inst16.count_rst_5 ));
    CascadeMux I__1437 (
            .O(N__15295),
            .I(N__15291));
    CascadeMux I__1436 (
            .O(N__15294),
            .I(N__15288));
    InMux I__1435 (
            .O(N__15291),
            .I(N__15285));
    InMux I__1434 (
            .O(N__15288),
            .I(N__15282));
    LocalMux I__1433 (
            .O(N__15285),
            .I(N__15279));
    LocalMux I__1432 (
            .O(N__15282),
            .I(\b2v_inst16.un4_count_1_cry_4_THRU_CO ));
    Odrv4 I__1431 (
            .O(N__15279),
            .I(\b2v_inst16.un4_count_1_cry_4_THRU_CO ));
    CascadeMux I__1430 (
            .O(N__15274),
            .I(\b2v_inst16.count_rst_10_cascade_ ));
    InMux I__1429 (
            .O(N__15271),
            .I(N__15268));
    LocalMux I__1428 (
            .O(N__15268),
            .I(\b2v_inst16.count_4_5 ));
    InMux I__1427 (
            .O(N__15265),
            .I(N__15259));
    InMux I__1426 (
            .O(N__15264),
            .I(N__15256));
    InMux I__1425 (
            .O(N__15263),
            .I(N__15253));
    InMux I__1424 (
            .O(N__15262),
            .I(N__15250));
    LocalMux I__1423 (
            .O(N__15259),
            .I(N__15247));
    LocalMux I__1422 (
            .O(N__15256),
            .I(\b2v_inst16.countZ0Z_5 ));
    LocalMux I__1421 (
            .O(N__15253),
            .I(\b2v_inst16.countZ0Z_5 ));
    LocalMux I__1420 (
            .O(N__15250),
            .I(\b2v_inst16.countZ0Z_5 ));
    Odrv4 I__1419 (
            .O(N__15247),
            .I(\b2v_inst16.countZ0Z_5 ));
    InMux I__1418 (
            .O(N__15238),
            .I(N__15232));
    InMux I__1417 (
            .O(N__15237),
            .I(N__15232));
    LocalMux I__1416 (
            .O(N__15232),
            .I(N__15229));
    Odrv4 I__1415 (
            .O(N__15229),
            .I(\b2v_inst16.count_rst ));
    InMux I__1414 (
            .O(N__15226),
            .I(N__15223));
    LocalMux I__1413 (
            .O(N__15223),
            .I(\b2v_inst16.count_4_10 ));
    InMux I__1412 (
            .O(N__15220),
            .I(N__15214));
    InMux I__1411 (
            .O(N__15219),
            .I(N__15214));
    LocalMux I__1410 (
            .O(N__15214),
            .I(\b2v_inst16.count_rst_11 ));
    InMux I__1409 (
            .O(N__15211),
            .I(N__15208));
    LocalMux I__1408 (
            .O(N__15208),
            .I(\b2v_inst16.count_4_6 ));
    InMux I__1407 (
            .O(N__15205),
            .I(bfn_1_16_0_));
    InMux I__1406 (
            .O(N__15202),
            .I(\b2v_inst20.counter_1_cry_25 ));
    InMux I__1405 (
            .O(N__15199),
            .I(\b2v_inst20.counter_1_cry_26 ));
    InMux I__1404 (
            .O(N__15196),
            .I(\b2v_inst20.counter_1_cry_27 ));
    InMux I__1403 (
            .O(N__15193),
            .I(\b2v_inst20.counter_1_cry_28 ));
    InMux I__1402 (
            .O(N__15190),
            .I(\b2v_inst20.counter_1_cry_29 ));
    InMux I__1401 (
            .O(N__15187),
            .I(\b2v_inst20.counter_1_cry_30 ));
    CascadeMux I__1400 (
            .O(N__15184),
            .I(\b2v_inst16.countZ0Z_0_cascade_ ));
    InMux I__1399 (
            .O(N__15181),
            .I(\b2v_inst20.counter_1_cry_15 ));
    InMux I__1398 (
            .O(N__15178),
            .I(bfn_1_15_0_));
    InMux I__1397 (
            .O(N__15175),
            .I(\b2v_inst20.counter_1_cry_17 ));
    InMux I__1396 (
            .O(N__15172),
            .I(\b2v_inst20.counter_1_cry_18 ));
    InMux I__1395 (
            .O(N__15169),
            .I(\b2v_inst20.counter_1_cry_19 ));
    InMux I__1394 (
            .O(N__15166),
            .I(\b2v_inst20.counter_1_cry_20 ));
    InMux I__1393 (
            .O(N__15163),
            .I(\b2v_inst20.counter_1_cry_21 ));
    InMux I__1392 (
            .O(N__15160),
            .I(\b2v_inst20.counter_1_cry_22 ));
    InMux I__1391 (
            .O(N__15157),
            .I(\b2v_inst20.counter_1_cry_23 ));
    InMux I__1390 (
            .O(N__15154),
            .I(\b2v_inst20.counter_1_cry_6 ));
    InMux I__1389 (
            .O(N__15151),
            .I(\b2v_inst20.counter_1_cry_7 ));
    InMux I__1388 (
            .O(N__15148),
            .I(bfn_1_14_0_));
    InMux I__1387 (
            .O(N__15145),
            .I(\b2v_inst20.counter_1_cry_9 ));
    InMux I__1386 (
            .O(N__15142),
            .I(\b2v_inst20.counter_1_cry_10 ));
    InMux I__1385 (
            .O(N__15139),
            .I(\b2v_inst20.counter_1_cry_11 ));
    InMux I__1384 (
            .O(N__15136),
            .I(\b2v_inst20.counter_1_cry_12 ));
    InMux I__1383 (
            .O(N__15133),
            .I(\b2v_inst20.counter_1_cry_13 ));
    InMux I__1382 (
            .O(N__15130),
            .I(\b2v_inst20.counter_1_cry_14 ));
    InMux I__1381 (
            .O(N__15127),
            .I(N__15123));
    InMux I__1380 (
            .O(N__15126),
            .I(N__15120));
    LocalMux I__1379 (
            .O(N__15123),
            .I(N__15115));
    LocalMux I__1378 (
            .O(N__15120),
            .I(N__15115));
    Odrv4 I__1377 (
            .O(N__15115),
            .I(\b2v_inst11.un2_count_clk_17_0_o2_4 ));
    InMux I__1376 (
            .O(N__15112),
            .I(N__15109));
    LocalMux I__1375 (
            .O(N__15109),
            .I(\b2v_inst11.count_clk_0_11 ));
    InMux I__1374 (
            .O(N__15106),
            .I(N__15103));
    LocalMux I__1373 (
            .O(N__15103),
            .I(N__15100));
    Odrv4 I__1372 (
            .O(N__15100),
            .I(\b2v_inst11.count_clk_0_4 ));
    InMux I__1371 (
            .O(N__15097),
            .I(\b2v_inst20.counter_1_cry_1 ));
    InMux I__1370 (
            .O(N__15094),
            .I(\b2v_inst20.counter_1_cry_2 ));
    InMux I__1369 (
            .O(N__15091),
            .I(\b2v_inst20.counter_1_cry_3 ));
    InMux I__1368 (
            .O(N__15088),
            .I(\b2v_inst20.counter_1_cry_4 ));
    InMux I__1367 (
            .O(N__15085),
            .I(\b2v_inst20.counter_1_cry_5 ));
    CascadeMux I__1366 (
            .O(N__15082),
            .I(\b2v_inst11.count_clk_en_cascade_ ));
    InMux I__1365 (
            .O(N__15079),
            .I(N__15076));
    LocalMux I__1364 (
            .O(N__15076),
            .I(\b2v_inst11.count_clk_0_13 ));
    InMux I__1363 (
            .O(N__15073),
            .I(N__15070));
    LocalMux I__1362 (
            .O(N__15070),
            .I(\b2v_inst11.count_clk_0_15 ));
    CascadeMux I__1361 (
            .O(N__15067),
            .I(N__15064));
    InMux I__1360 (
            .O(N__15064),
            .I(N__15061));
    LocalMux I__1359 (
            .O(N__15061),
            .I(\b2v_inst11.count_clk_0_12 ));
    InMux I__1358 (
            .O(N__15058),
            .I(N__15055));
    LocalMux I__1357 (
            .O(N__15055),
            .I(\b2v_inst11.count_clk_0_10 ));
    CascadeMux I__1356 (
            .O(N__15052),
            .I(\b2v_inst11.count_clkZ0Z_10_cascade_ ));
    InMux I__1355 (
            .O(N__15049),
            .I(N__15046));
    LocalMux I__1354 (
            .O(N__15046),
            .I(N__15043));
    Odrv4 I__1353 (
            .O(N__15043),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2 ));
    InMux I__1352 (
            .O(N__15040),
            .I(N__15037));
    LocalMux I__1351 (
            .O(N__15037),
            .I(\b2v_inst11.count_clk_RNIVS8U1Z0Z_14 ));
    CascadeMux I__1350 (
            .O(N__15034),
            .I(N__15031));
    InMux I__1349 (
            .O(N__15031),
            .I(N__15028));
    LocalMux I__1348 (
            .O(N__15028),
            .I(\b2v_inst11.N_428 ));
    InMux I__1347 (
            .O(N__15025),
            .I(N__15022));
    LocalMux I__1346 (
            .O(N__15022),
            .I(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0 ));
    InMux I__1345 (
            .O(N__15019),
            .I(N__15016));
    LocalMux I__1344 (
            .O(N__15016),
            .I(\b2v_inst11.N_175 ));
    CascadeMux I__1343 (
            .O(N__15013),
            .I(\b2v_inst11.N_175_cascade_ ));
    InMux I__1342 (
            .O(N__15010),
            .I(N__15007));
    LocalMux I__1341 (
            .O(N__15007),
            .I(\b2v_inst11.N_190 ));
    CascadeMux I__1340 (
            .O(N__15004),
            .I(\b2v_inst11.N_190_cascade_ ));
    InMux I__1339 (
            .O(N__15001),
            .I(N__14998));
    LocalMux I__1338 (
            .O(N__14998),
            .I(\b2v_inst11.un2_count_clk_17_0_o3_0_4 ));
    CascadeMux I__1337 (
            .O(N__14995),
            .I(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ));
    CascadeMux I__1336 (
            .O(N__14992),
            .I(\b2v_inst11.N_379_cascade_ ));
    CascadeMux I__1335 (
            .O(N__14989),
            .I(N__14986));
    InMux I__1334 (
            .O(N__14986),
            .I(N__14983));
    LocalMux I__1333 (
            .O(N__14983),
            .I(SLP_S3n_ibuf_RNIF6NLZ0));
    InMux I__1332 (
            .O(N__14980),
            .I(N__14974));
    InMux I__1331 (
            .O(N__14979),
            .I(N__14974));
    LocalMux I__1330 (
            .O(N__14974),
            .I(N__14971));
    Odrv4 I__1329 (
            .O(N__14971),
            .I(\b2v_inst11.N_379 ));
    CascadeMux I__1328 (
            .O(N__14968),
            .I(N__14965));
    InMux I__1327 (
            .O(N__14965),
            .I(N__14962));
    LocalMux I__1326 (
            .O(N__14962),
            .I(\b2v_inst11.count_clk_RNI_0Z0Z_13 ));
    CascadeMux I__1325 (
            .O(N__14959),
            .I(\b2v_inst11.g3_cascade_ ));
    CascadeMux I__1324 (
            .O(N__14956),
            .I(\b2v_inst11.g1_0_1_cascade_ ));
    CascadeMux I__1323 (
            .O(N__14953),
            .I(\b2v_inst11.N_7_3_0_cascade_ ));
    CascadeMux I__1322 (
            .O(N__14950),
            .I(\b2v_inst11.g2_1_0_0_cascade_ ));
    InMux I__1321 (
            .O(N__14947),
            .I(N__14944));
    LocalMux I__1320 (
            .O(N__14944),
            .I(\b2v_inst11.g2_2_0 ));
    InMux I__1319 (
            .O(N__14941),
            .I(N__14938));
    LocalMux I__1318 (
            .O(N__14938),
            .I(N__14935));
    Span4Mux_v I__1317 (
            .O(N__14935),
            .I(N__14932));
    Odrv4 I__1316 (
            .O(N__14932),
            .I(\b2v_inst11.g2_1_0 ));
    InMux I__1315 (
            .O(N__14929),
            .I(N__14926));
    LocalMux I__1314 (
            .O(N__14926),
            .I(\b2v_inst11.g0_12_0 ));
    InMux I__1313 (
            .O(N__14923),
            .I(N__14920));
    LocalMux I__1312 (
            .O(N__14920),
            .I(\b2v_inst16.delayed_vddq_pwrgd_en ));
    CascadeMux I__1311 (
            .O(N__14917),
            .I(N__14913));
    InMux I__1310 (
            .O(N__14916),
            .I(N__14908));
    InMux I__1309 (
            .O(N__14913),
            .I(N__14908));
    LocalMux I__1308 (
            .O(N__14908),
            .I(\b2v_inst16.delayed_vddq_pwrgdZ0 ));
    CascadeMux I__1307 (
            .O(N__14905),
            .I(\b2v_inst16.delayed_vddq_pwrgd_en_cascade_ ));
    IoInMux I__1306 (
            .O(N__14902),
            .I(N__14899));
    LocalMux I__1305 (
            .O(N__14899),
            .I(N__14896));
    IoSpan4Mux I__1304 (
            .O(N__14896),
            .I(N__14893));
    IoSpan4Mux I__1303 (
            .O(N__14893),
            .I(N__14890));
    Odrv4 I__1302 (
            .O(N__14890),
            .I(b2v_inst16_un2_vpp_en_0_i));
    IoInMux I__1301 (
            .O(N__14887),
            .I(N__14884));
    LocalMux I__1300 (
            .O(N__14884),
            .I(N__14881));
    Span4Mux_s0_h I__1299 (
            .O(N__14881),
            .I(N__14878));
    Odrv4 I__1298 (
            .O(N__14878),
            .I(\b2v_inst200.count_enZ0 ));
    InMux I__1297 (
            .O(N__14875),
            .I(N__14871));
    InMux I__1296 (
            .O(N__14874),
            .I(N__14868));
    LocalMux I__1295 (
            .O(N__14871),
            .I(N__14865));
    LocalMux I__1294 (
            .O(N__14868),
            .I(N__14862));
    Odrv12 I__1293 (
            .O(N__14865),
            .I(\b2v_inst16.count_rst_7 ));
    Odrv4 I__1292 (
            .O(N__14862),
            .I(\b2v_inst16.count_rst_7 ));
    CascadeMux I__1291 (
            .O(N__14857),
            .I(\b2v_inst16.count_en_cascade_ ));
    InMux I__1290 (
            .O(N__14854),
            .I(N__14851));
    LocalMux I__1289 (
            .O(N__14851),
            .I(\b2v_inst16.count_4_2 ));
    CascadeMux I__1288 (
            .O(N__14848),
            .I(N__14845));
    InMux I__1287 (
            .O(N__14845),
            .I(N__14838));
    InMux I__1286 (
            .O(N__14844),
            .I(N__14838));
    InMux I__1285 (
            .O(N__14843),
            .I(N__14835));
    LocalMux I__1284 (
            .O(N__14838),
            .I(\b2v_inst16.countZ0Z_7 ));
    LocalMux I__1283 (
            .O(N__14835),
            .I(\b2v_inst16.countZ0Z_7 ));
    InMux I__1282 (
            .O(N__14830),
            .I(N__14824));
    InMux I__1281 (
            .O(N__14829),
            .I(N__14824));
    LocalMux I__1280 (
            .O(N__14824),
            .I(\b2v_inst16.un4_count_1_cry_6_THRU_CO ));
    InMux I__1279 (
            .O(N__14821),
            .I(\b2v_inst16.un4_count_1_cry_6 ));
    InMux I__1278 (
            .O(N__14818),
            .I(\b2v_inst16.un4_count_1_cry_7 ));
    InMux I__1277 (
            .O(N__14815),
            .I(N__14810));
    InMux I__1276 (
            .O(N__14814),
            .I(N__14805));
    InMux I__1275 (
            .O(N__14813),
            .I(N__14805));
    LocalMux I__1274 (
            .O(N__14810),
            .I(N__14802));
    LocalMux I__1273 (
            .O(N__14805),
            .I(\b2v_inst16.countZ0Z_9 ));
    Odrv4 I__1272 (
            .O(N__14802),
            .I(\b2v_inst16.countZ0Z_9 ));
    InMux I__1271 (
            .O(N__14797),
            .I(N__14791));
    InMux I__1270 (
            .O(N__14796),
            .I(N__14791));
    LocalMux I__1269 (
            .O(N__14791),
            .I(N__14788));
    Odrv4 I__1268 (
            .O(N__14788),
            .I(\b2v_inst16.un4_count_1_cry_8_THRU_CO ));
    InMux I__1267 (
            .O(N__14785),
            .I(bfn_1_4_0_));
    InMux I__1266 (
            .O(N__14782),
            .I(\b2v_inst16.un4_count_1_cry_9 ));
    InMux I__1265 (
            .O(N__14779),
            .I(N__14773));
    InMux I__1264 (
            .O(N__14778),
            .I(N__14773));
    LocalMux I__1263 (
            .O(N__14773),
            .I(N__14770));
    Odrv4 I__1262 (
            .O(N__14770),
            .I(\b2v_inst16.un4_count_1_cry_10_THRU_CO ));
    InMux I__1261 (
            .O(N__14767),
            .I(\b2v_inst16.un4_count_1_cry_10 ));
    InMux I__1260 (
            .O(N__14764),
            .I(\b2v_inst16.un4_count_1_cry_11 ));
    InMux I__1259 (
            .O(N__14761),
            .I(\b2v_inst16.un4_count_1_cry_12 ));
    InMux I__1258 (
            .O(N__14758),
            .I(\b2v_inst16.un4_count_1_cry_13 ));
    InMux I__1257 (
            .O(N__14755),
            .I(\b2v_inst16.un4_count_1_cry_14 ));
    CascadeMux I__1256 (
            .O(N__14752),
            .I(\b2v_inst16.count_rst_12_cascade_ ));
    CascadeMux I__1255 (
            .O(N__14749),
            .I(\b2v_inst16.countZ0Z_7_cascade_ ));
    InMux I__1254 (
            .O(N__14746),
            .I(N__14743));
    LocalMux I__1253 (
            .O(N__14743),
            .I(\b2v_inst16.count_4_7 ));
    InMux I__1252 (
            .O(N__14740),
            .I(\b2v_inst16.un4_count_1_cry_1 ));
    InMux I__1251 (
            .O(N__14737),
            .I(N__14731));
    InMux I__1250 (
            .O(N__14736),
            .I(N__14731));
    LocalMux I__1249 (
            .O(N__14731),
            .I(N__14728));
    Odrv4 I__1248 (
            .O(N__14728),
            .I(\b2v_inst16.un4_count_1_cry_2_THRU_CO ));
    InMux I__1247 (
            .O(N__14725),
            .I(\b2v_inst16.un4_count_1_cry_2 ));
    InMux I__1246 (
            .O(N__14722),
            .I(\b2v_inst16.un4_count_1_cry_3 ));
    InMux I__1245 (
            .O(N__14719),
            .I(\b2v_inst16.un4_count_1_cry_4 ));
    InMux I__1244 (
            .O(N__14716),
            .I(\b2v_inst16.un4_count_1_cry_5 ));
    CascadeMux I__1243 (
            .O(N__14713),
            .I(\b2v_inst16.countZ0Z_8_cascade_ ));
    InMux I__1242 (
            .O(N__14710),
            .I(N__14707));
    LocalMux I__1241 (
            .O(N__14707),
            .I(\b2v_inst16.count_4_8 ));
    CascadeMux I__1240 (
            .O(N__14704),
            .I(\b2v_inst16.count_rst_8_cascade_ ));
    CascadeMux I__1239 (
            .O(N__14701),
            .I(\b2v_inst16.countZ0Z_3_cascade_ ));
    InMux I__1238 (
            .O(N__14698),
            .I(N__14695));
    LocalMux I__1237 (
            .O(N__14695),
            .I(\b2v_inst16.count_4_3 ));
    CascadeMux I__1236 (
            .O(N__14692),
            .I(\b2v_inst16.countZ0Z_9_cascade_ ));
    InMux I__1235 (
            .O(N__14689),
            .I(N__14686));
    LocalMux I__1234 (
            .O(N__14686),
            .I(\b2v_inst16.count_rst_14 ));
    InMux I__1233 (
            .O(N__14683),
            .I(N__14680));
    LocalMux I__1232 (
            .O(N__14680),
            .I(\b2v_inst16.count_4_9 ));
    CascadeMux I__1231 (
            .O(N__14677),
            .I(\b2v_inst16.count_rst_0_cascade_ ));
    CascadeMux I__1230 (
            .O(N__14674),
            .I(\b2v_inst16.countZ0Z_11_cascade_ ));
    InMux I__1229 (
            .O(N__14671),
            .I(N__14668));
    LocalMux I__1228 (
            .O(N__14668),
            .I(\b2v_inst16.count_4_11 ));
    defparam IN_MUX_bfv_12_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_1_0_));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(\b2v_inst6.un2_count_1_cry_8 ),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\b2v_inst5.un2_count_1_cry_8 ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_9_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_2_0_ (
            .carryinitin(\b2v_inst36.un2_count_1_cry_8 ),
            .carryinitout(bfn_9_2_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(b2v_inst20_un4_counter_7),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_8 ),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_16 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\b2v_inst20.counter_1_cry_24 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(\b2v_inst16.un4_count_1_cry_8 ),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(\b2v_inst11.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\b2v_inst11.un1_count_cry_8 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\b2v_inst11.un1_count_clk_2_cry_8 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_5_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_1_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_7 ),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\b2v_inst200.un2_count_1_cry_15 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\b2v_inst11.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    ICE_GB \b2v_inst200.count_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__14887),
            .GLOBALBUFFEROUTPUT(\b2v_inst200.count_en_g ));
    ICE_GB N_606_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__27603),
            .GLOBALBUFFEROUTPUT(N_606_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_1_0 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_c_RNIQPK3_LC_1_1_0  (
            .in0(N__15882),
            .in1(N__14778),
            .in2(N__16053),
            .in3(N__15452),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIDGU31_11_LC_1_1_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIDGU31_11_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIDGU31_11_LC_1_1_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst16.count_RNIDGU31_11_LC_1_1_1  (
            .in0(N__20937),
            .in1(_gnd_net_),
            .in2(N__14677),
            .in3(N__14671),
            .lcout(\b2v_inst16.countZ0Z_11 ),
            .ltout(\b2v_inst16.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_11_LC_1_1_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_11_LC_1_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_11_LC_1_1_2 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_11_LC_1_1_2  (
            .in0(N__15883),
            .in1(N__16037),
            .in2(N__14674),
            .in3(N__14779),
            .lcout(\b2v_inst16.count_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36609),
            .ce(N__20949),
            .sr(N__20799));
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNIPM3K1_8_LC_1_1_3  (
            .in0(N__20936),
            .in1(N__14710),
            .in2(_gnd_net_),
            .in3(N__15307),
            .lcout(\b2v_inst16.countZ0Z_8 ),
            .ltout(\b2v_inst16.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_8_LC_1_1_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_8_LC_1_1_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_8_LC_1_1_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst16.count_8_LC_1_1_4  (
            .in0(N__15884),
            .in1(N__16038),
            .in2(N__14713),
            .in3(N__15322),
            .lcout(\b2v_inst16.count_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36609),
            .ce(N__20949),
            .sr(N__20799));
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_1_5 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_1_5 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_c_RNIBINE_LC_1_1_5  (
            .in0(N__14736),
            .in1(N__16030),
            .in2(N__15391),
            .in3(N__15881),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIF7UJ1_3_LC_1_1_6  (
            .in0(_gnd_net_),
            .in1(N__14698),
            .in2(N__14704),
            .in3(N__20935),
            .lcout(\b2v_inst16.countZ0Z_3 ),
            .ltout(\b2v_inst16.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_3_LC_1_1_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_3_LC_1_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_3_LC_1_1_7 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.count_3_LC_1_1_7  (
            .in0(N__14737),
            .in1(N__16034),
            .in2(N__14701),
            .in3(N__15885),
            .lcout(\b2v_inst16.count_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36609),
            .ce(N__20949),
            .sr(N__20799));
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_1_2_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIRP4K1_9_LC_1_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNIRP4K1_9_LC_1_2_0  (
            .in0(N__20941),
            .in1(N__14683),
            .in2(_gnd_net_),
            .in3(N__14689),
            .lcout(\b2v_inst16.countZ0Z_9 ),
            .ltout(\b2v_inst16.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_5_LC_1_2_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_5_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_5_LC_1_2_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst16.count_RNI_5_LC_1_2_1  (
            .in0(N__15262),
            .in1(N__14844),
            .in2(N__14692),
            .in3(N__15344),
            .lcout(\b2v_inst16.count_4_i_a3_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_2_2 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_2_2 .LUT_INIT=16'b0001000000100000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_c_RNIHUTE_LC_1_2_2  (
            .in0(N__14814),
            .in1(N__15888),
            .in2(N__16054),
            .in3(N__14796),
            .lcout(\b2v_inst16.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_9_LC_1_2_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_9_LC_1_2_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_9_LC_1_2_3 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst16.count_9_LC_1_2_3  (
            .in0(N__14797),
            .in1(N__16044),
            .in2(N__15898),
            .in3(N__14813),
            .lcout(\b2v_inst16.count_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36601),
            .ce(N__20928),
            .sr(N__20785));
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_4 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_4 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_c_RNIFQRE_LC_1_2_4  (
            .in0(N__16039),
            .in1(N__15887),
            .in2(N__14848),
            .in3(N__14829),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_2_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNINJ2K1_7_LC_1_2_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNINJ2K1_7_LC_1_2_5  (
            .in0(_gnd_net_),
            .in1(N__14746),
            .in2(N__14752),
            .in3(N__20940),
            .lcout(\b2v_inst16.countZ0Z_7 ),
            .ltout(\b2v_inst16.countZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_7_LC_1_2_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_7_LC_1_2_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_7_LC_1_2_6 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \b2v_inst16.count_7_LC_1_2_6  (
            .in0(N__16043),
            .in1(N__15890),
            .in2(N__14749),
            .in3(N__14830),
            .lcout(\b2v_inst16.count_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36601),
            .ce(N__20928),
            .sr(N__20785));
    defparam \b2v_inst16.count_5_LC_1_2_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_5_LC_1_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_5_LC_1_2_7 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst16.count_5_LC_1_2_7  (
            .in0(N__15889),
            .in1(N__15263),
            .in2(N__15294),
            .in3(N__16045),
            .lcout(\b2v_inst16.count_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36601),
            .ce(N__20928),
            .sr(N__20785));
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_1_3_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_LC_1_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__15582),
            .in2(N__15709),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_3_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_3_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_1_c_RNIAGME_LC_1_3_1  (
            .in0(N__16036),
            .in1(N__15519),
            .in2(_gnd_net_),
            .in3(N__14740),
            .lcout(\b2v_inst16.count_rst_7 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_1 ),
            .carryout(\b2v_inst16.un4_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_1_3_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_1_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_2_THRU_LUT4_0_LC_1_3_2  (
            .in0(_gnd_net_),
            .in1(N__15389),
            .in2(_gnd_net_),
            .in3(N__14725),
            .lcout(\b2v_inst16.un4_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_2 ),
            .carryout(\b2v_inst16.un4_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_1_3_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_1_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_THRU_LUT4_0_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__15632),
            .in2(_gnd_net_),
            .in3(N__14722),
            .lcout(\b2v_inst16.un4_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_3 ),
            .carryout(\b2v_inst16.un4_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_1_3_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_1_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_THRU_LUT4_0_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__15265),
            .in2(_gnd_net_),
            .in3(N__14719),
            .lcout(\b2v_inst16.un4_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_4 ),
            .carryout(\b2v_inst16.un4_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_3_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_3_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_5_c_RNIEOQE_LC_1_3_5  (
            .in0(N__16035),
            .in1(N__15564),
            .in2(_gnd_net_),
            .in3(N__14716),
            .lcout(\b2v_inst16.count_rst_11 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_5 ),
            .carryout(\b2v_inst16.un4_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_1_3_6 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_1_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_6_THRU_LUT4_0_LC_1_3_6  (
            .in0(_gnd_net_),
            .in1(N__14843),
            .in2(_gnd_net_),
            .in3(N__14821),
            .lcout(\b2v_inst16.un4_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_6 ),
            .carryout(\b2v_inst16.un4_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_1_3_7 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_1_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_THRU_LUT4_0_LC_1_3_7  (
            .in0(_gnd_net_),
            .in1(N__15348),
            .in2(_gnd_net_),
            .in3(N__14818),
            .lcout(\b2v_inst16.un4_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_7 ),
            .carryout(\b2v_inst16.un4_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_1_4_0 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_1_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_8_THRU_LUT4_0_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__14815),
            .in2(_gnd_net_),
            .in3(N__14785),
            .lcout(\b2v_inst16.un4_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(\b2v_inst16.un4_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_4_1 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_4_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_9_c_RNII0VE_LC_1_4_1  (
            .in0(N__16055),
            .in1(_gnd_net_),
            .in2(N__15540),
            .in3(N__14782),
            .lcout(\b2v_inst16.count_rst ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_9 ),
            .carryout(\b2v_inst16.un4_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_1_4_2 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_1_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_10_THRU_LUT4_0_LC_1_4_2  (
            .in0(_gnd_net_),
            .in1(N__15456),
            .in2(_gnd_net_),
            .in3(N__14767),
            .lcout(\b2v_inst16.un4_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_10 ),
            .carryout(\b2v_inst16.un4_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIFJV31_LC_1_4_3 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIFJV31_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_11_c_RNIFJV31_LC_1_4_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_11_c_RNIFJV31_LC_1_4_3  (
            .in0(N__16056),
            .in1(N__15552),
            .in2(_gnd_net_),
            .in3(N__14764),
            .lcout(\b2v_inst16.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_11 ),
            .carryout(\b2v_inst16.un4_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_4_4 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_4_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_12_c_RNISTM3_LC_1_4_4  (
            .in0(N__16023),
            .in1(N__15360),
            .in2(_gnd_net_),
            .in3(N__14761),
            .lcout(\b2v_inst16.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_12 ),
            .carryout(\b2v_inst16.un4_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_4_5 .C_ON=1'b1;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_4_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_13_c_RNITVN3_LC_1_4_5  (
            .in0(N__16057),
            .in1(N__15397),
            .in2(_gnd_net_),
            .in3(N__14758),
            .lcout(\b2v_inst16.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst16.un4_count_1_cry_13 ),
            .carryout(\b2v_inst16.un4_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_4_6 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_4_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_14_c_RNIU1P3_LC_1_4_6  (
            .in0(N__16024),
            .in1(N__15481),
            .in2(_gnd_net_),
            .in3(N__14755),
            .lcout(\b2v_inst16.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIKN901_12_LC_1_4_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIKN901_12_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIKN901_12_LC_1_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNIKN901_12_LC_1_4_7  (
            .in0(N__20962),
            .in1(N__20913),
            .in2(_gnd_net_),
            .in3(N__20973),
            .lcout(\b2v_inst16.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_2_LC_1_5_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_2_LC_1_5_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_2_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_2_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14874),
            .lcout(\b2v_inst16.count_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36588),
            .ce(N__20943),
            .sr(N__20763));
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_1_6_0 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_1_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_LC_1_6_0 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_LC_1_6_0  (
            .in0(N__15803),
            .in1(N__14923),
            .in2(N__14917),
            .in3(N__15777),
            .lcout(\b2v_inst16.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36585),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI2ABP4_0_LC_1_6_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI2ABP4_0_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI2ABP4_0_LC_1_6_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst16.curr_state_RNI2ABP4_0_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__15757),
            .in2(_gnd_net_),
            .in3(N__36406),
            .lcout(\b2v_inst16.delayed_vddq_pwrgd_en ),
            .ltout(\b2v_inst16.delayed_vddq_pwrgd_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNI8SES8_LC_1_6_2 .C_ON=1'b0;
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNI8SES8_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.delayed_vddq_pwrgd_RNI8SES8_LC_1_6_2 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \b2v_inst16.delayed_vddq_pwrgd_RNI8SES8_LC_1_6_2  (
            .in0(N__14916),
            .in1(N__21202),
            .in2(N__14905),
            .in3(N__15907),
            .lcout(b2v_inst16_un2_vpp_en_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_en_LC_1_6_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_en_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_en_LC_1_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_en_LC_1_6_3  (
            .in0(_gnd_net_),
            .in1(N__36404),
            .in2(_gnd_net_),
            .in3(N__22623),
            .lcout(\b2v_inst200.count_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GPIO_FPGA_SoC_4_ibuf_RNINPGR_LC_1_6_4.C_ON=1'b0;
    defparam GPIO_FPGA_SoC_4_ibuf_RNINPGR_LC_1_6_4.SEQ_MODE=4'b0000;
    defparam GPIO_FPGA_SoC_4_ibuf_RNINPGR_LC_1_6_4.LUT_INIT=16'b0010000000000000;
    LogicCell40 GPIO_FPGA_SoC_4_ibuf_RNINPGR_LC_1_6_4 (
            .in0(N__24390),
            .in1(N__24643),
            .in2(N__24148),
            .in3(N__16102),
            .lcout(N_15_i_0_a4_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_1_6_5 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIKEBL_1_LC_1_6_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \b2v_inst16.curr_state_RNIKEBL_1_LC_1_6_5  (
            .in0(N__15975),
            .in1(N__15802),
            .in2(_gnd_net_),
            .in3(N__36405),
            .lcout(\b2v_inst16.count_en ),
            .ltout(\b2v_inst16.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_1_6_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNID4TJ1_2_LC_1_6_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst16.count_RNID4TJ1_2_LC_1_6_6  (
            .in0(N__14875),
            .in1(_gnd_net_),
            .in2(N__14857),
            .in3(N__14854),
            .lcout(\b2v_inst16.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI_0_LC_1_6_7 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI_0_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI_0_LC_1_6_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst16.curr_state_RNI_0_LC_1_6_7  (
            .in0(N__15976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.N_2987_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI863D_6_LC_1_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI863D_6_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI863D_6_LC_1_7_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \b2v_inst11.count_clk_RNI863D_6_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__24162),
            .in2(_gnd_net_),
            .in3(N__26612),
            .lcout(),
            .ltout(\b2v_inst11.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIDGAL3_0_LC_1_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDGAL3_0_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDGAL3_0_LC_1_7_2 .LUT_INIT=16'b1101110011111111;
    LogicCell40 \b2v_inst11.func_state_RNIDGAL3_0_LC_1_7_2  (
            .in0(N__24389),
            .in1(N__16090),
            .in2(N__14959),
            .in3(N__23904),
            .lcout(),
            .ltout(\b2v_inst11.g1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI24DD8_7_LC_1_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI24DD8_7_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI24DD8_7_LC_1_7_3 .LUT_INIT=16'b0111111101010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI24DD8_7_LC_1_7_3  (
            .in0(N__14947),
            .in1(N__26789),
            .in2(N__14956),
            .in3(N__25859),
            .lcout(\b2v_inst11.dutycycle_RNI24DD8Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIF6NL_7_LC_1_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIF6NL_7_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIF6NL_7_LC_1_7_4 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIF6NL_7_LC_1_7_4  (
            .in0(N__26790),
            .in1(N__23722),
            .in2(N__24166),
            .in3(N__14929),
            .lcout(),
            .ltout(\b2v_inst11.N_7_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI608H1_7_LC_1_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI608H1_7_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI608H1_7_LC_1_7_5 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \b2v_inst11.dutycycle_RNI608H1_7_LC_1_7_5  (
            .in0(N__14941),
            .in1(N__23164),
            .in2(N__14953),
            .in3(N__26611),
            .lcout(),
            .ltout(\b2v_inst11.g2_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIMMPP2_7_LC_1_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIMMPP2_7_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIMMPP2_7_LC_1_7_6 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \b2v_inst11.dutycycle_RNIMMPP2_7_LC_1_7_6  (
            .in0(N__23165),
            .in1(N__26791),
            .in2(N__14950),
            .in3(N__23903),
            .lcout(\b2v_inst11.g2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNINPGR_7_LC_1_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNINPGR_7_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNINPGR_7_LC_1_7_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \b2v_inst11.dutycycle_RNINPGR_7_LC_1_7_7  (
            .in0(N__15919),
            .in1(N__24642),
            .in2(N__26831),
            .in3(N__23166),
            .lcout(\b2v_inst11.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI70K8_0_0_LC_1_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI70K8_0_0_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI70K8_0_0_LC_1_8_2 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \b2v_inst11.func_state_RNI70K8_0_0_LC_1_8_2  (
            .in0(N__23182),
            .in1(N__24387),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.g0_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S3n_ibuf_RNI9HQH3_LC_1_8_7.C_ON=1'b0;
    defparam SLP_S3n_ibuf_RNI9HQH3_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam SLP_S3n_ibuf_RNI9HQH3_LC_1_8_7.LUT_INIT=16'b0111111100110011;
    LogicCell40 SLP_S3n_ibuf_RNI9HQH3_LC_1_8_7 (
            .in0(N__23880),
            .in1(N__33782),
            .in2(N__14989),
            .in3(N__17590),
            .lcout(SLP_S3n_ibuf_RNI9HQHZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_4_LC_1_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_4_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_4_LC_1_9_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \b2v_inst11.count_clk_RNI_4_LC_1_9_0  (
            .in0(N__16287),
            .in1(N__17875),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_1_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_2_LC_1_9_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_2_LC_1_9_1  (
            .in0(N__18430),
            .in1(N__18361),
            .in2(N__14995),
            .in3(N__17904),
            .lcout(\b2v_inst11.N_379 ),
            .ltout(\b2v_inst11.N_379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_1_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_1_LC_1_9_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_1_LC_1_9_2  (
            .in0(N__16374),
            .in1(N__15049),
            .in2(N__14992),
            .in3(N__15019),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_7_LC_1_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_7_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_7_LC_1_9_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst11.count_clk_RNI_7_LC_1_9_3  (
            .in0(N__14980),
            .in1(N__15010),
            .in2(_gnd_net_),
            .in3(N__16572),
            .lcout(\b2v_inst11.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_2_LC_1_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_2_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_2_LC_1_9_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \b2v_inst11.count_clk_RNI_2_LC_1_9_4  (
            .in0(N__16286),
            .in1(N__17903),
            .in2(N__18429),
            .in3(N__18356),
            .lcout(\b2v_inst11.un2_count_clk_17_0_o3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S3n_ibuf_RNIF6NL_LC_1_9_5.C_ON=1'b0;
    defparam SLP_S3n_ibuf_RNIF6NL_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam SLP_S3n_ibuf_RNIF6NL_LC_1_9_5.LUT_INIT=16'b0001000100000000;
    LogicCell40 SLP_S3n_ibuf_RNIF6NL_LC_1_9_5 (
            .in0(N__30295),
            .in1(N__24388),
            .in2(_gnd_net_),
            .in3(N__24127),
            .lcout(SLP_S3n_ibuf_RNIF6NLZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVS8U1_13_LC_1_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVS8U1_13_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVS8U1_13_LC_1_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst11.count_clk_RNIVS8U1_13_LC_1_9_6  (
            .in0(N__15040),
            .in1(N__14979),
            .in2(N__14968),
            .in3(N__15127),
            .lcout(\b2v_inst11.count_clk_RNIVS8U1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINPGR_1_1_LC_1_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINPGR_1_1_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINPGR_1_1_LC_1_9_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \b2v_inst11.func_state_RNINPGR_1_1_LC_1_9_7  (
            .in0(N__24511),
            .in1(N__24212),
            .in2(N__26641),
            .in3(N__16174),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_13_LC_1_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_13_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_13_LC_1_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_13_LC_1_10_0  (
            .in0(N__16567),
            .in1(N__16369),
            .in2(N__18322),
            .in3(N__16445),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_5_LC_1_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_5_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_5_LC_1_10_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_5_LC_1_10_1  (
            .in0(N__18259),
            .in1(N__18320),
            .in2(_gnd_net_),
            .in3(N__16568),
            .lcout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI3BJF_4_LC_1_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI3BJF_4_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI3BJF_4_LC_1_10_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \b2v_inst11.count_clk_RNI3BJF_4_LC_1_10_2  (
            .in0(N__16886),
            .in1(N__16273),
            .in2(N__18084),
            .in3(N__15106),
            .lcout(\b2v_inst11.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVS8U1_14_LC_1_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVS8U1_14_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVS8U1_14_LC_1_10_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \b2v_inst11.count_clk_RNIVS8U1_14_LC_1_10_3  (
            .in0(N__18258),
            .in1(N__16407),
            .in2(N__16222),
            .in3(N__16341),
            .lcout(\b2v_inst11.count_clk_RNIVS8U1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI608H1_1_LC_1_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI608H1_1_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI608H1_1_LC_1_10_4 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \b2v_inst11.func_state_RNI608H1_1_LC_1_10_4  (
            .in0(N__24512),
            .in1(N__23698),
            .in2(N__15034),
            .in3(N__15025),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_13_LC_1_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_13_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_13_LC_1_10_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI_13_LC_1_10_5  (
            .in0(N__16330),
            .in1(N__16406),
            .in2(N__16449),
            .in3(N__15126),
            .lcout(\b2v_inst11.N_175 ),
            .ltout(\b2v_inst11.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_1_LC_1_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_1_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_1_LC_1_10_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \b2v_inst11.count_clk_RNI_1_LC_1_10_6  (
            .in0(N__16368),
            .in1(N__18257),
            .in2(N__15013),
            .in3(N__18316),
            .lcout(\b2v_inst11.N_190 ),
            .ltout(\b2v_inst11.N_190_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_6_LC_1_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_6_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_6_LC_1_10_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \b2v_inst11.count_clk_RNI_6_LC_1_10_7  (
            .in0(N__16566),
            .in1(N__17870),
            .in2(N__15004),
            .in3(N__15001),
            .lcout(\b2v_inst11.N_3038_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_14_LC_1_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_14_LC_1_11_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_14_LC_1_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_14_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16927),
            .lcout(\b2v_inst11.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__18082),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIMATB8_0_LC_1_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIMATB8_0_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIMATB8_0_LC_1_11_1 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \b2v_inst11.func_state_RNIMATB8_0_LC_1_11_1  (
            .in0(N__17959),
            .in1(N__25858),
            .in2(N__23179),
            .in3(N__16078),
            .lcout(\b2v_inst11.count_clk_en ),
            .ltout(\b2v_inst11.count_clk_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI3T3F_13_LC_1_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI3T3F_13_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI3T3F_13_LC_1_11_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst11.count_clk_RNI3T3F_13_LC_1_11_2  (
            .in0(N__16429),
            .in1(_gnd_net_),
            .in2(N__15082),
            .in3(N__15079),
            .lcout(\b2v_inst11.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_13_LC_1_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_13_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_13_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_13_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16428),
            .lcout(\b2v_inst11.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__18082),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_15_LC_1_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_15_LC_1_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_15_LC_1_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_15_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16794),
            .lcout(\b2v_inst11.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__18082),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI736F_15_LC_1_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI736F_15_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI736F_15_LC_1_11_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst11.count_clk_RNI736F_15_LC_1_11_6  (
            .in0(N__18083),
            .in1(_gnd_net_),
            .in2(N__16795),
            .in3(N__15073),
            .lcout(\b2v_inst11.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_2_LC_1_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_2_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_2_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_2_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18384),
            .lcout(\b2v_inst11.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36582),
            .ce(N__18082),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI1Q2F_12_LC_1_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI1Q2F_12_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI1Q2F_12_LC_1_12_0 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \b2v_inst11.count_clk_RNI1Q2F_12_LC_1_12_0  (
            .in0(N__16865),
            .in1(N__18054),
            .in2(N__15067),
            .in3(N__16462),
            .lcout(\b2v_inst11.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_12_LC_1_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_12_LC_1_12_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_12_LC_1_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_clk_12_LC_1_12_1  (
            .in0(N__16461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16870),
            .lcout(\b2v_inst11.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36584),
            .ce(N__18107),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_10_LC_1_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_10_LC_1_12_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_10_LC_1_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_clk_10_LC_1_12_2  (
            .in0(N__16868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16512),
            .lcout(\b2v_inst11.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36584),
            .ce(N__18107),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIMAMA_10_LC_1_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIMAMA_10_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIMAMA_10_LC_1_12_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_clk_RNIMAMA_10_LC_1_12_3  (
            .in0(N__18055),
            .in1(N__15058),
            .in2(N__16516),
            .in3(N__16866),
            .lcout(\b2v_inst11.count_clkZ0Z_10 ),
            .ltout(\b2v_inst11.count_clkZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_15_LC_1_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_15_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_15_LC_1_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI_15_LC_1_12_4  (
            .in0(N__16501),
            .in1(N__16474),
            .in2(N__15052),
            .in3(N__16899),
            .lcout(\b2v_inst11.un2_count_clk_17_0_o2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVM1F_11_LC_1_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVM1F_11_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVM1F_11_LC_1_12_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_clk_RNIVM1F_11_LC_1_12_5  (
            .in0(N__18056),
            .in1(N__15112),
            .in2(N__16489),
            .in3(N__16867),
            .lcout(\b2v_inst11.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_11_LC_1_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_11_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_11_LC_1_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_clk_11_LC_1_12_6  (
            .in0(N__16869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16485),
            .lcout(\b2v_inst11.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36584),
            .ce(N__18107),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_4_LC_1_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_4_LC_1_12_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_4_LC_1_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_clk_4_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(N__16266),
            .in2(_gnd_net_),
            .in3(N__16871),
            .lcout(\b2v_inst11.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36584),
            .ce(N__18107),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_c_LC_1_13_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_c_LC_1_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_c_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__20326),
            .in2(N__18748),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\b2v_inst20.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__18595),
            .in2(_gnd_net_),
            .in3(N__15097),
            .lcout(\b2v_inst20.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_1 ),
            .carryout(\b2v_inst20.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(N__18454),
            .in2(_gnd_net_),
            .in3(N__15094),
            .lcout(\b2v_inst20.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_2 ),
            .carryout(\b2v_inst20.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__18676),
            .in2(_gnd_net_),
            .in3(N__15091),
            .lcout(\b2v_inst20.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_3 ),
            .carryout(\b2v_inst20.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4  (
            .in0(_gnd_net_),
            .in1(N__20374),
            .in2(_gnd_net_),
            .in3(N__15088),
            .lcout(\b2v_inst20.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_4 ),
            .carryout(\b2v_inst20.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst20.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__20350),
            .in2(_gnd_net_),
            .in3(N__15085),
            .lcout(\b2v_inst20.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_5 ),
            .carryout(\b2v_inst20.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_7_LC_1_13_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_7_LC_1_13_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_7_LC_1_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_7_LC_1_13_6  (
            .in0(_gnd_net_),
            .in1(N__20388),
            .in2(_gnd_net_),
            .in3(N__15154),
            .lcout(\b2v_inst20.counterZ0Z_7 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_6 ),
            .carryout(\b2v_inst20.counter_1_cry_7 ),
            .clk(N__36587),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_8_LC_1_13_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_8_LC_1_13_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_8_LC_1_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_8_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__16741),
            .in2(_gnd_net_),
            .in3(N__15151),
            .lcout(\b2v_inst20.counterZ0Z_8 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_7 ),
            .carryout(\b2v_inst20.counter_1_cry_8 ),
            .clk(N__36587),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_9_LC_1_14_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_9_LC_1_14_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_9_LC_1_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_9_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__16768),
            .in2(_gnd_net_),
            .in3(N__15148),
            .lcout(\b2v_inst20.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\b2v_inst20.counter_1_cry_9 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_10_LC_1_14_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_10_LC_1_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_10_LC_1_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_10_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__16755),
            .in2(_gnd_net_),
            .in3(N__15145),
            .lcout(\b2v_inst20.counterZ0Z_10 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_9 ),
            .carryout(\b2v_inst20.counter_1_cry_10 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_11_LC_1_14_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_11_LC_1_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_11_LC_1_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_11_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__16780),
            .in2(_gnd_net_),
            .in3(N__15142),
            .lcout(\b2v_inst20.counterZ0Z_11 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_10 ),
            .carryout(\b2v_inst20.counter_1_cry_11 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_12_LC_1_14_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_12_LC_1_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_12_LC_1_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_12_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(N__16690),
            .in2(_gnd_net_),
            .in3(N__15139),
            .lcout(\b2v_inst20.counterZ0Z_12 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_11 ),
            .carryout(\b2v_inst20.counter_1_cry_12 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_13_LC_1_14_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_13_LC_1_14_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_13_LC_1_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_13_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__16704),
            .in2(_gnd_net_),
            .in3(N__15136),
            .lcout(\b2v_inst20.counterZ0Z_13 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_12 ),
            .carryout(\b2v_inst20.counter_1_cry_13 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_14_LC_1_14_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_14_LC_1_14_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_14_LC_1_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_14_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__16717),
            .in2(_gnd_net_),
            .in3(N__15133),
            .lcout(\b2v_inst20.counterZ0Z_14 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_13 ),
            .carryout(\b2v_inst20.counter_1_cry_14 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_15_LC_1_14_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_15_LC_1_14_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_15_LC_1_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_15_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__16729),
            .in2(_gnd_net_),
            .in3(N__15130),
            .lcout(\b2v_inst20.counterZ0Z_15 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_14 ),
            .carryout(\b2v_inst20.counter_1_cry_15 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_16_LC_1_14_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_16_LC_1_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_16_LC_1_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_16_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__16639),
            .in2(_gnd_net_),
            .in3(N__15181),
            .lcout(\b2v_inst20.counterZ0Z_16 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_15 ),
            .carryout(\b2v_inst20.counter_1_cry_16 ),
            .clk(N__36590),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_17_LC_1_15_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_17_LC_1_15_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_17_LC_1_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_17_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__16666),
            .in2(_gnd_net_),
            .in3(N__15178),
            .lcout(\b2v_inst20.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\b2v_inst20.counter_1_cry_17 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_18_LC_1_15_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_18_LC_1_15_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_18_LC_1_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_18_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__16653),
            .in2(_gnd_net_),
            .in3(N__15175),
            .lcout(\b2v_inst20.counterZ0Z_18 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_17 ),
            .carryout(\b2v_inst20.counter_1_cry_18 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_19_LC_1_15_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_19_LC_1_15_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_19_LC_1_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_19_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__16678),
            .in2(_gnd_net_),
            .in3(N__15172),
            .lcout(\b2v_inst20.counterZ0Z_19 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_18 ),
            .carryout(\b2v_inst20.counter_1_cry_19 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_20_LC_1_15_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_20_LC_1_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_20_LC_1_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_20_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__16588),
            .in2(_gnd_net_),
            .in3(N__15169),
            .lcout(\b2v_inst20.counterZ0Z_20 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_19 ),
            .carryout(\b2v_inst20.counter_1_cry_20 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_21_LC_1_15_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_21_LC_1_15_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_21_LC_1_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_21_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__16615),
            .in2(_gnd_net_),
            .in3(N__15166),
            .lcout(\b2v_inst20.counterZ0Z_21 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_20 ),
            .carryout(\b2v_inst20.counter_1_cry_21 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_22_LC_1_15_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_22_LC_1_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_22_LC_1_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_22_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__16602),
            .in2(_gnd_net_),
            .in3(N__15163),
            .lcout(\b2v_inst20.counterZ0Z_22 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_21 ),
            .carryout(\b2v_inst20.counter_1_cry_22 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_23_LC_1_15_6 .C_ON=1'b1;
    defparam \b2v_inst20.counter_23_LC_1_15_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_23_LC_1_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_23_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__16627),
            .in2(_gnd_net_),
            .in3(N__15160),
            .lcout(\b2v_inst20.counterZ0Z_23 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_22 ),
            .carryout(\b2v_inst20.counter_1_cry_23 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_24_LC_1_15_7 .C_ON=1'b1;
    defparam \b2v_inst20.counter_24_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_24_LC_1_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_24_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__17011),
            .in2(_gnd_net_),
            .in3(N__15157),
            .lcout(\b2v_inst20.counterZ0Z_24 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_23 ),
            .carryout(\b2v_inst20.counter_1_cry_24 ),
            .clk(N__36596),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_25_LC_1_16_0 .C_ON=1'b1;
    defparam \b2v_inst20.counter_25_LC_1_16_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_25_LC_1_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_25_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__17038),
            .in2(_gnd_net_),
            .in3(N__15205),
            .lcout(\b2v_inst20.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\b2v_inst20.counter_1_cry_25 ),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_26_LC_1_16_1 .C_ON=1'b1;
    defparam \b2v_inst20.counter_26_LC_1_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_26_LC_1_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_26_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__17025),
            .in2(_gnd_net_),
            .in3(N__15202),
            .lcout(\b2v_inst20.counterZ0Z_26 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_25 ),
            .carryout(\b2v_inst20.counter_1_cry_26 ),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_27_LC_1_16_2 .C_ON=1'b1;
    defparam \b2v_inst20.counter_27_LC_1_16_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_27_LC_1_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_27_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__17050),
            .in2(_gnd_net_),
            .in3(N__15199),
            .lcout(\b2v_inst20.counterZ0Z_27 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_26 ),
            .carryout(\b2v_inst20.counter_1_cry_27 ),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_28_LC_1_16_3 .C_ON=1'b1;
    defparam \b2v_inst20.counter_28_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_28_LC_1_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_28_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__17068),
            .in2(_gnd_net_),
            .in3(N__15196),
            .lcout(\b2v_inst20.counterZ0Z_28 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_27 ),
            .carryout(\b2v_inst20.counter_1_cry_28 ),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_29_LC_1_16_4 .C_ON=1'b1;
    defparam \b2v_inst20.counter_29_LC_1_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_29_LC_1_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_29_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__17095),
            .in2(_gnd_net_),
            .in3(N__15193),
            .lcout(\b2v_inst20.counterZ0Z_29 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_28 ),
            .carryout(\b2v_inst20.counter_1_cry_29 ),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_30_LC_1_16_5 .C_ON=1'b1;
    defparam \b2v_inst20.counter_30_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_30_LC_1_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst20.counter_30_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__17082),
            .in2(_gnd_net_),
            .in3(N__15190),
            .lcout(\b2v_inst20.counterZ0Z_30 ),
            .ltout(),
            .carryin(\b2v_inst20.counter_1_cry_29 ),
            .carryout(\b2v_inst20.counter_1_cry_30 ),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_31_LC_1_16_6 .C_ON=1'b0;
    defparam \b2v_inst20.counter_31_LC_1_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_31_LC_1_16_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.counter_31_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(N__17107),
            .in2(_gnd_net_),
            .in3(N__15187),
            .lcout(\b2v_inst20.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36600),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_1_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI1I651_0_LC_2_1_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNI1I651_0_LC_2_1_0  (
            .in0(N__15676),
            .in1(N__20932),
            .in2(_gnd_net_),
            .in3(N__15301),
            .lcout(\b2v_inst16.countZ0Z_0 ),
            .ltout(\b2v_inst16.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_0_LC_2_1_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_LC_2_1_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \b2v_inst16.count_RNI_0_LC_2_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15184),
            .in3(N__15727),
            .lcout(\b2v_inst16.N_416 ),
            .ltout(\b2v_inst16.N_416_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_1_2 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_1_2 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_7_c_RNIGSSE_LC_2_1_2  (
            .in0(N__16029),
            .in1(N__15349),
            .in2(N__15325),
            .in3(N__15321),
            .lcout(\b2v_inst16.count_rst_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_0_0_LC_2_1_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_0_0_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_0_0_LC_2_1_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst16.count_RNI_0_0_LC_2_1_3  (
            .in0(N__15698),
            .in1(N__16027),
            .in2(_gnd_net_),
            .in3(N__15726),
            .lcout(\b2v_inst16.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_4_c_RNIDMPE_LC_2_1_4  (
            .in0(N__16028),
            .in1(N__15264),
            .in2(N__15295),
            .in3(N__15886),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst16.count_RNIJD0K1_5_LC_2_1_5  (
            .in0(N__20933),
            .in1(_gnd_net_),
            .in2(N__15274),
            .in3(N__15271),
            .lcout(\b2v_inst16.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_2_1_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_2_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI4M8F1_10_LC_2_1_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNI4M8F1_10_LC_2_1_6  (
            .in0(N__15226),
            .in1(N__20934),
            .in2(_gnd_net_),
            .in3(N__15237),
            .lcout(\b2v_inst16.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_10_LC_2_1_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_10_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_10_LC_2_1_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_10_LC_2_1_7  (
            .in0(N__15238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36615),
            .ce(N__20942),
            .sr(N__20798));
    defparam \b2v_inst16.count_RNILG1K1_6_LC_2_2_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILG1K1_6_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILG1K1_6_LC_2_2_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst16.count_RNILG1K1_6_LC_2_2_0  (
            .in0(N__15211),
            .in1(N__15219),
            .in2(_gnd_net_),
            .in3(N__20938),
            .lcout(\b2v_inst16.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_6_LC_2_2_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_6_LC_2_2_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_6_LC_2_2_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_6_LC_2_2_1  (
            .in0(N__15220),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36610),
            .ce(N__20945),
            .sr(N__20797));
    defparam \b2v_inst16.count_RNILS241_15_LC_2_2_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNILS241_15_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNILS241_15_LC_2_2_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst16.count_RNILS241_15_LC_2_2_2  (
            .in0(N__15433),
            .in1(N__15418),
            .in2(_gnd_net_),
            .in3(N__20939),
            .lcout(\b2v_inst16.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_15_LC_2_2_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_15_LC_2_2_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_15_LC_2_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_15_LC_2_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15432),
            .lcout(\b2v_inst16.count_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36610),
            .ce(N__20945),
            .sr(N__20797));
    defparam \b2v_inst200.count_RNI3TN71_12_LC_2_2_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3TN71_12_LC_2_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNI3TN71_12_LC_2_2_4  (
            .in0(N__25212),
            .in1(N__17143),
            .in2(_gnd_net_),
            .in3(N__18904),
            .lcout(\b2v_inst200.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73351_5_LC_2_2_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73351_5_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73351_5_LC_2_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI73351_5_LC_2_2_5  (
            .in0(N__17128),
            .in1(N__25210),
            .in2(_gnd_net_),
            .in3(N__18802),
            .lcout(\b2v_inst200.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9551_7_LC_2_2_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9551_7_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9551_7_LC_2_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst200.count_RNIB9551_7_LC_2_2_6  (
            .in0(N__25211),
            .in1(N__17119),
            .in2(_gnd_net_),
            .in3(N__18778),
            .lcout(\b2v_inst200.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_14_LC_2_3_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_14_LC_2_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_14_LC_2_3_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst16.count_14_LC_2_3_0  (
            .in0(N__15406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.count_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__20944),
            .sr(N__20796));
    defparam \b2v_inst16.count_RNIJP141_14_LC_2_3_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIJP141_14_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIJP141_14_LC_2_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNIJP141_14_LC_2_3_1  (
            .in0(N__15412),
            .in1(N__20912),
            .in2(_gnd_net_),
            .in3(N__15405),
            .lcout(\b2v_inst16.countZ0Z_14 ),
            .ltout(\b2v_inst16.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_13_LC_2_3_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_13_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_13_LC_2_3_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \b2v_inst16.count_RNI_13_LC_2_3_2  (
            .in0(N__15633),
            .in1(N__15390),
            .in2(N__15364),
            .in3(N__15361),
            .lcout(\b2v_inst16.count_4_i_a3_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIHM041_13_LC_2_3_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIHM041_13_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIHM041_13_LC_2_3_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNIHM041_13_LC_2_3_3  (
            .in0(N__15592),
            .in1(N__20911),
            .in2(_gnd_net_),
            .in3(N__15600),
            .lcout(\b2v_inst16.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_3_4 .C_ON=1'b0;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_3_4 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.un4_count_1_cry_3_c_RNICKOE_LC_2_3_4  (
            .in0(N__15618),
            .in1(N__16025),
            .in2(N__15637),
            .in3(N__15895),
            .lcout(),
            .ltout(\b2v_inst16.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_2_3_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIHAVJ1_4_LC_2_3_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst16.count_RNIHAVJ1_4_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(N__15607),
            .in2(N__15640),
            .in3(N__20910),
            .lcout(\b2v_inst16.countZ0Z_4 ),
            .ltout(\b2v_inst16.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_4_LC_2_3_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_4_LC_2_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_4_LC_2_3_6 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst16.count_4_LC_2_3_6  (
            .in0(N__15619),
            .in1(N__16026),
            .in2(N__15610),
            .in3(N__15896),
            .lcout(\b2v_inst16.count_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__20944),
            .sr(N__20796));
    defparam \b2v_inst16.count_13_LC_2_3_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_13_LC_2_3_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_13_LC_2_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_13_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15601),
            .lcout(\b2v_inst16.count_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36602),
            .ce(N__20944),
            .sr(N__20796));
    defparam \b2v_inst16.count_RNI2J651_0_1_LC_2_4_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2J651_0_1_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2J651_0_1_LC_2_4_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst16.count_RNI2J651_0_1_LC_2_4_0  (
            .in0(N__15502),
            .in1(N__20882),
            .in2(_gnd_net_),
            .in3(N__15490),
            .lcout(\b2v_inst16.un4_count_1_axb_1 ),
            .ltout(\b2v_inst16.un4_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI_1_LC_2_4_1 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI_1_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI_1_LC_2_4_1 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \b2v_inst16.count_RNI_1_LC_2_4_1  (
            .in0(N__15712),
            .in1(_gnd_net_),
            .in2(N__15586),
            .in3(N__15982),
            .lcout(\b2v_inst16.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_1_LC_2_4_2 .C_ON=1'b0;
    defparam \b2v_inst16.count_1_LC_2_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_1_LC_2_4_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst16.count_1_LC_2_4_2  (
            .in0(N__15983),
            .in1(N__15710),
            .in2(_gnd_net_),
            .in3(N__15583),
            .lcout(\b2v_inst16.count_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36597),
            .ce(N__20914),
            .sr(N__20789));
    defparam \b2v_inst16.count_RNIKN901_0_12_LC_2_4_3 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIKN901_0_12_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIKN901_0_12_LC_2_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst16.count_RNIKN901_0_12_LC_2_4_3  (
            .in0(N__15571),
            .in1(N__15553),
            .in2(N__15541),
            .in3(N__15520),
            .lcout(\b2v_inst16.count_4_i_a3_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI2J651_1_LC_2_4_4 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2J651_1_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2J651_1_LC_2_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst16.count_RNI2J651_1_LC_2_4_4  (
            .in0(N__20915),
            .in1(N__15501),
            .in2(_gnd_net_),
            .in3(N__15489),
            .lcout(),
            .ltout(\b2v_inst16.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNI2J651_2_1_LC_2_4_5 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNI2J651_2_1_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNI2J651_2_1_LC_2_4_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst16.count_RNI2J651_2_1_LC_2_4_5  (
            .in0(N__15477),
            .in1(_gnd_net_),
            .in2(N__15463),
            .in3(N__15460),
            .lcout(),
            .ltout(\b2v_inst16.count_4_i_a3_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_RNIMAG52_12_LC_2_4_6 .C_ON=1'b0;
    defparam \b2v_inst16.count_RNIMAG52_12_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.count_RNIMAG52_12_LC_2_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst16.count_RNIMAG52_12_LC_2_4_6  (
            .in0(N__15751),
            .in1(N__15742),
            .in2(N__15736),
            .in3(N__15733),
            .lcout(\b2v_inst16.N_414 ),
            .ltout(\b2v_inst16.N_414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_0_LC_2_4_7 .C_ON=1'b0;
    defparam \b2v_inst16.count_0_LC_2_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_0_LC_2_4_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst16.count_0_LC_2_4_7  (
            .in0(N__15711),
            .in1(_gnd_net_),
            .in2(N__15679),
            .in3(N__15984),
            .lcout(\b2v_inst16.count_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36597),
            .ce(N__20914),
            .sr(N__20789));
    defparam \b2v_inst11.count_off_RNI5BGAF_1_LC_2_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI5BGAF_1_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI5BGAF_1_LC_2_5_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.count_off_RNI5BGAF_1_LC_2_5_0  (
            .in0(N__19318),
            .in1(N__15655),
            .in2(N__19485),
            .in3(N__15664),
            .lcout(\b2v_inst11.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4AGAF_0_LC_2_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4AGAF_0_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4AGAF_0_LC_2_5_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst11.count_off_RNI4AGAF_0_LC_2_5_1  (
            .in0(N__17170),
            .in1(N__19431),
            .in2(N__15649),
            .in3(N__19317),
            .lcout(\b2v_inst11.count_offZ0Z_0 ),
            .ltout(\b2v_inst11.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_1_LC_2_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_1_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_1_LC_2_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.count_off_RNI_1_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15667),
            .in3(N__19145),
            .lcout(\b2v_inst11.count_off_RNIZ0Z_1 ),
            .ltout(\b2v_inst11.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_1_LC_2_5_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_1_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_1_LC_2_5_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.count_off_1_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15658),
            .in3(N__19323),
            .lcout(\b2v_inst11.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36592),
            .ce(N__19484),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_0_LC_2_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_0_LC_2_5_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_0_LC_2_5_4 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \b2v_inst11.count_off_0_LC_2_5_4  (
            .in0(N__19320),
            .in1(N__17171),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36592),
            .ce(N__19484),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_10_LC_2_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_10_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_10_LC_2_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_10_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__17241),
            .in2(_gnd_net_),
            .in3(N__19321),
            .lcout(\b2v_inst11.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36592),
            .ce(N__19484),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIRKFDF_10_LC_2_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIRKFDF_10_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIRKFDF_10_LC_2_5_6 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \b2v_inst11.count_off_RNIRKFDF_10_LC_2_5_6  (
            .in0(N__19319),
            .in1(N__15913),
            .in2(N__19486),
            .in3(N__17242),
            .lcout(\b2v_inst11.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_13_LC_2_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_13_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_13_LC_2_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_13_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(N__17373),
            .in2(_gnd_net_),
            .in3(N__19322),
            .lcout(\b2v_inst11.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36592),
            .ce(N__19484),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI3B692_0_0_LC_2_6_0 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI3B692_0_0_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI3B692_0_0_LC_2_6_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \b2v_inst16.curr_state_RNI3B692_0_0_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__15773),
            .in2(_gnd_net_),
            .in3(N__15807),
            .lcout(\b2v_inst16.N_1440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI3B692_0_LC_2_6_1 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI3B692_0_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI3B692_0_LC_2_6_1 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \b2v_inst16.curr_state_RNI3B692_0_LC_2_6_1  (
            .in0(N__21140),
            .in1(N__35904),
            .in2(N__15811),
            .in3(N__15817),
            .lcout(\b2v_inst16.curr_state_RNI3B692Z0Z_0 ),
            .ltout(\b2v_inst16.curr_state_RNI3B692Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_1_LC_2_6_2 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_1_LC_2_6_2 .LUT_INIT=16'b0100000011101010;
    LogicCell40 \b2v_inst16.curr_state_1_LC_2_6_2  (
            .in0(N__15809),
            .in1(N__21142),
            .in2(N__15901),
            .in3(N__15897),
            .lcout(\b2v_inst16.curr_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36589),
            .ce(N__36369),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIERV34_0_0_LC_2_6_3 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIERV34_0_0_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIERV34_0_0_LC_2_6_3 .LUT_INIT=16'b1100110001011111;
    LogicCell40 \b2v_inst16.curr_state_RNIERV34_0_0_LC_2_6_3  (
            .in0(N__21139),
            .in1(N__15894),
            .in2(N__15778),
            .in3(N__15810),
            .lcout(),
            .ltout(\b2v_inst16.curr_state_7_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI7NCI4_1_LC_2_6_4 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI7NCI4_1_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI7NCI4_1_LC_2_6_4 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \b2v_inst16.curr_state_RNI7NCI4_1_LC_2_6_4  (
            .in0(N__35903),
            .in1(_gnd_net_),
            .in2(N__15829),
            .in3(N__15826),
            .lcout(\b2v_inst16.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst16.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_0_LC_2_6_5 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_0_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst16.curr_state_0_LC_2_6_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \b2v_inst16.curr_state_0_LC_2_6_5  (
            .in0(N__21141),
            .in1(_gnd_net_),
            .in2(N__15820),
            .in3(_gnd_net_),
            .lcout(\b2v_inst16.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36589),
            .ce(N__36369),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNIERV34_0_LC_2_6_6 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNIERV34_0_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNIERV34_0_LC_2_6_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \b2v_inst16.curr_state_RNIERV34_0_LC_2_6_6  (
            .in0(N__15808),
            .in1(N__15772),
            .in2(_gnd_net_),
            .in3(N__21138),
            .lcout(\b2v_inst16.N_268 ),
            .ltout(\b2v_inst16.N_268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_RNI68A74_0_LC_2_6_7 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_RNI68A74_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_RNI68A74_0_LC_2_6_7 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \b2v_inst16.curr_state_RNI68A74_0_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16060),
            .in3(N__35902),
            .lcout(\b2v_inst16.N_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNILCR74_0_LC_2_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNILCR74_0_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNILCR74_0_LC_2_7_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \b2v_inst11.func_state_RNILCR74_0_LC_2_7_0  (
            .in0(N__16113),
            .in1(N__17834),
            .in2(N__16141),
            .in3(N__16213),
            .lcout(\b2v_inst11.N_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_0_LC_2_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_0_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_0_LC_2_7_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_0_LC_2_7_1  (
            .in0(N__24397),
            .in1(N__24641),
            .in2(_gnd_net_),
            .in3(N__23381),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_2_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_2_7_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_0_LC_2_7_2  (
            .in0(N__21201),
            .in1(N__23704),
            .in2(N__15925),
            .in3(N__17746),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_329_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIF6NL_9_LC_2_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIF6NL_9_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIF6NL_9_LC_2_7_3 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \b2v_inst11.count_off_RNIF6NL_9_LC_2_7_3  (
            .in0(N__24393),
            .in1(N__24149),
            .in2(N__17752),
            .in3(N__23382),
            .lcout(\b2v_inst11.N_340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINPGR_2_1_LC_2_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINPGR_2_1_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINPGR_2_1_LC_2_7_4 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \b2v_inst11.func_state_RNINPGR_2_1_LC_2_7_4  (
            .in0(N__24640),
            .in1(N__24396),
            .in2(N__24161),
            .in3(N__27142),
            .lcout(),
            .ltout(\b2v_inst11.func_state_RNINPGR_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI608H1_0_1_LC_2_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI608H1_0_1_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI608H1_0_1_LC_2_7_5 .LUT_INIT=16'b0000111100011111;
    LogicCell40 \b2v_inst11.func_state_RNI608H1_0_1_LC_2_7_5  (
            .in0(N__23705),
            .in1(N__26632),
            .in2(N__15922),
            .in3(N__23426),
            .lcout(\b2v_inst11.func_state_RNI608H1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_2_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_2_7_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_s_1_LC_2_7_6  (
            .in0(N__24150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24394),
            .lcout(b2v_inst11_dutycycle_1_0_iv_0_o3_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_0_LC_2_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_0_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_0_LC_2_7_7 .LUT_INIT=16'b0011011100111111;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_0_LC_2_7_7  (
            .in0(N__24395),
            .in1(N__24151),
            .in2(N__23720),
            .in3(N__19849),
            .lcout(\b2v_inst11.g0_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_2_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_2_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_1_LC_2_8_0  (
            .in0(N__16114),
            .in1(N__23887),
            .in2(N__18718),
            .in3(N__16189),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_o_N_330_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_2_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_2_8_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_1_LC_2_8_1  (
            .in0(N__23702),
            .in1(N__16084),
            .in2(N__16144),
            .in3(N__16134),
            .lcout(),
            .ltout(\b2v_inst11.un1_func_state25_6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_en_LC_2_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_en_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_en_LC_2_8_2 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \b2v_inst11.count_off_en_LC_2_8_2  (
            .in0(N__17575),
            .in1(N__16123),
            .in2(N__16117),
            .in3(N__27722),
            .lcout(\b2v_inst11.count_off_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIC9BO3_1_LC_2_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIC9BO3_1_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIC9BO3_1_LC_2_8_3 .LUT_INIT=16'b1111111110001100;
    LogicCell40 \b2v_inst11.func_state_RNIC9BO3_1_LC_2_8_3  (
            .in0(N__24469),
            .in1(N__24213),
            .in2(N__35938),
            .in3(N__16195),
            .lcout(\b2v_inst11.N_430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_0_LC_2_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_0_LC_2_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.func_state_RNI_1_0_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__23701),
            .in2(_gnd_net_),
            .in3(N__19841),
            .lcout(\b2v_inst11.func_state_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_1_LC_2_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_1_LC_2_8_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_1_LC_2_8_5  (
            .in0(N__23703),
            .in1(_gnd_net_),
            .in2(N__27149),
            .in3(N__29398),
            .lcout(N_236_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIEJ1N1_0_LC_2_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIEJ1N1_0_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIEJ1N1_0_LC_2_8_6 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \b2v_inst11.func_state_RNIEJ1N1_0_LC_2_8_6  (
            .in0(N__24639),
            .in1(N__18496),
            .in2(N__24519),
            .in3(N__19842),
            .lcout(\b2v_inst11.g1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_2_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_2_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_2_LC_2_8_7  (
            .in0(N__23886),
            .in1(N__18717),
            .in2(N__27148),
            .in3(N__17745),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_331_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIH4KN3_0_LC_2_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIH4KN3_0_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIH4KN3_0_LC_2_9_0 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \b2v_inst11.func_state_RNIH4KN3_0_LC_2_9_0  (
            .in0(N__24606),
            .in1(N__33781),
            .in2(N__16069),
            .in3(N__16162),
            .lcout(\b2v_inst11.count_clk_en_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_0_1_LC_2_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_0_1_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_0_1_LC_2_9_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_0_1_LC_2_9_1  (
            .in0(N__26941),
            .in1(N__23696),
            .in2(N__23390),
            .in3(N__17741),
            .lcout(\b2v_inst11.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIMFI92_1_LC_2_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIMFI92_1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIMFI92_1_LC_2_9_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.count_clk_RNIMFI92_1_LC_2_9_2  (
            .in0(N__17798),
            .in1(N__22496),
            .in2(_gnd_net_),
            .in3(N__16187),
            .lcout(\b2v_inst11.un1_count_off_0_sqmuxa_4_i_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI5M9V2_9_LC_2_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI5M9V2_9_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI5M9V2_9_LC_2_9_3 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \b2v_inst11.count_off_RNI5M9V2_9_LC_2_9_3  (
            .in0(N__23068),
            .in1(N__16204),
            .in2(N__27150),
            .in3(N__17799),
            .lcout(\b2v_inst11.func_state_1_ss0_i_0_o3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI8JP5_1_LC_2_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI8JP5_1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI8JP5_1_LC_2_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.count_clk_RNI8JP5_1_LC_2_9_4  (
            .in0(N__24605),
            .in1(N__16188),
            .in2(N__17751),
            .in3(N__21672),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_1_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_9_LC_2_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_9_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_9_LC_2_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.count_off_RNI_9_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17740),
            .lcout(\b2v_inst11.count_off_RNIZ0Z_9 ),
            .ltout(\b2v_inst11.count_off_RNIZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_1_LC_2_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_1_LC_2_9_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.func_state_RNI_1_1_LC_2_9_6  (
            .in0(N__23695),
            .in1(_gnd_net_),
            .in2(N__16168),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.func_state_RNI_1Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNI_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_3_0_LC_2_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_3_0_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_3_0_LC_2_9_7 .LUT_INIT=16'b0000010100000111;
    LogicCell40 \b2v_inst11.func_state_RNI_3_0_LC_2_9_7  (
            .in0(N__19843),
            .in1(N__23697),
            .in2(N__16165),
            .in3(N__17797),
            .lcout(\b2v_inst11.un1_func_state25_4_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_LC_2_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_LC_2_10_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_LC_2_10_0  (
            .in0(N__16878),
            .in1(N__16370),
            .in2(_gnd_net_),
            .in3(N__16334),
            .lcout(),
            .ltout(\b2v_inst11.count_clk_RNIZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI2UQ9_1_LC_2_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI2UQ9_1_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI2UQ9_1_LC_2_10_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI2UQ9_1_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__16150),
            .in2(N__16156),
            .in3(N__18048),
            .lcout(\b2v_inst11.count_clkZ0Z_1 ),
            .ltout(\b2v_inst11.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_1_LC_2_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_1_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_1_LC_2_10_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst11.count_clk_1_LC_2_10_2  (
            .in0(N__16879),
            .in1(_gnd_net_),
            .in2(N__16153),
            .in3(N__16336),
            .lcout(\b2v_inst11.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36583),
            .ce(N__18118),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_0_LC_2_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_0_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_0_LC_2_10_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.count_clk_0_LC_2_10_3  (
            .in0(N__16335),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16880),
            .lcout(\b2v_inst11.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36583),
            .ce(N__18118),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI1TQ9_0_LC_2_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI1TQ9_0_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI1TQ9_0_LC_2_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_clk_RNI1TQ9_0_LC_2_10_4  (
            .in0(N__18050),
            .in1(N__16246),
            .in2(_gnd_net_),
            .in3(N__16228),
            .lcout(\b2v_inst11.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI9KMF_7_LC_2_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI9KMF_7_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI9KMF_7_LC_2_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI9KMF_7_LC_2_10_5  (
            .in0(N__16543),
            .in1(N__16240),
            .in2(_gnd_net_),
            .in3(N__18049),
            .lcout(\b2v_inst11.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_7_LC_2_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_7_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_7_LC_2_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_7_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16542),
            .lcout(\b2v_inst11.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36583),
            .ce(N__18118),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICQPCF_6_LC_2_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICQPCF_6_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICQPCF_6_LC_2_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_off_RNICQPCF_6_LC_2_10_7  (
            .in0(N__19072),
            .in1(N__19458),
            .in2(_gnd_net_),
            .in3(N__19567),
            .lcout(\b2v_inst11.un3_count_off_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_2_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_2_11_0 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_o3_2_LC_2_11_0  (
            .in0(N__23878),
            .in1(N__24366),
            .in2(_gnd_net_),
            .in3(N__24132),
            .lcout(),
            .ltout(\b2v_inst11.N_168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNICGI84_0_LC_2_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNICGI84_0_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNICGI84_0_LC_2_11_1 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \b2v_inst11.func_state_RNICGI84_0_LC_2_11_1  (
            .in0(N__24500),
            .in1(N__35892),
            .in2(N__16234),
            .in3(N__16381),
            .lcout(\b2v_inst11.func_state_RNICGI84_0_0 ),
            .ltout(\b2v_inst11.func_state_RNICGI84_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_2_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_0_LC_2_11_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_0_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16231),
            .in3(N__16337),
            .lcout(\b2v_inst11.count_clk_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_0_0_LC_2_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_0_0_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_0_0_LC_2_11_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_0_0_LC_2_11_3  (
            .in0(N__26942),
            .in1(N__23365),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.func_state_RNIVS8U1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI505F_14_LC_2_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI505F_14_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI505F_14_LC_2_11_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst11.count_clk_RNI505F_14_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__16926),
            .in2(N__18068),
            .in3(N__16393),
            .lcout(\b2v_inst11.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIN9J12_1_LC_2_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIN9J12_1_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIN9J12_1_LC_2_11_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.func_state_RNIN9J12_1_LC_2_11_5  (
            .in0(N__24211),
            .in1(N__23877),
            .in2(N__24515),
            .in3(N__35891),
            .lcout(\b2v_inst11.N_338 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI608H1_0_LC_2_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI608H1_0_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI608H1_0_LC_2_11_6 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \b2v_inst11.func_state_RNI608H1_0_LC_2_11_6  (
            .in0(N__17750),
            .in1(N__23699),
            .in2(N__19840),
            .in3(N__16387),
            .lcout(\b2v_inst11.un1_count_clk_1_sqmuxa_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_0_1_LC_2_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_0_1_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_0_1_LC_2_11_7 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_0_1_LC_2_11_7  (
            .in0(N__23700),
            .in1(N__23366),
            .in2(N__29400),
            .in3(N__23472),
            .lcout(b2v_inst11_un1_dutycycle_172_m3_amcf1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_2_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_LC_2_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__16375),
            .in2(N__16342),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_2_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_2_12_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5M5_LC_2_12_1  (
            .in0(N__16877),
            .in1(N__18360),
            .in2(_gnd_net_),
            .in3(N__16297),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_1_c_RNIS5MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_1 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_2_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_2_12_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7N5_LC_2_12_2  (
            .in0(N__16872),
            .in1(N__17905),
            .in2(_gnd_net_),
            .in3(N__16294),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_2_c_RNIT7NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_2 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_2_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_2_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9O5_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__16291),
            .in2(_gnd_net_),
            .in3(N__16252),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_3_c_RNIU9OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_3 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_2_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_2_12_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBP5_LC_2_12_4  (
            .in0(N__16873),
            .in1(N__18321),
            .in2(_gnd_net_),
            .in3(N__16249),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_4_c_RNIVBPZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_4 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_2_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_2_12_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQ5_LC_2_12_5  (
            .in0(N__16875),
            .in1(N__17874),
            .in2(_gnd_net_),
            .in3(N__16576),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_5_c_RNI0EQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_5 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_2_12_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_2_12_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GR5_LC_2_12_6  (
            .in0(N__16874),
            .in1(N__16573),
            .in2(_gnd_net_),
            .in3(N__16531),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_6_c_RNI1GRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_6 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_2_12_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_2_12_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_7_c_RNI2IS5_LC_2_12_7  (
            .in0(N__16876),
            .in1(N__18428),
            .in2(_gnd_net_),
            .in3(N__16528),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_7_c_RNI2ISZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_2_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_2_13_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KT5_LC_2_13_0  (
            .in0(N__16885),
            .in1(N__18256),
            .in2(_gnd_net_),
            .in3(N__16525),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_8_c_RNI3KTZ0Z5 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_2_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_2_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MU5_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__16522),
            .in2(_gnd_net_),
            .in3(N__16504),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_9_c_RNI4MUZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_9_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_2_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_2_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AA_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__16500),
            .in2(_gnd_net_),
            .in3(N__16477),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_10_c_RNIC1AAZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_10_cZ0 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_2_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_2_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BA_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__16473),
            .in2(_gnd_net_),
            .in3(N__16453),
            .lcout(\b2v_inst11.un1_count_clk_2_cry_11_c_RNID3BAZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_11 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_2_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_2_13_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_12_c_RNIE5CA_LC_2_13_4  (
            .in0(N__16884),
            .in1(N__16450),
            .in2(_gnd_net_),
            .in3(N__16414),
            .lcout(\b2v_inst11.count_clk_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_12 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_2_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_2_13_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_13_c_RNIF7DA_LC_2_13_5  (
            .in0(N__16887),
            .in1(N__16411),
            .in2(_gnd_net_),
            .in3(N__16906),
            .lcout(\b2v_inst11.count_clk_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_clk_2_cry_13 ),
            .carryout(\b2v_inst11.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_2_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_2_13_6 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \b2v_inst11.un1_count_clk_2_cry_14_c_RNIG9EA_LC_2_13_6  (
            .in0(N__16903),
            .in1(_gnd_net_),
            .in2(N__16888),
            .in3(N__16798),
            .lcout(\b2v_inst11.count_clk_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_9_LC_2_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_9_LC_2_13_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_9_LC_2_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst11.count_clk_9_LC_2_13_7  (
            .in0(N__18279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36591),
            .ce(N__18091),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_2_14_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_RNO_LC_2_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_2_c_RNO_LC_2_14_0  (
            .in0(N__16779),
            .in1(N__16767),
            .in2(N__16756),
            .in3(N__16740),
            .lcout(\b2v_inst20.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_2_14_1 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_RNO_LC_2_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_3_c_RNO_LC_2_14_1  (
            .in0(N__16728),
            .in1(N__16716),
            .in2(N__16705),
            .in3(N__16689),
            .lcout(\b2v_inst20.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_2_14_2 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_RNO_LC_2_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_4_c_RNO_LC_2_14_2  (
            .in0(N__16677),
            .in1(N__16665),
            .in2(N__16654),
            .in3(N__16638),
            .lcout(\b2v_inst20.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_2_14_3 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_RNO_LC_2_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_5_c_RNO_LC_2_14_3  (
            .in0(N__16626),
            .in1(N__16614),
            .in2(N__16603),
            .in3(N__16587),
            .lcout(\b2v_inst20.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_4_1_LC_2_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_4_1_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_4_1_LC_2_14_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_4_1_LC_2_14_5  (
            .in0(N__19947),
            .in1(N__23879),
            .in2(_gnd_net_),
            .in3(N__29388),
            .lcout(func_state_RNIVS8U1_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.un1_vddq_en_LC_2_14_6 .C_ON=1'b0;
    defparam \b2v_inst16.un1_vddq_en_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.un1_vddq_en_LC_2_14_6 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \b2v_inst16.un1_vddq_en_LC_2_14_6  (
            .in0(N__21199),
            .in1(N__16981),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(VDDQ_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_LC_2_15_0 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_0_c_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_LC_2_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__18520),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\b2v_inst20.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_LC_2_15_1 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_1_c_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_LC_2_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__20302),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_0 ),
            .carryout(\b2v_inst20.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_2_c_LC_2_15_2 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_2_c_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_2_c_LC_2_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_2_c_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16957),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_1 ),
            .carryout(\b2v_inst20.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_3_c_LC_2_15_3 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_3_c_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_3_c_LC_2_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_3_c_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16948),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_2 ),
            .carryout(\b2v_inst20.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_4_c_LC_2_15_4 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_4_c_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_4_c_LC_2_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_4_c_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__16939),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_3 ),
            .carryout(\b2v_inst20.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_5_c_LC_2_15_5 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_5_c_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_5_c_LC_2_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_5_c_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__16933),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_4 ),
            .carryout(\b2v_inst20.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_LC_2_15_6 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_6_c_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_LC_2_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_6_c_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__16999),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_5 ),
            .carryout(\b2v_inst20.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_LC_2_15_7 .C_ON=1'b1;
    defparam \b2v_inst20.un4_counter_7_c_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_LC_2_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_7_c_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__17056),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst20.un4_counter_6 ),
            .carryout(b2v_inst20_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_2_16_0.C_ON=1'b0;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_2_16_0.SEQ_MODE=4'b0000;
    defparam b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_2_16_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 b2v_inst20_un4_counter_7_THRU_LUT4_0_LC_2_16_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17110),
            .lcout(b2v_inst20_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_2_16_5 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_7_c_RNO_LC_2_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_7_c_RNO_LC_2_16_5  (
            .in0(N__17106),
            .in1(N__17094),
            .in2(N__17083),
            .in3(N__17067),
            .lcout(\b2v_inst20.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_2_16_6 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_6_c_RNO_LC_2_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst20.un4_counter_6_c_RNO_LC_2_16_6  (
            .in0(N__17049),
            .in1(N__17037),
            .in2(N__17026),
            .in3(N__17010),
            .lcout(\b2v_inst20.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_1_LC_4_1_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_1_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_1_LC_4_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst200.count_RNI_1_LC_4_1_0  (
            .in0(N__18829),
            .in1(N__18853),
            .in2(N__18571),
            .in3(N__18544),
            .lcout(\b2v_inst200.un25_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIP16E1_1_LC_4_1_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIP16E1_1_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIP16E1_1_LC_4_1_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNIP16E1_1_LC_4_1_1  (
            .in0(N__18555),
            .in1(N__16993),
            .in2(_gnd_net_),
            .in3(N__25206),
            .lcout(\b2v_inst200.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_1_LC_4_1_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_1_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_1_LC_4_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_1_LC_4_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18556),
            .lcout(\b2v_inst200.count_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36627),
            .ce(N__25154),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QV41_2_LC_4_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QV41_2_LC_4_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNI1QV41_2_LC_4_1_3  (
            .in0(N__16987),
            .in1(N__18531),
            .in2(_gnd_net_),
            .in3(N__25207),
            .lcout(\b2v_inst200.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_2_LC_4_1_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_2_LC_4_1_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_2_LC_4_1_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_2_LC_4_1_4  (
            .in0(N__18532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36627),
            .ce(N__25154),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI3T051_3_LC_4_1_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI3T051_3_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI3T051_3_LC_4_1_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI3T051_3_LC_4_1_5  (
            .in0(N__17149),
            .in1(N__25208),
            .in2(_gnd_net_),
            .in3(N__18840),
            .lcout(\b2v_inst200.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_3_LC_4_1_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_3_LC_4_1_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_3_LC_4_1_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst200.count_3_LC_4_1_6  (
            .in0(N__18841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36627),
            .ce(N__25154),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50251_4_LC_4_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50251_4_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50251_4_LC_4_1_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI50251_4_LC_4_1_7  (
            .in0(N__17134),
            .in1(N__25209),
            .in2(_gnd_net_),
            .in3(N__18816),
            .lcout(\b2v_inst200.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_12_LC_4_2_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_12_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_12_LC_4_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_12_LC_4_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18903),
            .lcout(\b2v_inst200.count_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36623),
            .ce(N__25153),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_13_LC_4_2_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_13_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_13_LC_4_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_13_LC_4_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20644),
            .lcout(\b2v_inst200.count_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36623),
            .ce(N__25153),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_4_LC_4_2_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_4_LC_4_2_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_4_LC_4_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_4_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18817),
            .lcout(\b2v_inst200.count_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36623),
            .ce(N__25153),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_5_LC_4_2_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_5_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_5_LC_4_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_5_LC_4_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18798),
            .lcout(\b2v_inst200.count_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36623),
            .ce(N__25153),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_7_LC_4_2_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_7_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_7_LC_4_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_7_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18774),
            .lcout(\b2v_inst200.count_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36623),
            .ce(N__25153),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_17_LC_4_2_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_17_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_17_LC_4_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_17_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18865),
            .lcout(\b2v_inst200.count_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36623),
            .ce(N__25153),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICFRGF_15_LC_4_3_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICFRGF_15_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICFRGF_15_LC_4_3_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_off_RNICFRGF_15_LC_4_3_0  (
            .in0(N__19533),
            .in1(N__17221),
            .in2(N__19351),
            .in3(N__17328),
            .lcout(\b2v_inst11.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_15_LC_4_3_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_15_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_15_LC_4_3_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.count_off_15_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17332),
            .in3(N__19347),
            .lcout(\b2v_inst11.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36617),
            .ce(N__19536),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI89PGF_13_LC_4_3_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI89PGF_13_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI89PGF_13_LC_4_3_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst11.count_off_RNI89PGF_13_LC_4_3_2  (
            .in0(N__19531),
            .in1(N__17215),
            .in2(N__17377),
            .in3(N__19348),
            .lcout(\b2v_inst11.count_offZ0Z_13 ),
            .ltout(\b2v_inst11.count_offZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI_15_LC_4_3_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI_15_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI_15_LC_4_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_off_RNI_15_LC_4_3_3  (
            .in0(N__18934),
            .in1(N__17191),
            .in2(N__17203),
            .in3(N__17346),
            .lcout(\b2v_inst11.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_8_LC_4_3_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_8_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_8_LC_4_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_8_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__17256),
            .in2(_gnd_net_),
            .in3(N__19350),
            .lcout(\b2v_inst11.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36617),
            .ce(N__19536),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIG0SCF_8_LC_4_3_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIG0SCF_8_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIG0SCF_8_LC_4_3_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \b2v_inst11.count_off_RNIG0SCF_8_LC_4_3_5  (
            .in0(N__19349),
            .in1(N__17200),
            .in2(N__17260),
            .in3(N__19532),
            .lcout(\b2v_inst11.count_offZ0Z_8 ),
            .ltout(\b2v_inst11.count_offZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIETQCF_0_7_LC_4_3_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIETQCF_0_7_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIETQCF_0_7_LC_4_3_6 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \b2v_inst11.count_off_RNIETQCF_0_7_LC_4_3_6  (
            .in0(N__19549),
            .in1(N__19534),
            .in2(N__17194),
            .in3(N__19216),
            .lcout(\b2v_inst11.un34_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIETQCF_7_LC_4_3_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIETQCF_7_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIETQCF_7_LC_4_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_off_RNIETQCF_7_LC_4_3_7  (
            .in0(N__19535),
            .in1(N__19548),
            .in2(_gnd_net_),
            .in3(N__19215),
            .lcout(\b2v_inst11.un3_count_off_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_4_4_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_LC_4_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__19149),
            .in2(N__17190),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_4_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_4_4_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_4_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_RNIU152_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__18913),
            .in2(_gnd_net_),
            .in3(N__17155),
            .lcout(\b2v_inst11.un3_count_off_1_cry_1_c_RNIUZ0Z152 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_1 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_4_4_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_4_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_2_c_RNIV362_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__19012),
            .in2(_gnd_net_),
            .in3(N__17152),
            .lcout(\b2v_inst11.un3_count_off_1_cry_2_c_RNIVZ0Z362 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_2 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_4_4_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_4_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_3_c_RNI0672_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__19006),
            .in2(_gnd_net_),
            .in3(N__17302),
            .lcout(\b2v_inst11.un3_count_off_1_cry_3_c_RNIZ0Z0672 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_3 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_4_4_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_4_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_4_c_RNI1882_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(N__19164),
            .in2(_gnd_net_),
            .in3(N__17299),
            .lcout(\b2v_inst11.un3_count_off_1_cry_4_c_RNIZ0Z1882 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_4 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_4_4_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_4_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_5_c_RNI2A92_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(N__17296),
            .in2(_gnd_net_),
            .in3(N__17281),
            .lcout(\b2v_inst11.un3_count_off_1_cry_5_c_RNI2AZ0Z92 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_5 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_4_4_6 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_4_4_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_6_c_RNI3CA2_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17278),
            .in3(N__17269),
            .lcout(\b2v_inst11.un3_count_off_1_cry_6_c_RNI3CAZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_6 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_4_4_7 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_4_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_7_c_RNI4EB2_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__17266),
            .in2(_gnd_net_),
            .in3(N__17248),
            .lcout(\b2v_inst11.un3_count_off_1_cry_7_c_RNI4EBZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_7 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_4_5_0 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_4_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_8_c_RNI5GC2_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__19021),
            .in2(_gnd_net_),
            .in3(N__17245),
            .lcout(\b2v_inst11.un3_count_off_1_cry_8_c_RNI5GCZ0Z2 ),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\b2v_inst11.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_4_5_1 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_4_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_9_c_RNI6ID2_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__17454),
            .in2(_gnd_net_),
            .in3(N__17227),
            .lcout(\b2v_inst11.un3_count_off_1_cry_9_c_RNI6IDZ0Z2 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_9 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_4_5_2 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_4_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_10_c_RNIEVK5_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__17317),
            .in2(_gnd_net_),
            .in3(N__17224),
            .lcout(\b2v_inst11.un3_count_off_1_cry_10_c_RNIEVKZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_10 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_4_5_3 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_4_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_11_c_RNIF1M5_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__17472),
            .in2(_gnd_net_),
            .in3(N__17389),
            .lcout(\b2v_inst11.un3_count_off_1_cry_11_c_RNIF1MZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_11 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_4_5_4 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_4_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_12_c_RNIG3N5_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__17386),
            .in2(_gnd_net_),
            .in3(N__17356),
            .lcout(\b2v_inst11.un3_count_off_1_cry_12_c_RNIG3NZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_12 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_4_5_5 .C_ON=1'b1;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_4_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_13_c_RNIH5O5_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__18933),
            .in2(_gnd_net_),
            .in3(N__17353),
            .lcout(\b2v_inst11.un3_count_off_1_cry_13_c_RNIH5OZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un3_count_off_1_cry_13 ),
            .carryout(\b2v_inst11.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_4_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_4_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_14_c_RNII7P5_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__17350),
            .in2(_gnd_net_),
            .in3(N__17335),
            .lcout(\b2v_inst11.un3_count_off_1_cry_14_c_RNII7PZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIJE0A4_LC_4_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIJE0A4_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_1_c_RNIJE0A4_LC_4_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_1_c_RNIJE0A4_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(N__19186),
            .in2(_gnd_net_),
            .in3(N__19343),
            .lcout(\b2v_inst11.count_off_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_12_LC_4_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_12_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_12_LC_4_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_12_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__17493),
            .in2(_gnd_net_),
            .in3(N__19341),
            .lcout(\b2v_inst11.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36599),
            .ce(N__19517),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI43NGF_11_LC_4_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI43NGF_11_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI43NGF_11_LC_4_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_off_RNI43NGF_11_LC_4_6_1  (
            .in0(N__17311),
            .in1(N__17409),
            .in2(_gnd_net_),
            .in3(N__19516),
            .lcout(\b2v_inst11.un3_count_off_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI3CGD4_LC_4_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI3CGD4_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_10_c_RNI3CGD4_LC_4_6_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_10_c_RNI3CGD4_LC_4_6_2  (
            .in0(N__17419),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19342),
            .lcout(\b2v_inst11.count_off_1_11 ),
            .ltout(\b2v_inst11.count_off_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI43NGF_0_11_LC_4_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI43NGF_0_11_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI43NGF_0_11_LC_4_6_3 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \b2v_inst11.count_off_RNI43NGF_0_11_LC_4_6_3  (
            .in0(N__17473),
            .in1(N__17410),
            .in2(N__17305),
            .in3(N__19518),
            .lcout(\b2v_inst11.un34_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI66OGF_12_LC_4_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI66OGF_12_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI66OGF_12_LC_4_6_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.count_off_RNI66OGF_12_LC_4_6_4  (
            .in0(N__19515),
            .in1(N__17494),
            .in2(N__17482),
            .in3(N__19339),
            .lcout(\b2v_inst11.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNII3TCF_0_9_LC_4_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNII3TCF_0_9_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNII3TCF_0_9_LC_4_6_5 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \b2v_inst11.count_off_RNII3TCF_0_9_LC_4_6_5  (
            .in0(N__19036),
            .in1(N__19042),
            .in2(N__17461),
            .in3(N__19519),
            .lcout(),
            .ltout(\b2v_inst11.un34_clk_100khz_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIQTKGS2_9_LC_4_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIQTKGS2_9_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIQTKGS2_9_LC_4_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_off_RNIQTKGS2_9_LC_4_6_6  (
            .in0(N__17437),
            .in1(N__19099),
            .in2(N__17431),
            .in3(N__17428),
            .lcout(\b2v_inst11.count_off_RNIQTKGS2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_11_LC_4_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_11_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_11_LC_4_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_11_LC_4_6_7  (
            .in0(N__19340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17418),
            .lcout(\b2v_inst11.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36599),
            .ce(N__19517),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_7_LC_4_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_7_LC_4_7_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_7_LC_4_7_0 .LUT_INIT=16'b1010001100110011;
    LogicCell40 \b2v_inst11.dutycycle_7_LC_4_7_0  (
            .in0(N__17554),
            .in1(N__17395),
            .in2(N__23043),
            .in3(N__17539),
            .lcout(\b2v_inst11.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36594),
            .ce(),
            .sr(N__25981));
    defparam \b2v_inst11.dutycycle_RNI863D_2_LC_4_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI863D_2_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI863D_2_LC_4_7_1 .LUT_INIT=16'b0111011101011111;
    LogicCell40 \b2v_inst11.dutycycle_RNI863D_2_LC_4_7_1  (
            .in0(N__24103),
            .in1(N__23694),
            .in2(N__27151),
            .in3(N__30298),
            .lcout(),
            .ltout(\b2v_inst11.g4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIGT0G4_2_LC_4_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIGT0G4_2_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIGT0G4_2_LC_4_7_2 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \b2v_inst11.dutycycle_RNIGT0G4_2_LC_4_7_2  (
            .in0(N__22991),
            .in1(N__24622),
            .in2(N__17401),
            .in3(N__33784),
            .lcout(\b2v_inst11.g1_0_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIVTQU_LC_4_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIVTQU_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIVTQU_LC_4_7_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIVTQU_LC_4_7_3  (
            .in0(N__24392),
            .in1(N__21481),
            .in2(N__24128),
            .in3(N__23693),
            .lcout(),
            .ltout(\b2v_inst11.g0_17_N_3L3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIVGS13_7_LC_4_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIVGS13_7_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIVGS13_7_LC_4_7_4 .LUT_INIT=16'b0001101110111011;
    LogicCell40 \b2v_inst11.dutycycle_RNIVGS13_7_LC_4_7_4  (
            .in0(N__27724),
            .in1(N__17553),
            .in2(N__17398),
            .in3(N__23894),
            .lcout(\b2v_inst11.dutycycle_RNIVGS13Z0Z_7 ),
            .ltout(\b2v_inst11.dutycycle_RNIVGS13Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIJI0UD_7_LC_4_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIJI0UD_7_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIJI0UD_7_LC_4_7_5 .LUT_INIT=16'b1000101100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNIJI0UD_7_LC_4_7_5  (
            .in0(N__17552),
            .in1(N__17538),
            .in2(N__17524),
            .in3(N__22987),
            .lcout(\b2v_inst11.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_ss0_i_0_x2_LC_4_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_ss0_i_0_x2_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_1_ss0_i_0_x2_LC_4_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.func_state_1_ss0_i_0_x2_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(N__24391),
            .in2(_gnd_net_),
            .in3(N__24104),
            .lcout(\b2v_inst11.N_160_i ),
            .ltout(\b2v_inst11.N_160_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_5_1_LC_4_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_5_1_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_5_1_LC_4_7_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_5_1_LC_4_7_7  (
            .in0(N__23895),
            .in1(N__23376),
            .in2(N__17521),
            .in3(N__17842),
            .lcout(\b2v_inst11.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_1_LC_4_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_1_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_1_LC_4_8_0 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_1_LC_4_8_0  (
            .in0(N__23714),
            .in1(N__23482),
            .in2(N__23907),
            .in3(N__21419),
            .lcout(\b2v_inst11.N_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_4_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_3_LC_4_8_1 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_3_LC_4_8_1  (
            .in0(N__28756),
            .in1(N__21602),
            .in2(N__29539),
            .in3(N__26977),
            .lcout(g0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIUPHS3_6_LC_4_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIUPHS3_6_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIUPHS3_6_LC_4_8_2 .LUT_INIT=16'b0101010111111100;
    LogicCell40 \b2v_inst11.dutycycle_RNIUPHS3_6_LC_4_8_2  (
            .in0(N__17560),
            .in1(N__25840),
            .in2(N__19195),
            .in3(N__19639),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIERM9C_2_LC_4_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIERM9C_2_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIERM9C_2_LC_4_8_3 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \b2v_inst11.dutycycle_RNIERM9C_2_LC_4_8_3  (
            .in0(N__22986),
            .in1(N__17518),
            .in2(N__17509),
            .in3(N__33783),
            .lcout(\b2v_inst11.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_4_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_8_LC_4_8_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_8_LC_4_8_4  (
            .in0(N__26188),
            .in1(N__26329),
            .in2(_gnd_net_),
            .in3(N__29526),
            .lcout(\b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNISM1B4_6_LC_4_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNISM1B4_6_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNISM1B4_6_LC_4_8_5 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNISM1B4_6_LC_4_8_5  (
            .in0(N__18508),
            .in1(N__17506),
            .in2(N__26197),
            .in3(N__23899),
            .lcout(\b2v_inst11.N_231_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_3_LC_4_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_3_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_3_LC_4_8_6 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_3_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28758),
            .in3(N__29525),
            .lcout(\b2v_inst11.N_354 ),
            .ltout(\b2v_inst11.N_354_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_1_LC_4_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_1_LC_4_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_1_LC_4_8_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_1_LC_4_8_7  (
            .in0(N__29399),
            .in1(N__21603),
            .in2(N__17593),
            .in3(N__26976),
            .lcout(b2v_inst11_g0_i_m2_i_a6_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_LC_4_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_LC_4_9_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_LC_4_9_0  (
            .in0(N__23356),
            .in1(N__19728),
            .in2(N__19847),
            .in3(N__20038),
            .lcout(\b2v_inst11.N_159 ),
            .ltout(\b2v_inst11.N_159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_6_0_LC_4_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_6_0_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_6_0_LC_4_9_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.func_state_RNI_6_0_LC_4_9_1  (
            .in0(N__20695),
            .in1(_gnd_net_),
            .in2(N__17581),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI7J1P_0_LC_4_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI7J1P_0_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI7J1P_0_LC_4_9_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst11.func_state_RNI7J1P_0_LC_4_9_2  (
            .in0(N__24361),
            .in1(N__24052),
            .in2(N__19848),
            .in3(N__35897),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m0_0_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIT2K23_1_LC_4_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIT2K23_1_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIT2K23_1_LC_4_9_3 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \b2v_inst11.func_state_RNIT2K23_1_LC_4_9_3  (
            .in0(N__17727),
            .in1(N__22498),
            .in2(N__17578),
            .in3(N__23716),
            .lcout(\b2v_inst11.func_state_1_m0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_4_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_4_9_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst11.un1_func_state25_6_0_o_b2v_inst11_un1_func_state25_6_0_a3_LC_4_9_4  (
            .in0(N__27064),
            .in1(N__20697),
            .in2(N__26947),
            .in3(N__20040),
            .lcout(\b2v_inst11.un1_func_state25_6_0_o_N_313_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI_0_6_LC_4_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI_0_6_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI_0_6_LC_4_9_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_clk_RNI_0_6_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__27063),
            .in2(_gnd_net_),
            .in3(N__26587),
            .lcout(\b2v_inst11.N_19_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIF6NL_6_LC_4_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIF6NL_6_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIF6NL_6_LC_4_9_6 .LUT_INIT=16'b1010101110101111;
    LogicCell40 \b2v_inst11.count_clk_RNIF6NL_6_LC_4_9_6  (
            .in0(N__23499),
            .in1(N__20696),
            .in2(N__26633),
            .in3(N__20039),
            .lcout(),
            .ltout(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIVS8U1_6_LC_4_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIVS8U1_6_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIVS8U1_6_LC_4_9_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \b2v_inst11.count_clk_RNIVS8U1_6_LC_4_9_7  (
            .in0(N__22036),
            .in1(N__20293),
            .in2(N__17563),
            .in3(N__22120),
            .lcout(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_5_1_LC_4_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_5_1_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_5_1_LC_4_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_5_1_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__24190),
            .in2(_gnd_net_),
            .in3(N__23322),
            .lcout(\b2v_inst11.func_state_RNI_5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_2_1_LC_4_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_2_1_LC_4_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNI_2_1_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23638),
            .lcout(\b2v_inst11.func_state_RNI_2Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNI_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_4_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_6_LC_4_10_2 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_6_LC_4_10_2  (
            .in0(N__27102),
            .in1(N__20694),
            .in2(N__17638),
            .in3(N__19726),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m2s2_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICME96_6_LC_4_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICME96_6_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICME96_6_LC_4_10_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \b2v_inst11.dutycycle_RNICME96_6_LC_4_10_3  (
            .in0(N__23060),
            .in1(N__17635),
            .in2(N__17623),
            .in3(N__17620),
            .lcout(\b2v_inst11.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_6_LC_4_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_6_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_6_LC_4_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_6_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__19727),
            .in2(_gnd_net_),
            .in3(N__20693),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_5Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIOSKL1_6_LC_4_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIOSKL1_6_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIOSKL1_6_LC_4_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIOSKL1_6_LC_4_10_5  (
            .in0(N__21665),
            .in1(N__24102),
            .in2(N__17608),
            .in3(N__23852),
            .lcout(),
            .ltout(\b2v_inst11.N_306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIH3TI8_6_LC_4_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIH3TI8_6_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIH3TI8_6_LC_4_10_6 .LUT_INIT=16'b0000010011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIH3TI8_6_LC_4_10_6  (
            .in0(N__19738),
            .in1(N__17605),
            .in2(N__17596),
            .in3(N__23059),
            .lcout(\b2v_inst11.dutycycle_e_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_1_1_LC_4_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_1_1_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_1_1_LC_4_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_1_1_LC_4_10_7  (
            .in0(N__23125),
            .in1(N__23639),
            .in2(N__23519),
            .in3(N__26568),
            .lcout(\b2v_inst11.un1_clk_100khz_43_and_i_0_ccf1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI5M9V2_0_LC_4_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI5M9V2_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI5M9V2_0_LC_4_11_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \b2v_inst11.func_state_RNI5M9V2_0_LC_4_11_0  (
            .in0(N__17763),
            .in1(N__22483),
            .in2(N__23375),
            .in3(N__19760),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m2_am_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIR5S85_1_LC_4_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIR5S85_1_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIR5S85_1_LC_4_11_1 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \b2v_inst11.func_state_RNIR5S85_1_LC_4_11_1  (
            .in0(N__17841),
            .in1(N__23061),
            .in2(N__17809),
            .in3(N__17806),
            .lcout(),
            .ltout(\b2v_inst11.func_state_RNIR5S85Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIMLUM9_0_LC_4_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIMLUM9_0_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIMLUM9_0_LC_4_11_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \b2v_inst11.func_state_RNIMLUM9_0_LC_4_11_2  (
            .in0(N__17661),
            .in1(_gnd_net_),
            .in2(N__17782),
            .in3(N__19879),
            .lcout(\b2v_inst11.func_state_1_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI7762C_0_LC_4_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI7762C_0_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI7762C_0_LC_4_11_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \b2v_inst11.func_state_RNI7762C_0_LC_4_11_3  (
            .in0(N__17948),
            .in1(N__21164),
            .in2(N__17776),
            .in3(N__17646),
            .lcout(\b2v_inst11.func_state ),
            .ltout(\b2v_inst11.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_2_0_LC_4_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_2_0_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_2_0_LC_4_11_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.func_state_RNI_2_0_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17779),
            .in3(_gnd_net_),
            .lcout(func_state_RNI_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_LC_4_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_LC_4_11_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_0_LC_4_11_5 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.func_state_0_LC_4_11_5  (
            .in0(N__17775),
            .in1(N__21165),
            .in2(N__17955),
            .in3(N__17647),
            .lcout(\b2v_inst11.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36593),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_0_0_LC_4_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_0_0_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_0_0_LC_4_11_6 .LUT_INIT=16'b0101011111111111;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_0_0_LC_4_11_6  (
            .in0(N__17764),
            .in1(N__17736),
            .in2(N__17662),
            .in3(N__19761),
            .lcout(),
            .ltout(\b2v_inst11.func_state_1_m2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIOIMG7_1_LC_4_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIOIMG7_1_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIOIMG7_1_LC_4_11_7 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \b2v_inst11.func_state_RNIOIMG7_1_LC_4_11_7  (
            .in0(N__19896),
            .in1(N__17674),
            .in2(N__17665),
            .in3(N__17657),
            .lcout(\b2v_inst11.func_state_1_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_1_LC_4_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_1_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.func_state_1_LC_4_12_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst11.func_state_1_LC_4_12_0  (
            .in0(N__21177),
            .in1(N__17947),
            .in2(N__17971),
            .in3(N__17923),
            .lcout(\b2v_inst11.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36598),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_4_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_4_12_1 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_0_o3_1_LC_4_12_1  (
            .in0(N__22035),
            .in1(N__20289),
            .in2(N__23532),
            .in3(N__22114),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_0_o3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_fast_RNITMQQ5_LC_4_12_2 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_RNITMQQ5_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_fast_RNITMQQ5_LC_4_12_2 .LUT_INIT=16'b1101110111111100;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_RNITMQQ5_LC_4_12_2  (
            .in0(N__27163),
            .in1(N__19988),
            .in2(N__17986),
            .in3(N__19964),
            .lcout(N_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_1_1_LC_4_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_1_1_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_1_1_LC_4_12_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_1_1_LC_4_12_3  (
            .in0(N__26634),
            .in1(N__23857),
            .in2(N__23533),
            .in3(N__23632),
            .lcout(\b2v_inst11.N_326_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_en_0_LC_4_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_en_0_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_en_0_LC_4_12_4 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \b2v_inst11.count_clk_en_0_LC_4_12_4  (
            .in0(N__24920),
            .in1(N__24845),
            .in2(N__24101),
            .in3(N__33725),
            .lcout(\b2v_inst11.count_clk_enZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_4_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.VCCST_EN_i_0_o3_0_LC_4_12_5 .LUT_INIT=16'b0001111111011111;
    LogicCell40 \b2v_inst11.VCCST_EN_i_0_o3_0_LC_4_12_5  (
            .in0(N__21987),
            .in1(N__35820),
            .in2(N__24100),
            .in3(N__22113),
            .lcout(VCCST_EN_i_0_o3_0),
            .ltout(VCCST_EN_i_0_o3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI6BE8E_1_LC_4_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI6BE8E_1_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI6BE8E_1_LC_4_12_6 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \b2v_inst11.func_state_RNI6BE8E_1_LC_4_12_6  (
            .in0(N__17967),
            .in1(N__17946),
            .in2(N__17926),
            .in3(N__17922),
            .lcout(func_state_RNI6BE8E_0_1),
            .ltout(func_state_RNI6BE8E_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_1_LC_4_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_1_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_1_LC_4_12_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \b2v_inst11.func_state_RNI_1_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17914),
            .in3(N__23349),
            .lcout(\b2v_inst11.N_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIU6GN_7_LC_4_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIU6GN_7_LC_4_13_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \b2v_inst11.count_RNIU6GN_7_LC_4_13_0  (
            .in0(N__24691),
            .in1(N__35827),
            .in2(_gnd_net_),
            .in3(N__17911),
            .lcout(\b2v_inst11.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_7_LC_4_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_7_LC_4_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_7_LC_4_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_7_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24690),
            .lcout(\b2v_inst11.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36603),
            .ce(N__36363),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI18IF_3_LC_4_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI18IF_3_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI18IF_3_LC_4_13_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst11.count_clk_RNI18IF_3_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__18232),
            .in2(N__18114),
            .in3(N__18214),
            .lcout(\b2v_inst11.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI7HLF_6_LC_4_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI7HLF_6_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI7HLF_6_LC_4_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNI7HLF_6_LC_4_13_3  (
            .in0(N__18178),
            .in1(N__18154),
            .in2(_gnd_net_),
            .in3(N__18106),
            .lcout(\b2v_inst11.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIBNNF_8_LC_4_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIBNNF_8_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIBNNF_8_LC_4_13_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \b2v_inst11.count_clk_RNIBNNF_8_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__18148),
            .in2(N__18112),
            .in3(N__18124),
            .lcout(\b2v_inst11.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIV4HF_2_LC_4_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIV4HF_2_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIV4HF_2_LC_4_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIV4HF_2_LC_4_13_5  (
            .in0(N__18391),
            .in1(N__18373),
            .in2(_gnd_net_),
            .in3(N__18102),
            .lcout(\b2v_inst11.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI5EKF_5_LC_4_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI5EKF_5_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI5EKF_5_LC_4_13_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst11.count_clk_RNI5EKF_5_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__18184),
            .in2(N__18113),
            .in3(N__18208),
            .lcout(\b2v_inst11.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIDQOF_9_LC_4_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIDQOF_9_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIDQOF_9_LC_4_13_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_clk_RNIDQOF_9_LC_4_13_7  (
            .in0(N__18283),
            .in1(N__18268),
            .in2(_gnd_net_),
            .in3(N__18095),
            .lcout(\b2v_inst11.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_3_LC_4_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_3_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_3_LC_4_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_3_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18231),
            .lcout(\b2v_inst11.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36611),
            .ce(N__18111),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_5_LC_4_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_5_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_5_LC_4_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_5_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18207),
            .lcout(\b2v_inst11.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36611),
            .ce(N__18111),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_6_LC_4_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_6_LC_4_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_6_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_6_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18177),
            .lcout(\b2v_inst11.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36611),
            .ce(N__18111),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_8_LC_4_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_8_LC_4_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_clk_8_LC_4_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_clk_8_LC_4_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18147),
            .lcout(\b2v_inst11.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36611),
            .ce(N__18111),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_4_15_0 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_0_c_RNO_LC_4_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst20.un4_counter_0_c_RNO_LC_4_15_0  (
            .in0(N__18736),
            .in1(N__18587),
            .in2(N__18450),
            .in3(N__18668),
            .lcout(\b2v_inst20.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_4_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_4_15_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \b2v_inst11.func_state_0_sqmuxa_0_o3_LC_4_15_1  (
            .in0(N__24581),
            .in1(N__24924),
            .in2(N__24520),
            .in3(N__23757),
            .lcout(\b2v_inst11.func_state_0_sqmuxa_0_oZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINPGR_0_1_LC_4_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINPGR_0_1_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINPGR_0_1_LC_4_15_2 .LUT_INIT=16'b0100010011000100;
    LogicCell40 \b2v_inst11.func_state_RNINPGR_0_1_LC_4_15_2  (
            .in0(N__24318),
            .in1(N__23655),
            .in2(N__24056),
            .in3(N__24582),
            .lcout(),
            .ltout(\b2v_inst11.N_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI608H1_1_1_LC_4_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI608H1_1_1_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI608H1_1_1_LC_4_15_3 .LUT_INIT=16'b1111000111110011;
    LogicCell40 \b2v_inst11.func_state_RNI608H1_1_1_LC_4_15_3  (
            .in0(N__24021),
            .in1(N__24317),
            .in2(N__18511),
            .in3(N__26642),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1 ),
            .ltout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNITPOC2_0_LC_4_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNITPOC2_0_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNITPOC2_0_LC_4_15_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst11.func_state_RNITPOC2_0_LC_4_15_4  (
            .in0(N__18699),
            .in1(_gnd_net_),
            .in2(N__18499),
            .in3(N__19839),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_4_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNINPGR_1_LC_4_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNINPGR_1_LC_4_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNINPGR_1_LC_4_15_5 .LUT_INIT=16'b0010101000100010;
    LogicCell40 \b2v_inst11.func_state_RNINPGR_1_LC_4_15_5  (
            .in0(N__23656),
            .in1(N__24319),
            .in2(N__24604),
            .in3(N__24025),
            .lcout(\b2v_inst11.N_381_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_RNIQDE62_LC_4_15_6 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_RNIQDE62_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_RNIQDE62_LC_4_15_6 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \b2v_inst5.RSMRSTn_RNIQDE62_LC_4_15_6  (
            .in0(N__18484),
            .in1(N__21991),
            .in2(N__20287),
            .in3(N__22119),
            .lcout(N_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_3_LC_4_15_7 .C_ON=1'b0;
    defparam \b2v_inst20.counter_3_LC_4_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_3_LC_4_15_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_3_LC_4_15_7  (
            .in0(N__18466),
            .in1(N__18446),
            .in2(_gnd_net_),
            .in3(N__24849),
            .lcout(\b2v_inst20.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36616),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_0_LC_4_16_0 .C_ON=1'b0;
    defparam \b2v_inst20.counter_0_LC_4_16_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_0_LC_4_16_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \b2v_inst20.counter_0_LC_4_16_0  (
            .in0(N__24838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18741),
            .lcout(\b2v_inst20.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36622),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_1_LC_4_16_1 .C_ON=1'b0;
    defparam \b2v_inst20.counter_1_LC_4_16_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_1_LC_4_16_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_1_LC_4_16_1  (
            .in0(N__18740),
            .in1(N__20322),
            .in2(_gnd_net_),
            .in3(N__24841),
            .lcout(\b2v_inst20.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36622),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_4_16_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_4_16_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_0_0_6_LC_4_16_3  (
            .in0(N__24562),
            .in1(N__23991),
            .in2(_gnd_net_),
            .in3(N__24308),
            .lcout(\b2v_inst11.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_4_LC_4_16_4 .C_ON=1'b0;
    defparam \b2v_inst20.counter_4_LC_4_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_4_LC_4_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst20.counter_4_LC_4_16_4  (
            .in0(N__24837),
            .in1(N__18688),
            .in2(_gnd_net_),
            .in3(N__18672),
            .lcout(\b2v_inst20.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36622),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_5_LC_4_16_5 .C_ON=1'b0;
    defparam \b2v_inst20.counter_5_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_5_LC_4_16_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_5_LC_4_16_5  (
            .in0(N__18652),
            .in1(N__20370),
            .in2(_gnd_net_),
            .in3(N__24840),
            .lcout(\b2v_inst20.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36622),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_0_LC_4_16_6 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_0_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_0_LC_4_16_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_0_LC_4_16_6  (
            .in0(N__33688),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(delayed_vccin_vccinaux_ok_RNI8L1J7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_2_LC_4_16_7 .C_ON=1'b0;
    defparam \b2v_inst20.counter_2_LC_4_16_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_2_LC_4_16_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \b2v_inst20.counter_2_LC_4_16_7  (
            .in0(N__18607),
            .in1(N__18591),
            .in2(_gnd_net_),
            .in3(N__24839),
            .lcout(\b2v_inst20.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36622),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_0_0_LC_5_1_0 .C_ON=1'b1;
    defparam \b2v_inst200.count_RNIC03N_0_0_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_0_0_LC_5_1_0 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \b2v_inst200.count_RNIC03N_0_0_LC_5_1_0  (
            .in0(N__22317),
            .in1(N__20622),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_1_0 ),
            .ltout(),
            .carryin(bfn_5_1_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_1_cy ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_5_0_LC_5_1_1 .C_ON=1'b1;
    defparam \b2v_inst200.count_RNIC03N_5_0_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_5_0_LC_5_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.count_RNIC03N_5_0_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__18567),
            .in2(_gnd_net_),
            .in3(N__18547),
            .lcout(\b2v_inst200.count_RNIC03N_5Z0Z_0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_1_cy ),
            .carryout(\b2v_inst200.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_1_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_1_c_RNIJNSD_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(N__18543),
            .in2(_gnd_net_),
            .in3(N__18523),
            .lcout(\b2v_inst200.un2_count_1_cry_1_c_RNIJNSDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_1 ),
            .carryout(\b2v_inst200.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_1_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_2_c_RNIKPTD_LC_5_1_3  (
            .in0(_gnd_net_),
            .in1(N__18852),
            .in2(_gnd_net_),
            .in3(N__18832),
            .lcout(\b2v_inst200.un2_count_1_cry_2_c_RNIKPTDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_2 ),
            .carryout(\b2v_inst200.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_1_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_3_c_RNILRUD_LC_5_1_4  (
            .in0(_gnd_net_),
            .in1(N__18828),
            .in2(_gnd_net_),
            .in3(N__18805),
            .lcout(\b2v_inst200.un2_count_1_cry_3_c_RNILRUDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_3 ),
            .carryout(\b2v_inst200.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_1_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_4_c_RNIMTVD_LC_5_1_5  (
            .in0(_gnd_net_),
            .in1(N__20589),
            .in2(_gnd_net_),
            .in3(N__18784),
            .lcout(\b2v_inst200.un2_count_1_cry_4_c_RNIMTVDZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_4 ),
            .carryout(\b2v_inst200.un2_count_1_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_1_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_5_c_RNINV0E_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(N__20479),
            .in2(_gnd_net_),
            .in3(N__18781),
            .lcout(\b2v_inst200.un2_count_1_cry_5_c_RNINV0EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_5_cZ0 ),
            .carryout(\b2v_inst200.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_1_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_6_c_RNIO12E_LC_5_1_7  (
            .in0(_gnd_net_),
            .in1(N__20610),
            .in2(_gnd_net_),
            .in3(N__18760),
            .lcout(\b2v_inst200.un2_count_1_cry_6_c_RNIO12EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_6 ),
            .carryout(\b2v_inst200.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_7_c_RNIP33E_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__20469),
            .in2(_gnd_net_),
            .in3(N__18757),
            .lcout(\b2v_inst200.un2_count_1_cry_7_c_RNIP33EZ0 ),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_2_1 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_8_c_RNIQ54E_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__25258),
            .in2(_gnd_net_),
            .in3(N__18754),
            .lcout(\b2v_inst200.un2_count_1_cry_8_c_RNIQ54EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_8 ),
            .carryout(\b2v_inst200.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_2_2 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_2_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst200.un2_count_1_cry_9_c_RNIR75E_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20995),
            .in3(N__18751),
            .lcout(\b2v_inst200.un2_count_1_cry_9_c_RNIR75EZ0 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_9 ),
            .carryout(\b2v_inst200.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_2_3 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_10_c_RNI3A29_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__21079),
            .in2(_gnd_net_),
            .in3(N__18907),
            .lcout(\b2v_inst200.un2_count_1_cry_10_c_RNI3AZ0Z29 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_10 ),
            .carryout(\b2v_inst200.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_2_4 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_11_c_RNI4C39_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__20409),
            .in2(_gnd_net_),
            .in3(N__18889),
            .lcout(\b2v_inst200.un2_count_1_cry_11_c_RNI4CZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_11 ),
            .carryout(\b2v_inst200.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_2_5 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_12_c_RNI5E49_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__20632),
            .in2(_gnd_net_),
            .in3(N__18886),
            .lcout(\b2v_inst200.un2_count_1_cry_12_c_RNI5EZ0Z49 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_12 ),
            .carryout(\b2v_inst200.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_2_6 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_13_c_RNI6G59_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__20520),
            .in2(_gnd_net_),
            .in3(N__18883),
            .lcout(\b2v_inst200.un2_count_1_cry_13_c_RNI6GZ0Z59 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_13 ),
            .carryout(\b2v_inst200.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_5_2_7 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_5_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_14_c_RNI7I69_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__20562),
            .in2(_gnd_net_),
            .in3(N__18880),
            .lcout(\b2v_inst200.un2_count_1_cry_14_c_RNI7IZ0Z69 ),
            .ltout(),
            .carryin(\b2v_inst200.un2_count_1_cry_14 ),
            .carryout(\b2v_inst200.un2_count_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_0 .C_ON=1'b1;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst200.un2_count_1_cry_15_c_RNI8K79_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__21057),
            .in2(_gnd_net_),
            .in3(N__18877),
            .lcout(\b2v_inst200.un2_count_1_cry_15_c_RNI8KZ0Z79 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\b2v_inst200.un2_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_3_1 .C_ON=1'b0;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_3_1 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst200.un2_count_1_cry_16_c_RNI9M89_LC_5_3_1  (
            .in0(N__21073),
            .in1(N__22313),
            .in2(_gnd_net_),
            .in3(N__18874),
            .lcout(\b2v_inst200.un2_count_1_cry_16_c_RNI9MZ0Z89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDCT71_17_LC_5_3_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDCT71_17_LC_5_3_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIDCT71_17_LC_5_3_2  (
            .in0(N__18871),
            .in1(N__18864),
            .in2(_gnd_net_),
            .in3(N__25219),
            .lcout(\b2v_inst200.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIKG1A4_LC_5_4_0 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIKG1A4_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_2_c_RNIKG1A4_LC_5_4_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_2_c_RNIKG1A4_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__18990),
            .in2(_gnd_net_),
            .in3(N__19330),
            .lcout(\b2v_inst11.count_off_1_3 ),
            .ltout(\b2v_inst11.count_off_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI6HMCF_3_LC_5_4_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI6HMCF_3_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI6HMCF_3_LC_5_4_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_off_RNI6HMCF_3_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__18981),
            .in2(N__19015),
            .in3(N__19487),
            .lcout(\b2v_inst11.un3_count_off_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI8KNCF_4_LC_5_4_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI8KNCF_4_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI8KNCF_4_LC_5_4_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.count_off_RNI8KNCF_4_LC_5_4_2  (
            .in0(N__19488),
            .in1(N__18969),
            .in2(N__18961),
            .in3(N__19331),
            .lcout(\b2v_inst11.count_offZ0Z_4 ),
            .ltout(\b2v_inst11.count_offZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI6HMCF_0_3_LC_5_4_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI6HMCF_0_3_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI6HMCF_0_3_LC_5_4_3 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \b2v_inst11.count_off_RNI6HMCF_0_3_LC_5_4_3  (
            .in0(N__19000),
            .in1(N__18982),
            .in2(N__18994),
            .in3(N__19490),
            .lcout(\b2v_inst11.un34_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_3_LC_5_4_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_3_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_3_LC_5_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_3_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__18991),
            .in2(_gnd_net_),
            .in3(N__19335),
            .lcout(\b2v_inst11.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36619),
            .ce(N__19525),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_4_LC_5_4_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_4_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_4_LC_5_4_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_4_LC_5_4_5  (
            .in0(N__19333),
            .in1(_gnd_net_),
            .in2(N__18973),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36619),
            .ce(N__19525),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_14_LC_5_4_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_14_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_14_LC_5_4_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_14_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__18942),
            .in2(_gnd_net_),
            .in3(N__19334),
            .lcout(\b2v_inst11.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36619),
            .ce(N__19525),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIACQGF_14_LC_5_4_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIACQGF_14_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIACQGF_14_LC_5_4_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \b2v_inst11.count_off_RNIACQGF_14_LC_5_4_7  (
            .in0(N__19332),
            .in1(N__18952),
            .in2(N__18946),
            .in3(N__19489),
            .lcout(\b2v_inst11.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4ELCF_0_2_LC_5_5_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4ELCF_0_2_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4ELCF_0_2_LC_5_5_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \b2v_inst11.count_off_RNI4ELCF_0_2_LC_5_5_0  (
            .in0(N__19174),
            .in1(N__18921),
            .in2(N__19537),
            .in3(N__19165),
            .lcout(\b2v_inst11.un34_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4ELCF_2_LC_5_5_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4ELCF_2_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4ELCF_2_LC_5_5_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_off_RNI4ELCF_2_LC_5_5_1  (
            .in0(N__18922),
            .in1(N__19173),
            .in2(_gnd_net_),
            .in3(N__19494),
            .lcout(\b2v_inst11.un3_count_off_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_2_LC_5_5_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_2_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_2_LC_5_5_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_2_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__19185),
            .in2(_gnd_net_),
            .in3(N__19338),
            .lcout(\b2v_inst11.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36612),
            .ce(N__19526),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNIANOCF_5_LC_5_5_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNIANOCF_5_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNIANOCF_5_LC_5_5_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \b2v_inst11.count_off_RNIANOCF_5_LC_5_5_4  (
            .in0(N__19495),
            .in1(N__19092),
            .in2(N__19081),
            .in3(N__19336),
            .lcout(\b2v_inst11.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNICQPCF_0_6_LC_5_5_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNICQPCF_0_6_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNICQPCF_0_6_LC_5_5_5 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \b2v_inst11.count_off_RNICQPCF_0_6_LC_5_5_5  (
            .in0(N__19065),
            .in1(N__19563),
            .in2(N__19153),
            .in3(N__19530),
            .lcout(),
            .ltout(\b2v_inst11.un34_clk_100khz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNI4N0JT1_2_LC_5_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNI4N0JT1_2_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNI4N0JT1_2_LC_5_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst11.count_off_RNI4N0JT1_2_LC_5_5_6  (
            .in0(N__19123),
            .in1(N__19117),
            .in2(N__19111),
            .in3(N__19108),
            .lcout(\b2v_inst11.un34_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_5_LC_5_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_5_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_5_LC_5_5_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \b2v_inst11.count_off_5_LC_5_5_7  (
            .in0(N__19337),
            .in1(_gnd_net_),
            .in2(N__19093),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36612),
            .ce(N__19526),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_6_LC_5_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_6_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_6_LC_5_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.count_off_6_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__19579),
            .in2(_gnd_net_),
            .in3(N__19328),
            .lcout(\b2v_inst11.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36605),
            .ce(N__19521),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_9_LC_5_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_9_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_9_LC_5_6_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_9_LC_5_6_1  (
            .in0(N__19327),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19050),
            .lcout(\b2v_inst11.count_offZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36605),
            .ce(N__19521),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIQS7A4_LC_5_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIQS7A4_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_8_c_RNIQS7A4_LC_5_6_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_8_c_RNIQS7A4_LC_5_6_2  (
            .in0(N__19051),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19329),
            .lcout(\b2v_inst11.count_off_1_9 ),
            .ltout(\b2v_inst11.count_off_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_RNII3TCF_9_LC_5_6_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_RNII3TCF_9_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_off_RNII3TCF_9_LC_5_6_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_off_RNII3TCF_9_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__19035),
            .in2(N__19024),
            .in3(N__19520),
            .lcout(\b2v_inst11.un3_count_off_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNINM4A4_LC_5_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNINM4A4_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_5_c_RNINM4A4_LC_5_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_5_c_RNINM4A4_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__19578),
            .in2(_gnd_net_),
            .in3(N__19325),
            .lcout(\b2v_inst11.count_off_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_off_7_LC_5_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_off_7_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_off_7_LC_5_6_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.count_off_7_LC_5_6_5  (
            .in0(N__19326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19362),
            .lcout(\b2v_inst11.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36605),
            .ce(N__19521),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIOO5A4_LC_5_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIOO5A4_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un3_count_off_1_cry_6_c_RNIOO5A4_LC_5_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.un3_count_off_1_cry_6_c_RNIOO5A4_LC_5_6_6  (
            .in0(N__19363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19324),
            .lcout(\b2v_inst11.count_off_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_15_LC_5_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_15_LC_5_6_7  (
            .in0(N__29614),
            .in1(N__29731),
            .in2(_gnd_net_),
            .in3(N__22687),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIDGA72_LC_5_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIDGA72_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIDGA72_LC_5_7_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIDGA72_LC_5_7_0  (
            .in0(N__23452),
            .in1(N__21508),
            .in2(N__23906),
            .in3(N__23721),
            .lcout(\b2v_inst11.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_5_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_12_LC_5_7_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_12_LC_5_7_1  (
            .in0(N__29047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21402),
            .lcout(\b2v_inst11.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_LC_5_7_2 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_LC_5_7_2  (
            .in0(N__26328),
            .in1(N__29533),
            .in2(N__26196),
            .in3(N__26712),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_5_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_14_LC_5_7_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_14_LC_5_7_3  (
            .in0(N__29730),
            .in1(N__26452),
            .in2(N__26750),
            .in3(N__21108),
            .lcout(\b2v_inst11.un2_count_clk_17_0_a2_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_6_LC_5_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_6_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_6_LC_5_7_4 .LUT_INIT=16'b0101011101011111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_6_LC_5_7_4  (
            .in0(N__23380),
            .in1(N__19732),
            .in2(N__21869),
            .in3(N__20698),
            .lcout(\b2v_inst11.g0_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_1_LC_5_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_1_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_1_LC_5_7_6 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_1_LC_5_7_6  (
            .in0(N__21857),
            .in1(N__21271),
            .in2(N__21823),
            .in3(N__26650),
            .lcout(\b2v_inst11.dutycycle_RNI_9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_4_1_LC_5_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_4_1_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_4_1_LC_5_7_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.func_state_RNI_4_1_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(N__21819),
            .in2(_gnd_net_),
            .in3(N__21853),
            .lcout(\b2v_inst11.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI2T5T7_3_LC_5_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI2T5T7_3_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI2T5T7_3_LC_5_8_0 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \b2v_inst11.dutycycle_RNI2T5T7_3_LC_5_8_0  (
            .in0(N__23044),
            .in1(N__23229),
            .in2(N__19588),
            .in3(N__19603),
            .lcout(\b2v_inst11.dutycycle_eena_8 ),
            .ltout(\b2v_inst11.dutycycle_eena_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_3_LC_5_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_3_LC_5_8_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_3_LC_5_8_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \b2v_inst11.dutycycle_3_LC_5_8_1  (
            .in0(N__19624),
            .in1(N__19630),
            .in2(N__19633),
            .in3(N__27721),
            .lcout(\b2v_inst11.dutycycle_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36595),
            .ce(),
            .sr(N__25976));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNIBC872_LC_5_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNIBC872_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNIBC872_LC_5_8_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_c_RNIBC872_LC_5_8_2  (
            .in0(N__23835),
            .in1(N__23709),
            .in2(N__23521),
            .in3(N__21343),
            .lcout(\b2v_inst11.dutycycle_rst_7 ),
            .ltout(\b2v_inst11.dutycycle_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIP1UUA_3_LC_5_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIP1UUA_3_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIP1UUA_3_LC_5_8_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIP1UUA_3_LC_5_8_3  (
            .in0(N__19623),
            .in1(N__27720),
            .in2(N__19615),
            .in3(N__19612),
            .lcout(\b2v_inst11.dutycycleZ0Z_3 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_5_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_3_LC_5_8_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_3_LC_5_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19606),
            .in3(N__23157),
            .lcout(\b2v_inst11.un1_clk_100khz_43_and_i_0_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_2_1_LC_5_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_2_1_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_2_1_LC_5_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_2_1_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(N__23836),
            .in2(_gnd_net_),
            .in3(N__19597),
            .lcout(\b2v_inst11.un1_clk_100khz_43_and_i_0_c ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIVS8U1_12_LC_5_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIVS8U1_12_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIVS8U1_12_LC_5_8_6 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \b2v_inst11.dutycycle_RNIVS8U1_12_LC_5_8_6  (
            .in0(N__23837),
            .in1(N__23483),
            .in2(N__29048),
            .in3(N__23710),
            .lcout(),
            .ltout(\b2v_inst11.N_307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI9R6T4_12_LC_5_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI9R6T4_12_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI9R6T4_12_LC_5_8_7 .LUT_INIT=16'b0000001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI9R6T4_12_LC_5_8_7  (
            .in0(N__27723),
            .in1(N__19699),
            .in2(N__19702),
            .in3(N__23045),
            .lcout(\b2v_inst11.dutycycle_RNI9R6T4Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_2_LC_5_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_2_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_2_LC_5_9_0 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_2_LC_5_9_0  (
            .in0(N__23231),
            .in1(N__25816),
            .in2(N__21301),
            .in3(N__19651),
            .lcout(\b2v_inst11.N_234_N ),
            .ltout(\b2v_inst11.N_234_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI9R6T4_1_LC_5_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI9R6T4_1_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI9R6T4_1_LC_5_9_1 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \b2v_inst11.func_state_RNI9R6T4_1_LC_5_9_1  (
            .in0(N__23047),
            .in1(N__19693),
            .in2(N__19684),
            .in3(N__27719),
            .lcout(\b2v_inst11.func_state_RNI9R6T4Z0Z_1 ),
            .ltout(\b2v_inst11.func_state_RNI9R6T4Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIA3KA7_11_LC_5_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIA3KA7_11_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIA3KA7_11_LC_5_9_2 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \b2v_inst11.dutycycle_RNIA3KA7_11_LC_5_9_2  (
            .in0(N__21457),
            .in1(N__19668),
            .in2(N__19681),
            .in3(N__25817),
            .lcout(\b2v_inst11.dutycycleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_11_LC_5_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_11_LC_5_9_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_11_LC_5_9_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \b2v_inst11.dutycycle_11_LC_5_9_3  (
            .in0(N__25818),
            .in1(N__21456),
            .in2(N__19672),
            .in3(N__19678),
            .lcout(\b2v_inst11.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36586),
            .ce(),
            .sr(N__25948));
    defparam \b2v_inst11.dutycycle_RNI_2_LC_5_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_LC_5_9_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_LC_5_9_4  (
            .in0(N__26637),
            .in1(N__19660),
            .in2(N__21323),
            .in3(N__30279),
            .lcout(\b2v_inst11.un1_clk_100khz_42_and_i_o2_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_14_LC_5_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_14_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_14_LC_5_9_5 .LUT_INIT=16'b1100000011010101;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_14_LC_5_9_5  (
            .in0(N__25815),
            .in1(N__23230),
            .in2(N__29737),
            .in3(N__26636),
            .lcout(),
            .ltout(\b2v_inst11.N_155_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIMBHI8_14_LC_5_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_14_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_14_LC_5_9_6 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIMBHI8_14_LC_5_9_6  (
            .in0(N__27718),
            .in1(N__23132),
            .in2(N__19645),
            .in3(N__23046),
            .lcout(\b2v_inst11.dutycycle_en_11 ),
            .ltout(\b2v_inst11.dutycycle_en_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_14_LC_5_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_14_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_14_LC_5_9_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \b2v_inst11.dutycycle_14_LC_5_9_7  (
            .in0(N__25819),
            .in1(N__22710),
            .in2(N__19642),
            .in3(N__22741),
            .lcout(\b2v_inst11.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36586),
            .ce(),
            .sr(N__25948));
    defparam \b2v_inst11.func_state_RNIVS8U1_3_1_LC_5_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_3_1_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_3_1_LC_5_10_0 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_3_1_LC_5_10_0  (
            .in0(N__22031),
            .in1(N__20288),
            .in2(N__19858),
            .in3(N__22115),
            .lcout(func_state_RNIVS8U1_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI70K8_0_LC_5_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI70K8_0_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI70K8_0_LC_5_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.func_state_RNI70K8_0_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__24331),
            .in2(_gnd_net_),
            .in3(N__19762),
            .lcout(\b2v_inst11.N_305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIEIB72_LC_5_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIEIB72_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIEIB72_LC_5_10_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIEIB72_LC_5_10_2  (
            .in0(N__23715),
            .in1(N__21496),
            .in2(N__23520),
            .in3(N__23874),
            .lcout(\b2v_inst11.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_3_1_LC_5_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_3_1_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_3_1_LC_5_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.func_state_RNI_3_1_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21813),
            .lcout(\b2v_inst11.N_3060_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_LC_5_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_LC_5_10_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_LC_5_10_4  (
            .in0(N__21379),
            .in1(N__29344),
            .in2(_gnd_net_),
            .in3(N__26102),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_6 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_6_LC_5_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_6_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_6_LC_5_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_6_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19708),
            .in3(N__20699),
            .lcout(\b2v_inst11.N_426_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_5_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_3_LC_5_10_6 .LUT_INIT=16'b0000111001110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_3_LC_5_10_6  (
            .in0(N__28772),
            .in1(N__26337),
            .in2(N__26844),
            .in3(N__29482),
            .lcout(),
            .ltout(\b2v_inst11.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_9_LC_5_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_9_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_9_LC_5_10_7 .LUT_INIT=16'b1101101101000010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_9_LC_5_10_7  (
            .in0(N__26103),
            .in1(N__26448),
            .in2(N__19705),
            .in3(N__26830),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_5_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_5_11_0 .LUT_INIT=16'b0101011111011111;
    LogicCell40 \b2v_inst11.SYNTHESIZED_WIRE_2_i_0_o3_2_LC_5_11_0  (
            .in0(N__24328),
            .in1(N__20277),
            .in2(N__21986),
            .in3(N__22093),
            .lcout(N_15_i_0_a4_1_N_3L3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_5_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_5_11_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst11.dutycycle_1_0_iv_i_a2_6_LC_5_11_1  (
            .in0(N__24587),
            .in1(N__24934),
            .in2(N__24513),
            .in3(N__23853),
            .lcout(\b2v_inst11.N_382 ),
            .ltout(\b2v_inst11.N_382_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQ6_LC_5_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQ6_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQ6_LC_5_11_2 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQ6_LC_5_11_2  (
            .in0(N__23057),
            .in1(N__19912),
            .in2(N__19906),
            .in3(N__27078),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIQHGQZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNIF6NL_0_6_LC_5_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNIF6NL_0_6_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNIF6NL_0_6_LC_5_11_3 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \b2v_inst11.count_clk_RNIF6NL_0_6_LC_5_11_3  (
            .in0(N__23509),
            .in1(N__26649),
            .in2(N__20041),
            .in3(N__20706),
            .lcout(),
            .ltout(\b2v_inst11.g0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_clk_RNI5FOR1_6_LC_5_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_clk_RNI5FOR1_6_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_clk_RNI5FOR1_6_LC_5_11_4 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \b2v_inst11.count_clk_RNI5FOR1_6_LC_5_11_4  (
            .in0(N__21978),
            .in1(N__35896),
            .in2(N__19903),
            .in3(N__22095),
            .lcout(\b2v_inst11.un1_count_off_1_sqmuxa_8_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIRF2E4_0_LC_5_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIRF2E4_0_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIRF2E4_0_LC_5_11_5 .LUT_INIT=16'b0110111100001111;
    LogicCell40 \b2v_inst11.func_state_RNIRF2E4_0_LC_5_11_5  (
            .in0(N__24113),
            .in1(N__24330),
            .in2(N__19900),
            .in3(N__19756),
            .lcout(\b2v_inst11.func_state_RNIRF2E4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_6 .LUT_INIT=16'b1100100000001000;
    LogicCell40 \b2v_inst11.VCCST_EN_i_0_i_LC_5_11_6  (
            .in0(N__21977),
            .in1(N__24111),
            .in2(N__35929),
            .in3(N__22094),
            .lcout(VCCST_EN_i_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIF6NL_1_LC_5_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIF6NL_1_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIF6NL_1_LC_5_11_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \b2v_inst11.func_state_RNIF6NL_1_LC_5_11_7  (
            .in0(N__24112),
            .in1(N__24329),
            .in2(_gnd_net_),
            .in3(N__23587),
            .lcout(\b2v_inst11.un1_clk_100khz_2_i_o3_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIVS8U1_0_LC_5_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIVS8U1_0_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIVS8U1_0_LC_5_12_0 .LUT_INIT=16'b1110111011111100;
    LogicCell40 \b2v_inst11.func_state_RNIVS8U1_0_LC_5_12_0  (
            .in0(N__19813),
            .in1(N__26915),
            .in2(N__33617),
            .in3(N__23617),
            .lcout(\b2v_inst11.dutycycle_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI98672_LC_5_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI98672_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI98672_LC_5_12_1 .LUT_INIT=16'b1111101111110001;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_RNI98672_LC_5_12_1  (
            .in0(N__23618),
            .in1(N__21361),
            .in2(N__26931),
            .in3(N__19814),
            .lcout(\b2v_inst11.dutycycle_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI_0_0_LC_5_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI_0_0_LC_5_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst11.func_state_RNI_0_0_LC_5_12_2  (
            .in0(N__19815),
            .in1(N__20707),
            .in2(_gnd_net_),
            .in3(N__20021),
            .lcout(\b2v_inst11.func_state_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_0_LC_5_12_3 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_0_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_0_LC_5_12_3 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \b2v_inst5.curr_state_0_LC_5_12_3  (
            .in0(N__21944),
            .in1(N__25548),
            .in2(_gnd_net_),
            .in3(N__22096),
            .lcout(\b2v_inst5.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36604),
            .ce(N__36364),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI_0_LC_5_12_4 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI_0_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI_0_LC_5_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst5.curr_state_RNI_0_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21924),
            .lcout(\b2v_inst5.N_2897_i ),
            .ltout(\b2v_inst5.N_2897_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_5_12_5 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_LC_5_12_5 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(N__22098),
            .in2(N__19930),
            .in3(N__25547),
            .lcout(),
            .ltout(\b2v_inst5.m4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI1CVE1_0_LC_5_12_6 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI1CVE1_0_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI1CVE1_0_LC_5_12_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.curr_state_RNI1CVE1_0_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__19927),
            .in2(N__19921),
            .in3(N__35819),
            .lcout(\b2v_inst5.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.g0_8_LC_5_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.g0_8_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.g0_8_LC_5_12_7 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \b2v_inst11.g0_8_LC_5_12_7  (
            .in0(N__23510),
            .in1(N__21979),
            .in2(N__24932),
            .in3(N__22097),
            .lcout(\b2v_inst11.N_165_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_1_LC_5_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_1_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_1_LC_5_13_0 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_1_LC_5_13_0  (
            .in0(N__21420),
            .in1(N__21324),
            .in2(_gnd_net_),
            .in3(N__33321),
            .lcout(),
            .ltout(\b2v_inst11.g2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_12_LC_5_13_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_12_LC_5_13_1  (
            .in0(N__29049),
            .in1(N__33595),
            .in2(N__19918),
            .in3(N__26190),
            .lcout(\b2v_inst11.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNISSAOS1_5_LC_5_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNISSAOS1_5_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNISSAOS1_5_LC_5_13_2 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \b2v_inst11.dutycycle_RNISSAOS1_5_LC_5_13_2  (
            .in0(N__20146),
            .in1(N__20158),
            .in2(N__20167),
            .in3(N__27534),
            .lcout(dutycycle_RNISSAOS1_0_5),
            .ltout(dutycycle_RNISSAOS1_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_LC_5_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_LC_5_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19915),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_5 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_1_LC_5_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_1_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_1_LC_5_13_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_1_LC_5_13_4  (
            .in0(N__26192),
            .in1(N__33597),
            .in2(N__20044),
            .in3(N__33322),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.N_224_i_LC_5_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.N_224_i_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.N_224_i_LC_5_13_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.N_224_i_LC_5_13_5  (
            .in0(N__24484),
            .in1(N__35826),
            .in2(N__23905),
            .in3(N__24586),
            .lcout(\b2v_inst11.N_224_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_1_LC_5_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_1_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_1_LC_5_13_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_1_LC_5_13_6  (
            .in0(N__21421),
            .in1(N__29050),
            .in2(N__33353),
            .in3(N__21325),
            .lcout(),
            .ltout(\b2v_inst11.N_73_mux_i_i_o7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_LC_5_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_LC_5_13_7 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_LC_5_13_7  (
            .in0(N__33596),
            .in1(N__26635),
            .in2(N__20008),
            .in3(N__26191),
            .lcout(N_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI52GVC_5_LC_5_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI52GVC_5_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI52GVC_5_LC_5_14_0 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \b2v_inst11.dutycycle_RNI52GVC_5_LC_5_14_0  (
            .in0(N__20124),
            .in1(N__27688),
            .in2(N__27285),
            .in3(N__20005),
            .lcout(\b2v_inst11.N_73_mux_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIUNGA5_5_LC_5_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIUNGA5_5_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIUNGA5_5_LC_5_14_1 .LUT_INIT=16'b1011101100011011;
    LogicCell40 \b2v_inst11.dutycycle_RNIUNGA5_5_LC_5_14_1  (
            .in0(N__27687),
            .in1(N__20123),
            .in2(N__23058),
            .in3(N__20083),
            .lcout(\b2v_inst11.dutycycle_RNIUNGA5Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI4NJR6_5_LC_5_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI4NJR6_5_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI4NJR6_5_LC_5_14_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI4NJR6_5_LC_5_14_2  (
            .in0(N__20125),
            .in1(N__19990),
            .in2(N__20101),
            .in3(N__19965),
            .lcout(),
            .ltout(\b2v_inst11.N_73_mux_i_i_a7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI7JLNN_5_LC_5_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI7JLNN_5_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI7JLNN_5_LC_5_14_3 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI7JLNN_5_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__19999),
            .in2(N__19993),
            .in3(N__26053),
            .lcout(\b2v_inst11.N_73_mux_i_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_5_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_0_LC_5_14_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_0_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__19989),
            .in2(_gnd_net_),
            .in3(N__19966),
            .lcout(),
            .ltout(N_73_mux_i_i_a7_4_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_fast_RNIVS8U1_0_LC_5_14_5 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_RNIVS8U1_0_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_fast_RNIVS8U1_0_LC_5_14_5 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_RNIVS8U1_0_LC_5_14_5  (
            .in0(N__19951),
            .in1(N__23792),
            .in2(N__19933),
            .in3(N__29329),
            .lcout(),
            .ltout(N_73_mux_i_i_a7_4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI74U7G_5_LC_5_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI74U7G_5_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI74U7G_5_LC_5_14_6 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI74U7G_5_LC_5_14_6  (
            .in0(N__20122),
            .in1(N__27552),
            .in2(N__20170),
            .in3(N__20094),
            .lcout(\b2v_inst11.N_73_mux_i_i_1 ),
            .ltout(\b2v_inst11.N_73_mux_i_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_5_LC_5_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_5_LC_5_14_7 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_5_LC_5_14_7 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \b2v_inst11.dutycycle_5_LC_5_14_7  (
            .in0(N__20157),
            .in1(N__20145),
            .in2(N__20128),
            .in3(N__27535),
            .lcout(\b2v_inst11.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36618),
            .ce(),
            .sr(N__25937));
    defparam \b2v_inst11.func_state_RNIDGAL3_0_0_LC_5_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIDGAL3_0_0_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIDGAL3_0_0_LC_5_15_0 .LUT_INIT=16'b1111111101000111;
    LogicCell40 \b2v_inst11.func_state_RNIDGAL3_0_0_LC_5_15_0  (
            .in0(N__22066),
            .in1(N__20259),
            .in2(N__22021),
            .in3(N__20110),
            .lcout(\b2v_inst11.N_140_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_fast_RNIGMH81_LC_5_15_1 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_RNIGMH81_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_fast_RNIGMH81_LC_5_15_1 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_RNIGMH81_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__22009),
            .in2(N__20276),
            .in3(N__22065),
            .lcout(RSMRSTn_fast_RNIGMH81),
            .ltout(RSMRSTn_fast_RNIGMH81_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_rep1_RNIABFM6_LC_5_15_2 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_rep1_RNIABFM6_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.tmp_1_rep1_RNIABFM6_LC_5_15_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst20.tmp_1_rep1_RNIABFM6_LC_5_15_2  (
            .in0(N__20065),
            .in1(_gnd_net_),
            .in2(N__20104),
            .in3(N__20082),
            .lcout(N_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_LC_5_15_3 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_LC_5_15_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst20.tmp_1_LC_5_15_3  (
            .in0(N__24857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35887),
            .lcout(SYNTHESIZED_WIRE_1keep_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36624),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_rep1_RNI07F73_LC_5_15_4 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_rep1_RNI07F73_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.tmp_1_rep1_RNI07F73_LC_5_15_4 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \b2v_inst20.tmp_1_rep1_RNI07F73_LC_5_15_4  (
            .in0(N__24510),
            .in1(N__24580),
            .in2(N__24933),
            .in3(N__20081),
            .lcout(\b2v_inst20.tmp_1_rep1_RNI07FZ0Z73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.counter_6_LC_5_15_5 .C_ON=1'b0;
    defparam \b2v_inst20.counter_6_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.counter_6_LC_5_15_5 .LUT_INIT=16'b0000011000000110;
    LogicCell40 \b2v_inst20.counter_6_LC_5_15_5  (
            .in0(N__20059),
            .in1(N__20342),
            .in2(N__24864),
            .in3(_gnd_net_),
            .lcout(\b2v_inst20.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36624),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_5_15_6 .C_ON=1'b0;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst20.un4_counter_1_c_RNO_LC_5_15_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst20.un4_counter_1_c_RNO_LC_5_15_6  (
            .in0(N__20392),
            .in1(N__20366),
            .in2(N__20346),
            .in3(N__20318),
            .lcout(\b2v_inst20.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_fast_LC_5_15_7 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_fast_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_fast_LC_5_15_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst20.tmp_1_fast_LC_5_15_7  (
            .in0(N__20260),
            .in1(_gnd_net_),
            .in2(N__24865),
            .in3(_gnd_net_),
            .lcout(SYNTHESIZED_WIRE_1keep_3_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36624),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_ATP_RNIQFGQ_LC_5_16_0 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_ATP_RNIQFGQ_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.HDA_SDO_ATP_RNIQFGQ_LC_5_16_0 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \b2v_inst200.HDA_SDO_ATP_RNIQFGQ_LC_5_16_0  (
            .in0(N__35815),
            .in1(N__20215),
            .in2(N__20191),
            .in3(N__20203),
            .lcout(HDA_SDO_ATP_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_16_1 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI_0_LC_5_16_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst200.curr_state_RNI_0_LC_5_16_1  (
            .in0(N__22186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22229),
            .lcout(\b2v_inst200.N_205 ),
            .ltout(\b2v_inst200.N_205_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_16_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_16_2 .LUT_INIT=16'b1011101010111011;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_LC_5_16_2  (
            .in0(N__22595),
            .in1(N__20202),
            .in2(N__20209),
            .in3(N__33686),
            .lcout(G_2734),
            .ltout(G_2734_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNI52VB_2_LC_5_16_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNI52VB_2_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNI52VB_2_LC_5_16_3 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \b2v_inst200.curr_state_RNI52VB_2_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__20176),
            .in2(N__20206),
            .in3(N__35814),
            .lcout(\b2v_inst200.curr_stateZ0Z_2 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_16_4 .C_ON=1'b0;
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.HDA_SDO_ATP_LC_5_16_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \b2v_inst200.HDA_SDO_ATP_LC_5_16_4  (
            .in0(N__22230),
            .in1(_gnd_net_),
            .in2(N__20194),
            .in3(N__22190),
            .lcout(\b2v_inst200.HDA_SDO_ATP_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36628),
            .ce(N__36357),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_2_LC_5_16_6 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_2_LC_5_16_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_2_LC_5_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst200.curr_state_2_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20182),
            .lcout(\b2v_inst200.curr_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36628),
            .ce(N__36357),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_0_LC_5_16_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_0_LC_5_16_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_0_LC_5_16_7 .LUT_INIT=16'b1101110011001101;
    LogicCell40 \b2v_inst200.curr_state_0_LC_5_16_7  (
            .in0(N__33687),
            .in1(N__22249),
            .in2(N__22195),
            .in3(N__22231),
            .lcout(\b2v_inst200.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36628),
            .ce(N__36357),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIDC651_8_LC_6_1_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIDC651_8_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIDC651_8_LC_6_1_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst200.count_RNIDC651_8_LC_6_1_0  (
            .in0(N__25205),
            .in1(N__20431),
            .in2(N__22329),
            .in3(N__20439),
            .lcout(\b2v_inst200.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI96451_6_LC_6_1_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI96451_6_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI96451_6_LC_6_1_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst200.count_RNI96451_6_LC_6_1_1  (
            .in0(N__20457),
            .in1(N__22318),
            .in2(N__20449),
            .in3(N__25204),
            .lcout(\b2v_inst200.countZ0Z_6 ),
            .ltout(\b2v_inst200.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_6_LC_6_1_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_6_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_6_LC_6_1_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \b2v_inst200.count_RNI_6_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20473),
            .in3(N__20470),
            .lcout(\b2v_inst200.un25_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_6_LC_6_1_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_6_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_6_LC_6_1_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst200.count_6_LC_6_1_3  (
            .in0(N__20458),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22324),
            .lcout(\b2v_inst200.count_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36642),
            .ce(N__25158),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_8_LC_6_1_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_8_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_8_LC_6_1_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst200.count_8_LC_6_1_4  (
            .in0(N__22325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20440),
            .lcout(\b2v_inst200.count_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36642),
            .ce(N__25158),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_0_LC_6_1_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_0_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_0_LC_6_1_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst200.count_RNIC03N_0_LC_6_1_5  (
            .in0(N__20416),
            .in1(N__20425),
            .in2(_gnd_net_),
            .in3(N__25203),
            .lcout(\b2v_inst200.countZ0Z_0 ),
            .ltout(\b2v_inst200.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_0_LC_6_1_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_0_LC_6_1_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_0_LC_6_1_6 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \b2v_inst200.count_0_LC_6_1_6  (
            .in0(N__22322),
            .in1(_gnd_net_),
            .in2(N__20419),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36642),
            .ce(N__25158),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_16_LC_6_1_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_16_LC_6_1_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_16_LC_6_1_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_16_LC_6_1_7  (
            .in0(_gnd_net_),
            .in1(N__22323),
            .in2(_gnd_net_),
            .in3(N__20497),
            .lcout(\b2v_inst200.count_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36642),
            .ce(N__25158),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_9_LC_6_2_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_9_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_9_LC_6_2_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst200.count_RNI_9_LC_6_2_0  (
            .in0(_gnd_net_),
            .in1(N__25257),
            .in2(_gnd_net_),
            .in3(N__20410),
            .lcout(\b2v_inst200.un25_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI50P71_13_LC_6_2_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI50P71_13_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI50P71_13_LC_6_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst200.count_RNI50P71_13_LC_6_2_1  (
            .in0(N__20653),
            .in1(N__25216),
            .in2(_gnd_net_),
            .in3(N__20643),
            .lcout(\b2v_inst200.countZ0Z_13 ),
            .ltout(\b2v_inst200.countZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_1_0_LC_6_2_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_1_0_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_1_0_LC_6_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst200.count_RNIC03N_1_0_LC_6_2_2  (
            .in0(N__20521),
            .in1(N__20563),
            .in2(N__20626),
            .in3(N__20623),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_3_0_LC_6_2_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_3_0_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_3_0_LC_6_2_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst200.count_RNIC03N_3_0_LC_6_2_3  (
            .in0(N__20611),
            .in1(N__20590),
            .in2(N__20572),
            .in3(N__20569),
            .lcout(\b2v_inst200.un25_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_14_LC_6_2_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_14_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_14_LC_6_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_14_LC_6_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20536),
            .lcout(\b2v_inst200.count_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36636),
            .ce(N__25156),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI96R71_15_LC_6_2_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI96R71_15_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI96R71_15_LC_6_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI96R71_15_LC_6_2_5  (
            .in0(N__20550),
            .in1(N__20542),
            .in2(_gnd_net_),
            .in3(N__25218),
            .lcout(\b2v_inst200.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_15_LC_6_2_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_15_LC_6_2_6 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_15_LC_6_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_15_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20551),
            .lcout(\b2v_inst200.count_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36636),
            .ce(N__25156),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI73Q71_14_LC_6_2_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI73Q71_14_LC_6_2_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNI73Q71_14_LC_6_2_7  (
            .in0(N__20535),
            .in1(N__20527),
            .in2(_gnd_net_),
            .in3(N__25217),
            .lcout(\b2v_inst200.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIB9S71_16_LC_6_3_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIB9S71_16_LC_6_3_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \b2v_inst200.count_RNIB9S71_16_LC_6_3_0  (
            .in0(N__25215),
            .in1(N__20509),
            .in2(N__20496),
            .in3(N__22310),
            .lcout(\b2v_inst200.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_11_LC_6_3_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_11_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_11_LC_6_3_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst200.count_11_LC_6_3_1  (
            .in0(N__22312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21097),
            .lcout(\b2v_inst200.count_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36630),
            .ce(N__25155),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_10_LC_6_3_2 .C_ON=1'b0;
    defparam \b2v_inst200.count_10_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_10_LC_6_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.count_10_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__21012),
            .in2(_gnd_net_),
            .in3(N__22311),
            .lcout(\b2v_inst200.count_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36630),
            .ce(N__25155),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI1QM71_11_LC_6_3_3 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI1QM71_11_LC_6_3_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \b2v_inst200.count_RNI1QM71_11_LC_6_3_3  (
            .in0(N__22309),
            .in1(N__21096),
            .in2(N__21088),
            .in3(N__25214),
            .lcout(\b2v_inst200.countZ0Z_11 ),
            .ltout(\b2v_inst200.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_17_LC_6_3_4 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_17_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_17_LC_6_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNI_17_LC_6_3_4  (
            .in0(N__20994),
            .in1(N__21072),
            .in2(N__21061),
            .in3(N__21058),
            .lcout(),
            .ltout(\b2v_inst200.un25_clk_100khz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIC03N_6_0_LC_6_3_5 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIC03N_6_0_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIC03N_6_0_LC_6_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst200.count_RNIC03N_6_0_LC_6_3_5  (
            .in0(N__21046),
            .in1(N__21037),
            .in2(N__21025),
            .in3(N__21022),
            .lcout(\b2v_inst200.count_RNIC03N_6Z0Z_0 ),
            .ltout(\b2v_inst200.count_RNIC03N_6Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNI_0_LC_6_3_6 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNI_0_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNI_0_LC_6_3_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst200.count_RNI_0_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21016),
            .in3(_gnd_net_),
            .lcout(\b2v_inst200.count_RNI_0_0 ),
            .ltout(\b2v_inst200.count_RNI_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_6_3_7 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIOMPC1_10_LC_6_3_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \b2v_inst200.count_RNIOMPC1_10_LC_6_3_7  (
            .in0(N__21013),
            .in1(N__21004),
            .in2(N__20998),
            .in3(N__25213),
            .lcout(\b2v_inst200.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.count_12_LC_6_4_0 .C_ON=1'b0;
    defparam \b2v_inst16.count_12_LC_6_4_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst16.count_12_LC_6_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst16.count_12_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20980),
            .lcout(\b2v_inst16.count_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36626),
            .ce(N__20950),
            .sr(N__20800));
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_6_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_2_LC_6_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_2_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__30287),
            .in2(_gnd_net_),
            .in3(N__21280),
            .lcout(\b2v_inst11.N_366 ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__25444),
            .in2(N__21242),
            .in3(N__21262),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_2_c ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__28249),
            .in2(N__21244),
            .in3(N__21259),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_3_c ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__28231),
            .in2(N__32519),
            .in3(N__21256),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_4_c ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__28210),
            .in2(N__32520),
            .in3(N__21253),
            .lcout(\b2v_inst11.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_5_c ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_6_6_5  (
            .in0(N__31706),
            .in1(N__28192),
            .in2(N__21243),
            .in3(N__21250),
            .lcout(\b2v_inst11.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un152_sum_cry_6_c ),
            .carryout(\b2v_inst11.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__28408),
            .in2(_gnd_net_),
            .in3(N__21247),
            .lcout(\b2v_inst11.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_6_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_6_6_7  (
            .in0(N__32509),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_6_7_0 .C_ON=1'b0;
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_6_7_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \b2v_inst16.curr_state_1_sqmuxa_1_i_o3_0_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__21220),
            .in2(_gnd_net_),
            .in3(N__21200),
            .lcout(\b2v_inst16.N_208_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_LC_6_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_LC_6_7_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_LC_6_7_1  (
            .in0(N__26777),
            .in1(N__21378),
            .in2(N__21118),
            .in3(N__26647),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_6_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_10_LC_6_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_10_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__26326),
            .in2(_gnd_net_),
            .in3(N__29216),
            .lcout(),
            .ltout(\b2v_inst11.un2_count_clk_17_0_a2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_6_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_15_LC_6_7_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_15_LC_6_7_3  (
            .in0(N__28895),
            .in1(N__21334),
            .in2(N__21328),
            .in3(N__29612),
            .lcout(\b2v_inst11.N_363 ),
            .ltout(\b2v_inst11.N_363_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_6_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_15_LC_6_7_4 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_15_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__21297),
            .in2(N__21283),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_365 ),
            .ltout(\b2v_inst11.N_365_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_1_LC_6_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_6_1_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_1_LC_6_7_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_1_LC_6_7_5  (
            .in0(N__33613),
            .in1(N__26179),
            .in2(N__21274),
            .in3(N__33352),
            .lcout(\b2v_inst11.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_7_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \b2v_inst11.un1_count_clk_1_sqmuxa_0_o3_0_LC_6_7_6  (
            .in0(N__24365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24155),
            .lcout(N_161),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_6_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_6_LC_6_7_7 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_6_LC_6_7_7  (
            .in0(N__26776),
            .in1(N__29534),
            .in2(_gnd_net_),
            .in3(N__26178),
            .lcout(\b2v_inst11.g0_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_6_8_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_11_LC_6_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_11_LC_6_8_0  (
            .in0(N__29102),
            .in1(N__26301),
            .in2(N__21439),
            .in3(N__26800),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_6_8_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_8_LC_6_8_1 .LUT_INIT=16'b0101011101011111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_8_LC_6_8_1  (
            .in0(N__26299),
            .in1(N__29498),
            .in2(N__26832),
            .in3(N__26183),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_6_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_3_LC_6_8_2 .LUT_INIT=16'b1111100011100000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_3_LC_6_8_2  (
            .in0(N__28755),
            .in1(N__26798),
            .in2(N__29532),
            .in3(N__26300),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_6_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_8_3_LC_6_8_3 .LUT_INIT=16'b0001001100110111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_8_3_LC_6_8_3  (
            .in0(N__26445),
            .in1(N__29499),
            .in2(N__26327),
            .in3(N__28754),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_30_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_6_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_9_LC_6_8_4 .LUT_INIT=16'b1010111010001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_9_LC_6_8_4  (
            .in0(N__26184),
            .in1(N__26799),
            .in2(N__21442),
            .in3(N__26446),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_6_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_13_LC_6_8_5 .LUT_INIT=16'b0111010111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_13_LC_6_8_5  (
            .in0(N__28896),
            .in1(N__29198),
            .in2(N__21413),
            .in3(N__29037),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_6_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_9_LC_6_8_6 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_9_LC_6_8_6  (
            .in0(N__21430),
            .in1(N__26447),
            .in2(N__21424),
            .in3(N__21406),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_6_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_11_LC_6_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_11_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29101),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_7_1_LC_6_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_7_1_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_7_1_LC_6_9_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_7_1_LC_6_9_0  (
            .in0(N__33360),
            .in1(N__33621),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.dutycycle_RNI_7Z0Z_1 ),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABT8_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__33359),
            .in2(N__27132),
            .in3(N__21349),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_0_c_RNIABTZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI_LC_6_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI_LC_6_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNI_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__27108),
            .in2(N__30278),
            .in3(N__21346),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_1_c_RNIZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFV8_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__27059),
            .in2(N__28757),
            .in3(N__21337),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_2_c_RNICFVZ0Z8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_2 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDH09_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__29509),
            .in2(N__27104),
            .in3(N__21511),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_3_c_RNIDHZ0Z09 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_3 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_6_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_6_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJ19_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__27054),
            .in2(N__29389),
            .in3(N__21499),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_4_c_RNIEJZ0Z19 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_4_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_6_9_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_6_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFL29_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(N__26157),
            .in2(N__27103),
            .in3(N__21484),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_5_c_RNIFLZ0Z29 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_9_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGN39_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__27058),
            .in2(N__26842),
            .in3(N__21469),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_6_c_RNIGNZ0Z39 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHP49_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__27088),
            .in2(N__26336),
            .in3(N__21466),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_7_c_RNIHPZ0Z49 ),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIR59_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__26438),
            .in2(N__27129),
            .in3(N__21463),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_8_c_RNIIRZ0Z59 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_8_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJT69_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(N__27092),
            .in2(N__29215),
            .in3(N__21460),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_9_c_RNIJTZ0Z69 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_9 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNP5_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__29115),
            .in2(N__27130),
            .in3(N__21448),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_10_c_RNIRNPZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_10_cZ0 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQ5_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__27096),
            .in2(N__29046),
            .in3(N__21445),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_11_c_RNISPQZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_11 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRR5_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__28899),
            .in2(N__27131),
            .in3(N__21574),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_12_c_RNITRRZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_12 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_10_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTS5_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__27100),
            .in2(N__29725),
            .in3(N__21571),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_13_c_RNIUTSZ0Z5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_94_cry_13 ),
            .carryout(\b2v_inst11.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVT5_LC_6_10_7  (
            .in0(N__27101),
            .in1(N__29608),
            .in2(_gnd_net_),
            .in3(N__21568),
            .lcout(\b2v_inst11.un1_dutycycle_94_cry_14_c_RNIVVTZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_4_LC_6_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_4_LC_6_11_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_4_LC_6_11_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \b2v_inst11.dutycycle_4_LC_6_11_0  (
            .in0(N__21556),
            .in1(N__23053),
            .in2(N__21550),
            .in3(N__21523),
            .lcout(\b2v_inst11.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36606),
            .ce(),
            .sr(N__25972));
    defparam \b2v_inst11.dutycycle_RNIP7P13_4_LC_6_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIP7P13_4_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIP7P13_4_LC_6_11_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \b2v_inst11.dutycycle_RNIP7P13_4_LC_6_11_1  (
            .in0(N__27710),
            .in1(N__25811),
            .in2(N__21549),
            .in3(N__21565),
            .lcout(\b2v_inst11.dutycycle_RNIP7P13Z0Z_4 ),
            .ltout(\b2v_inst11.dutycycle_RNIP7P13Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIKF34B_4_LC_6_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIKF34B_4_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIKF34B_4_LC_6_11_2 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \b2v_inst11.dutycycle_RNIKF34B_4_LC_6_11_2  (
            .in0(N__21545),
            .in1(N__23051),
            .in2(N__21529),
            .in3(N__21522),
            .lcout(\b2v_inst11.dutycycleZ0Z_7 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_4_LC_6_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_4_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_4_LC_6_11_3 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_4_LC_6_11_3  (
            .in0(N__23167),
            .in1(N__23259),
            .in2(N__21526),
            .in3(N__23232),
            .lcout(\b2v_inst11.dutycycle_e_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_15_LC_6_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_15_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_15_LC_6_11_4 .LUT_INIT=16'b1010101100000011;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_15_LC_6_11_4  (
            .in0(N__23233),
            .in1(N__26648),
            .in2(N__25853),
            .in3(N__29613),
            .lcout(),
            .ltout(\b2v_inst11.N_158_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIMBHI8_15_LC_6_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_15_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_15_LC_6_11_5 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIMBHI8_15_LC_6_11_5  (
            .in0(N__23052),
            .in1(N__23175),
            .in2(N__21514),
            .in3(N__27664),
            .lcout(\b2v_inst11.dutycycle_en_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_6_LC_6_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_6_LC_6_11_6 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_6_LC_6_11_6 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \b2v_inst11.dutycycle_6_LC_6_11_6  (
            .in0(N__21691),
            .in1(N__21699),
            .in2(N__27700),
            .in3(N__21712),
            .lcout(\b2v_inst11.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36606),
            .ce(),
            .sr(N__25972));
    defparam \b2v_inst11.dutycycle_RNIQGT7G_6_LC_6_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIQGT7G_6_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIQGT7G_6_LC_6_11_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIQGT7G_6_LC_6_11_7  (
            .in0(N__21711),
            .in1(N__27663),
            .in2(N__21703),
            .in3(N__21690),
            .lcout(\b2v_inst11.dutycycleZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNIMJCJ5_1_LC_6_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNIMJCJ5_1_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNIMJCJ5_1_LC_6_12_0 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \b2v_inst11.func_state_RNIMJCJ5_1_LC_6_12_0  (
            .in0(_gnd_net_),
            .in1(N__24637),
            .in2(N__33754),
            .in3(N__21790),
            .lcout(),
            .ltout(\b2v_inst11.N_186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8E1K7_1_LC_6_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8E1K7_1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8E1K7_1_LC_6_12_1 .LUT_INIT=16'b0000111110111111;
    LogicCell40 \b2v_inst11.func_state_RNI8E1K7_1_LC_6_12_1  (
            .in0(N__21676),
            .in1(N__24125),
            .in2(N__21646),
            .in3(N__33729),
            .lcout(\b2v_inst11.N_117_f0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIVS8U1_6_LC_6_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIVS8U1_6_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIVS8U1_6_LC_6_12_2 .LUT_INIT=16'b1100110111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNIVS8U1_6_LC_6_12_2  (
            .in0(N__21643),
            .in1(N__25824),
            .in2(N__21877),
            .in3(N__23391),
            .lcout(\b2v_inst11.N_5572_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_12_1_LC_6_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_12_1_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_12_1_LC_6_12_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_12_1_LC_6_12_3  (
            .in0(N__21613),
            .in1(_gnd_net_),
            .in2(N__23395),
            .in3(N__21875),
            .lcout(),
            .ltout(b2v_inst11_g0_i_m2_i_a6_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SLP_S3n_ibuf_RNI4G1E7_LC_6_12_4.C_ON=1'b0;
    defparam SLP_S3n_ibuf_RNI4G1E7_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam SLP_S3n_ibuf_RNI4G1E7_LC_6_12_4.LUT_INIT=16'b0000000001000101;
    LogicCell40 SLP_S3n_ibuf_RNI4G1E7_LC_6_12_4 (
            .in0(N__21580),
            .in1(N__25823),
            .in2(N__21631),
            .in3(N__21628),
            .lcout(N_15_i_0_a4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_6_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_5_LC_6_12_5 .LUT_INIT=16'b0100010001100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_5_LC_6_12_5  (
            .in0(N__21612),
            .in1(N__21874),
            .in2(_gnd_net_),
            .in3(N__29330),
            .lcout(),
            .ltout(\b2v_inst11.g0_i_m2_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIS1UT1_5_LC_6_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIS1UT1_5_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIS1UT1_5_LC_6_12_6 .LUT_INIT=16'b0100101001000000;
    LogicCell40 \b2v_inst11.dutycycle_RNIS1UT1_5_LC_6_12_6  (
            .in0(N__21870),
            .in1(N__21589),
            .in2(N__21583),
            .in3(N__26876),
            .lcout(N_15_i_0_a4_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI4C1Q3_1_LC_6_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI4C1Q3_1_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI4C1Q3_1_LC_6_12_7 .LUT_INIT=16'b1111000011010001;
    LogicCell40 \b2v_inst11.func_state_RNI4C1Q3_1_LC_6_12_7  (
            .in0(N__21883),
            .in1(N__21876),
            .in2(N__21832),
            .in3(N__21812),
            .lcout(\b2v_inst11.un1_count_off_1_sqmuxa_8_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_0_LC_6_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_0_LC_6_13_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_0_LC_6_13_0 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \b2v_inst11.dutycycle_0_LC_6_13_0  (
            .in0(N__21778),
            .in1(N__27659),
            .in2(N__21769),
            .in3(N__21784),
            .lcout(\b2v_inst11.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36620),
            .ce(),
            .sr(N__25897));
    defparam \b2v_inst11.dutycycle_RNI8I5HB_0_LC_6_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI8I5HB_0_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI8I5HB_0_LC_6_13_1 .LUT_INIT=16'b0011001111111011;
    LogicCell40 \b2v_inst11.dutycycle_RNI8I5HB_0_LC_6_13_1  (
            .in0(N__33587),
            .in1(N__23026),
            .in2(N__33780),
            .in3(N__21751),
            .lcout(\b2v_inst11.dutycycle_eena ),
            .ltout(\b2v_inst11.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIG4U9E_0_LC_6_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIG4U9E_0_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIG4U9E_0_LC_6_13_2 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIG4U9E_0_LC_6_13_2  (
            .in0(N__21777),
            .in1(N__21765),
            .in2(N__21754),
            .in3(N__27658),
            .lcout(\b2v_inst11.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI8I5HB_1_LC_6_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI8I5HB_1_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI8I5HB_1_LC_6_13_3 .LUT_INIT=16'b0011001111111011;
    LogicCell40 \b2v_inst11.dutycycle_RNI8I5HB_1_LC_6_13_3  (
            .in0(N__33755),
            .in1(N__23025),
            .in2(N__33354),
            .in3(N__21750),
            .lcout(\b2v_inst11.dutycycle_eena_0 ),
            .ltout(\b2v_inst11.dutycycle_eena_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIRGRIE_1_LC_6_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIRGRIE_1_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIRGRIE_1_LC_6_13_4 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIRGRIE_1_LC_6_13_4  (
            .in0(N__21735),
            .in1(N__21720),
            .in2(N__21742),
            .in3(N__27657),
            .lcout(\b2v_inst11.dutycycle ),
            .ltout(\b2v_inst11.dutycycle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_1_LC_6_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_1_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_1_LC_6_13_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_1_LC_6_13_5  (
            .in0(N__33588),
            .in1(_gnd_net_),
            .in2(N__21739),
            .in3(N__29537),
            .lcout(\b2v_inst11.dutycycle_RNI_5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_1_LC_6_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_1_LC_6_13_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_1_LC_6_13_6 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \b2v_inst11.dutycycle_1_LC_6_13_6  (
            .in0(N__21736),
            .in1(N__21727),
            .in2(N__27714),
            .in3(N__21721),
            .lcout(\b2v_inst11.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36620),
            .ce(),
            .sr(N__25897));
    defparam \b2v_inst11.dutycycle_RNI_1_LC_6_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_LC_6_13_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_LC_6_13_7  (
            .in0(N__33586),
            .in1(N__29538),
            .in2(_gnd_net_),
            .in3(N__33320),
            .lcout(\b2v_inst11.g3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI_1_LC_6_14_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI_1_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI_1_LC_6_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst5.curr_state_RNI_1_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25569),
            .lcout(\b2v_inst5.curr_state_RNIZ0Z_1 ),
            .ltout(\b2v_inst5.curr_state_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIR6ES_0_LC_6_14_1 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIR6ES_0_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIR6ES_0_LC_6_14_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \b2v_inst5.curr_state_RNIR6ES_0_LC_6_14_1  (
            .in0(N__34721),
            .in1(_gnd_net_),
            .in2(N__22123),
            .in3(N__21925),
            .lcout(b2v_inst5_RSMRSTn_latmux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_fast_LC_6_14_2 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_LC_6_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.RSMRSTn_fast_LC_6_14_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_LC_6_14_2  (
            .in0(N__21928),
            .in1(N__34716),
            .in2(_gnd_net_),
            .in3(N__21904),
            .lcout(b2v_inst5_RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36625),
            .ce(N__36361),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_LC_6_14_3 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_LC_6_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.RSMRSTn_LC_6_14_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \b2v_inst5.RSMRSTn_LC_6_14_3  (
            .in0(N__21903),
            .in1(N__34712),
            .in2(_gnd_net_),
            .in3(N__21927),
            .lcout(RSMRSTn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36625),
            .ce(N__36361),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIFLPH1_1_LC_6_14_4 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIFLPH1_1_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIFLPH1_1_LC_6_14_4 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \b2v_inst5.curr_state_RNIFLPH1_1_LC_6_14_4  (
            .in0(N__21946),
            .in1(N__21901),
            .in2(N__34722),
            .in3(N__36403),
            .lcout(\b2v_inst5.curr_state_RNIFLPH1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNIJJOV_1_LC_6_14_5 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNIJJOV_1_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNIJJOV_1_LC_6_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.curr_state_RNIJJOV_1_LC_6_14_5  (
            .in0(N__21900),
            .in1(N__21945),
            .in2(N__34723),
            .in3(N__35745),
            .lcout(\b2v_inst5.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_6_14_6 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m6_i_LC_6_14_6 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m6_i_LC_6_14_6  (
            .in0(N__21926),
            .in1(N__21902),
            .in2(N__25555),
            .in3(N__34717),
            .lcout(\b2v_inst5.N_51 ),
            .ltout(\b2v_inst5.N_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_RNI2DVE1_1_LC_6_14_7 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_RNI2DVE1_1_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_RNI2DVE1_1_LC_6_14_7 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \b2v_inst5.curr_state_RNI2DVE1_1_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(N__35744),
            .in2(N__21886),
            .in3(N__30454),
            .lcout(\b2v_inst5.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI2DIN_9_LC_6_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI2DIN_9_LC_6_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNI2DIN_9_LC_6_15_0  (
            .in0(N__35813),
            .in1(N__22150),
            .in2(_gnd_net_),
            .in3(N__24669),
            .lcout(\b2v_inst11.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_9_LC_6_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_9_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_9_LC_6_15_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_9_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24673),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36629),
            .ce(N__36358),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIB49T_10_LC_6_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIB49T_10_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIB49T_10_LC_6_15_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNIB49T_10_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__22144),
            .in2(N__24658),
            .in3(N__35811),
            .lcout(\b2v_inst11.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_10_LC_6_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_10_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_10_LC_6_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_10_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24657),
            .lcout(\b2v_inst11.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36629),
            .ce(N__36358),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIK61M_11_LC_6_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIK61M_11_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIK61M_11_LC_6_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIK61M_11_LC_6_15_4  (
            .in0(N__35812),
            .in1(N__22138),
            .in2(_gnd_net_),
            .in3(N__24783),
            .lcout(\b2v_inst11.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_11_LC_6_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_11_LC_6_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_11_LC_6_15_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_11_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24787),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36629),
            .ce(N__36358),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIKNAN_2_LC_6_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIKNAN_2_LC_6_15_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNIKNAN_2_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(N__22132),
            .in2(N__24721),
            .in3(N__35810),
            .lcout(\b2v_inst11.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_2_LC_6_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_2_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_2_LC_6_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_2_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24720),
            .lcout(\b2v_inst11.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36629),
            .ce(N__36358),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_6_16_0 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_LC_6_16_0 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m8_i_LC_6_16_0  (
            .in0(N__22206),
            .in1(N__22192),
            .in2(N__22600),
            .in3(N__33684),
            .lcout(),
            .ltout(\b2v_inst200.N_56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNICM0V7_1_LC_6_16_1 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNICM0V7_1_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNICM0V7_1_LC_6_16_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.curr_state_RNICM0V7_1_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(N__22162),
            .in2(N__22126),
            .in3(N__35775),
            .lcout(\b2v_inst200.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_6_16_2 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_6_16_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a2_0_LC_6_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22333),
            .in3(N__22227),
            .lcout(N_411),
            .ltout(N_411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_6_16_3 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_6_16_3 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_0_LC_6_16_3  (
            .in0(N__22330),
            .in1(N__22264),
            .in2(N__22252),
            .in3(N__22207),
            .lcout(\b2v_inst200.m6_i_0 ),
            .ltout(\b2v_inst200.m6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_6_16_4 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m6_i_LC_6_16_4 .LUT_INIT=16'b1111000011111001;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m6_i_LC_6_16_4  (
            .in0(N__22194),
            .in1(N__22228),
            .in2(N__22243),
            .in3(N__33683),
            .lcout(),
            .ltout(\b2v_inst200.N_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_RNIGPR58_0_LC_6_16_5 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_RNIGPR58_0_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_RNIGPR58_0_LC_6_16_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst200.curr_state_RNIGPR58_0_LC_6_16_5  (
            .in0(_gnd_net_),
            .in1(N__22240),
            .in2(N__22234),
            .in3(N__35774),
            .lcout(\b2v_inst200.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst200.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_a3_0_LC_6_16_6 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_a3_0_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m8_i_a3_0_LC_6_16_6 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m8_i_a3_0_LC_6_16_6  (
            .in0(_gnd_net_),
            .in1(N__22191),
            .in2(N__22210),
            .in3(_gnd_net_),
            .lcout(N_412),
            .ltout(N_412_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_1_LC_6_16_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_1_LC_6_16_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.curr_state_1_LC_6_16_7 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \b2v_inst200.curr_state_1_LC_6_16_7  (
            .in0(N__33685),
            .in1(N__22596),
            .in2(N__22198),
            .in3(N__22193),
            .lcout(\b2v_inst200.curr_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36635),
            .ce(N__36356),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_4_LC_7_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_4_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_4_LC_7_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst36.count_RNI_4_LC_7_1_0  (
            .in0(N__27834),
            .in1(N__27802),
            .in2(N__27996),
            .in3(N__27762),
            .lcout(\b2v_inst36.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNINEG01_6_LC_7_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNINEG01_6_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNINEG01_6_LC_7_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNINEG01_6_LC_7_1_1  (
            .in0(N__22156),
            .in1(N__30696),
            .in2(_gnd_net_),
            .in3(N__27786),
            .lcout(\b2v_inst36.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_6_LC_7_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_6_LC_7_1_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_6_LC_7_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_6_LC_7_1_2  (
            .in0(N__27787),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36650),
            .ce(N__30699),
            .sr(N__30591));
    defparam \b2v_inst36.count_RNIHJCV_12_LC_7_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIHJCV_12_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIHJCV_12_LC_7_1_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIHJCV_12_LC_7_1_3  (
            .in0(N__22360),
            .in1(N__30698),
            .in2(_gnd_net_),
            .in3(N__27975),
            .lcout(\b2v_inst36.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIJ8E01_4_LC_7_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJ8E01_4_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJ8E01_4_LC_7_1_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst36.count_RNIJ8E01_4_LC_7_1_5  (
            .in0(N__27819),
            .in1(N__22372),
            .in2(_gnd_net_),
            .in3(N__30695),
            .lcout(\b2v_inst36.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_4_LC_7_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_4_LC_7_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_4_LC_7_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_4_LC_7_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27820),
            .lcout(\b2v_inst36.count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36650),
            .ce(N__30699),
            .sr(N__30591));
    defparam \b2v_inst36.count_RNITNJ01_9_LC_7_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNITNJ01_9_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNITNJ01_9_LC_7_1_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNITNJ01_9_LC_7_1_7  (
            .in0(N__22366),
            .in1(N__30697),
            .in2(_gnd_net_),
            .in3(N__27747),
            .lcout(\b2v_inst36.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_14_LC_7_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_14_LC_7_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_14_LC_7_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_14_LC_7_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27934),
            .lcout(\b2v_inst36.count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36644),
            .ce(N__30732),
            .sr(N__30587));
    defparam \b2v_inst36.count_9_LC_7_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_9_LC_7_2_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_9_LC_7_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_9_LC_7_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27748),
            .lcout(\b2v_inst36.count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36644),
            .ce(N__30732),
            .sr(N__30587));
    defparam \b2v_inst36.count_12_LC_7_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_12_LC_7_2_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_12_LC_7_2_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_12_LC_7_2_5  (
            .in0(N__27976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36644),
            .ce(N__30732),
            .sr(N__30587));
    defparam \b2v_inst36.curr_state_RNI8TT2_0_LC_7_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI8TT2_0_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI8TT2_0_LC_7_3_0 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \b2v_inst36.curr_state_RNI8TT2_0_LC_7_3_0  (
            .in0(N__22398),
            .in1(_gnd_net_),
            .in2(N__25354),
            .in3(N__25289),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_RNI8TT2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_RNIUDI9_LC_7_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_RNIUDI9_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.DSW_PWROK_RNIUDI9_LC_7_3_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst36.DSW_PWROK_RNIUDI9_LC_7_3_1  (
            .in0(N__22414),
            .in1(_gnd_net_),
            .in2(N__22354),
            .in3(N__35933),
            .lcout(DSW_PWROK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_0_LC_7_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_0_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_0_LC_7_3_2 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \b2v_inst36.curr_state_0_LC_7_3_2  (
            .in0(N__30845),
            .in1(N__22393),
            .in2(N__25352),
            .in3(N__25287),
            .lcout(\b2v_inst36.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36638),
            .ce(N__36367),
            .sr(_gnd_net_));
    defparam \b2v_inst36.DSW_PWROK_LC_7_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.DSW_PWROK_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.DSW_PWROK_LC_7_3_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \b2v_inst36.DSW_PWROK_LC_7_3_3  (
            .in0(N__25286),
            .in1(_gnd_net_),
            .in2(N__22399),
            .in3(N__25340),
            .lcout(\b2v_inst36.DSW_PWROK_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36638),
            .ce(N__36367),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_7_3_4 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m4_LC_7_3_4 .LUT_INIT=16'b0010001011000000;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m4_LC_7_3_4  (
            .in0(N__30844),
            .in1(N__22397),
            .in2(N__25353),
            .in3(N__25285),
            .lcout(),
            .ltout(\b2v_inst36.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI2MTL_0_LC_7_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI2MTL_0_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI2MTL_0_LC_7_3_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.curr_state_RNI2MTL_0_LC_7_3_5  (
            .in0(_gnd_net_),
            .in1(N__22408),
            .in2(N__22402),
            .in3(N__35932),
            .lcout(\b2v_inst36.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI_0_LC_7_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI_0_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI_0_LC_7_3_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst36.curr_state_RNI_0_LC_7_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22378),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.N_2939_i ),
            .ltout(\b2v_inst36.N_2939_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_7_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_7_1_0__m6_LC_7_3_7 .LUT_INIT=16'b0100000011100000;
    LogicCell40 \b2v_inst36.curr_state_7_1_0__m6_LC_7_3_7  (
            .in0(N__25288),
            .in1(N__25347),
            .in2(N__22375),
            .in3(N__30843),
            .lcout(\b2v_inst36.curr_state_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_11_LC_7_4_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_11_LC_7_4_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_11_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_11_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31444),
            .lcout(\b2v_inst5.count_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36631),
            .ce(N__31928),
            .sr(N__32173));
    defparam \b2v_inst5.count_12_LC_7_4_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_12_LC_7_4_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_12_LC_7_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_12_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31411),
            .lcout(\b2v_inst5.count_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36631),
            .ce(N__31928),
            .sr(N__32173));
    defparam \b2v_inst5.count_14_LC_7_4_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_14_LC_7_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_14_LC_7_4_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst5.count_14_LC_7_4_2  (
            .in0(_gnd_net_),
            .in1(N__31324),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36631),
            .ce(N__31928),
            .sr(N__32173));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_5_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__28657),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_5_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__25450),
            .in2(N__22507),
            .in3(N__22444),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_5_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__22671),
            .in2(N__22660),
            .in3(N__22441),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_5_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__32548),
            .in2(N__22558),
            .in3(N__22438),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_5_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__22546),
            .in2(N__32556),
            .in3(N__22435),
            .lcout(\b2v_inst11.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_5_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_5_5  (
            .in0(N__25474),
            .in1(N__22536),
            .in2(N__22426),
            .in3(N__22432),
            .lcout(\b2v_inst11.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un131_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_5_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22525),
            .in3(N__22429),
            .lcout(\b2v_inst11.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__22537),
            .in2(_gnd_net_),
            .in3(N__32547),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__28626),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__25495),
            .in2(N__25593),
            .in3(N__22417),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__25589),
            .in2(N__25435),
            .in3(N__22549),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__25642),
            .in2(N__32586),
            .in3(N__22540),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__32582),
            .in2(N__25633),
            .in3(N__22528),
            .lcout(\b2v_inst11.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_6_5  (
            .in0(N__32552),
            .in1(N__25621),
            .in2(N__25594),
            .in3(N__22516),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un124_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25612),
            .in3(N__22513),
            .lcout(\b2v_inst11.mult1_un124_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un124_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22510),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIPFFQ6_LC_7_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIPFFQ6_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIPFFQ6_LC_7_7_0 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_4_c_RNIPFFQ6_LC_7_7_0  (
            .in0(N__22497),
            .in1(N__23067),
            .in2(N__22456),
            .in3(N__27147),
            .lcout(b2v_inst11_dutycycle_set_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_7_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_7_7_1  (
            .in0(N__28677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_14_LC_7_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_14_LC_7_7_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_14_LC_7_7_2  (
            .in0(N__29726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22686),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_7_3  (
            .in0(N__22672),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32546),
            .lcout(\b2v_inst11.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_7_7_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_9_LC_7_7_5 .LUT_INIT=16'b1010100011101010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_9_LC_7_7_5  (
            .in0(N__26335),
            .in1(N__26449),
            .in2(N__26823),
            .in3(N__22648),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_13_LC_7_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_13_LC_7_7_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_13_LC_7_7_6  (
            .in0(N__26450),
            .in1(N__28900),
            .in2(N__22642),
            .in3(N__29223),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_7_7_7 .C_ON=1'b0;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_7_7_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst200.curr_state_13_2_0__m11_0_a3_0_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__22639),
            .in2(_gnd_net_),
            .in3(N__22627),
            .lcout(\b2v_inst200.m11_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIB6L91_LC_7_8_1 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIB6L91_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_c_RNIB6L91_LC_7_8_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_c_RNIB6L91_LC_7_8_1  (
            .in0(N__31491),
            .in1(N__31131),
            .in2(N__31152),
            .in3(N__32094),
            .lcout(\b2v_inst5.count_rst_10 ),
            .ltout(\b2v_inst5.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIP7CS2_4_LC_7_8_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIP7CS2_4_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIP7CS2_4_LC_7_8_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst5.count_RNIP7CS2_4_LC_7_8_2  (
            .in0(N__31835),
            .in1(_gnd_net_),
            .in2(N__22570),
            .in3(N__22770),
            .lcout(\b2v_inst5.un2_count_1_axb_4 ),
            .ltout(\b2v_inst5.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_4_LC_7_8_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_4_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_4_LC_7_8_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \b2v_inst5.count_4_LC_7_8_3  (
            .in0(N__31492),
            .in1(N__31132),
            .in2(N__22567),
            .in3(N__32096),
            .lcout(\b2v_inst5.count_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36608),
            .ce(N__31941),
            .sr(N__32135));
    defparam \b2v_inst5.count_8_LC_7_8_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_8_LC_7_8_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_8_LC_7_8_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst5.count_8_LC_7_8_4  (
            .in0(N__32095),
            .in1(N__31493),
            .in2(N__31066),
            .in3(N__31085),
            .lcout(\b2v_inst5.count_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36608),
            .ce(N__31941),
            .sr(N__32135));
    defparam \b2v_inst5.count_RNI1KGS2_8_LC_7_8_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI1KGS2_8_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI1KGS2_8_LC_7_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNI1KGS2_8_LC_7_8_5  (
            .in0(N__22564),
            .in1(N__31836),
            .in2(_gnd_net_),
            .in3(N__28282),
            .lcout(\b2v_inst5.countZ0Z_8 ),
            .ltout(\b2v_inst5.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIP7CS2_0_4_LC_7_8_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIP7CS2_0_4_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIP7CS2_0_4_LC_7_8_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \b2v_inst5.count_RNIP7CS2_0_4_LC_7_8_6  (
            .in0(N__31942),
            .in1(N__22780),
            .in2(N__22774),
            .in3(N__22771),
            .lcout(),
            .ltout(\b2v_inst5.un12_clk_100khz_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIAEONB_2_LC_7_8_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIAEONB_2_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIAEONB_2_LC_7_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.count_RNIAEONB_2_LC_7_8_7  (
            .in0(N__28294),
            .in1(N__28048),
            .in2(N__22762),
            .in3(N__31615),
            .lcout(\b2v_inst5.un12_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_7_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_9_LC_7_9_0 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_9_LC_7_9_0  (
            .in0(N__29491),
            .in1(N__26425),
            .in2(N__26836),
            .in3(N__26155),
            .lcout(),
            .ltout(\b2v_inst11.N_8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_7_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_10_LC_7_9_1 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_10_LC_7_9_1  (
            .in0(N__26308),
            .in1(N__26435),
            .in2(N__22759),
            .in3(N__29199),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_2Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_10_LC_7_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_10_LC_7_9_2 .LUT_INIT=16'b1011010101001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_10_LC_7_9_2  (
            .in0(N__29200),
            .in1(N__22756),
            .in2(N__22744),
            .in3(N__22693),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNITS10B_14_LC_7_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNITS10B_14_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNITS10B_14_LC_7_9_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst11.dutycycle_RNITS10B_14_LC_7_9_3  (
            .in0(N__22737),
            .in1(N__22726),
            .in2(N__22717),
            .in3(N__25864),
            .lcout(\b2v_inst11.dutycycleZ0Z_12 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_7_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_11_LC_7_9_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_11_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22696),
            .in3(N__29116),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_6_LC_7_9_5 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_6_LC_7_9_5  (
            .in0(N__26153),
            .in1(N__29490),
            .in2(_gnd_net_),
            .in3(N__26808),
            .lcout(\b2v_inst11.N_15_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_7_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_9_LC_7_9_6 .LUT_INIT=16'b0000001100111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_9_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__26426),
            .in2(N__29530),
            .in3(N__26154),
            .lcout(\b2v_inst11.dutycycle_RNI_3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_7_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_9_LC_7_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_9_LC_7_9_7  (
            .in0(N__26156),
            .in1(N__26436),
            .in2(N__29397),
            .in3(N__22849),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI5K4VA_9_LC_7_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI5K4VA_9_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI5K4VA_9_LC_7_10_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI5K4VA_9_LC_7_10_0  (
            .in0(N__25836),
            .in1(N__22809),
            .in2(N__22828),
            .in3(N__22834),
            .lcout(\b2v_inst11.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIRP00B_13_LC_7_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIRP00B_13_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIRP00B_13_LC_7_10_1 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \b2v_inst11.dutycycle_RNIRP00B_13_LC_7_10_1  (
            .in0(N__23271),
            .in1(N__22788),
            .in2(N__22801),
            .in3(N__25837),
            .lcout(\b2v_inst11.dutycycleZ0Z_8 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_13_LC_7_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_13_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_13_LC_7_10_2 .LUT_INIT=16'b1100000011010101;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_13_LC_7_10_2  (
            .in0(N__25835),
            .in1(N__23242),
            .in2(N__22843),
            .in3(N__26570),
            .lcout(),
            .ltout(\b2v_inst11.N_153_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIMBHI8_13_LC_7_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_13_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_13_LC_7_10_3 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIMBHI8_13_LC_7_10_3  (
            .in0(N__27671),
            .in1(N__23181),
            .in2(N__22840),
            .in3(N__23066),
            .lcout(\b2v_inst11.dutycycle_en_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_9_LC_7_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_9_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_9_LC_7_10_4 .LUT_INIT=16'b1100000011010101;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_9_LC_7_10_4  (
            .in0(N__25834),
            .in1(N__23241),
            .in2(N__26451),
            .in3(N__26569),
            .lcout(),
            .ltout(\b2v_inst11.N_156_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIMBHI8_9_LC_7_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_9_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_9_LC_7_10_5 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIMBHI8_9_LC_7_10_5  (
            .in0(N__27670),
            .in1(N__23180),
            .in2(N__22837),
            .in3(N__23065),
            .lcout(\b2v_inst11.dutycycle_e_1_9 ),
            .ltout(\b2v_inst11.dutycycle_e_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_9_LC_7_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_9_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_9_LC_7_10_6 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \b2v_inst11.dutycycle_9_LC_7_10_6  (
            .in0(N__25838),
            .in1(N__22824),
            .in2(N__22813),
            .in3(N__22810),
            .lcout(\b2v_inst11.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36607),
            .ce(),
            .sr(N__25946));
    defparam \b2v_inst11.dutycycle_13_LC_7_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_13_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_13_LC_7_10_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \b2v_inst11.dutycycle_13_LC_7_10_7  (
            .in0(N__22797),
            .in1(N__22789),
            .in2(N__23275),
            .in3(N__25839),
            .lcout(\b2v_inst11.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36607),
            .ce(),
            .sr(N__25946));
    defparam \b2v_inst11.dutycycle_RNI0084B_8_LC_7_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI0084B_8_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI0084B_8_LC_7_11_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \b2v_inst11.dutycycle_RNI0084B_8_LC_7_11_0  (
            .in0(N__23055),
            .in1(N__22880),
            .in2(N__22861),
            .in3(N__23076),
            .lcout(\b2v_inst11.dutycycleZ0Z_5 ),
            .ltout(\b2v_inst11.dutycycleZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_8_LC_7_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_8_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_8_LC_7_11_1 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_8_LC_7_11_1  (
            .in0(N__23234),
            .in1(N__23173),
            .in2(N__23263),
            .in3(N__23260),
            .lcout(\b2v_inst11.dutycycle_e_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNICDJJ5_10_LC_7_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_10_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNICDJJ5_10_LC_7_11_2 .LUT_INIT=16'b1100000011010101;
    LogicCell40 \b2v_inst11.dutycycle_RNICDJJ5_10_LC_7_11_2  (
            .in0(N__25860),
            .in1(N__23235),
            .in2(N__29217),
            .in3(N__26643),
            .lcout(),
            .ltout(\b2v_inst11.N_154_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIMBHI8_10_LC_7_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_10_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIMBHI8_10_LC_7_11_3 .LUT_INIT=16'b0010000010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIMBHI8_10_LC_7_11_3  (
            .in0(N__27672),
            .in1(N__23174),
            .in2(N__23083),
            .in3(N__23054),
            .lcout(\b2v_inst11.dutycycle_en_4 ),
            .ltout(\b2v_inst11.dutycycle_en_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIEOB3B_10_LC_7_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIEOB3B_10_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIEOB3B_10_LC_7_11_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIEOB3B_10_LC_7_11_4  (
            .in0(N__25861),
            .in1(N__22896),
            .in2(N__23080),
            .in3(N__22909),
            .lcout(\b2v_inst11.dutycycleZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_8_LC_7_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_8_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_8_LC_7_11_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \b2v_inst11.dutycycle_8_LC_7_11_5  (
            .in0(N__23077),
            .in1(N__22857),
            .in2(N__22885),
            .in3(N__23056),
            .lcout(\b2v_inst11.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36613),
            .ce(),
            .sr(N__25980));
    defparam \b2v_inst11.dutycycle_10_LC_7_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_10_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_10_LC_7_11_6 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \b2v_inst11.dutycycle_10_LC_7_11_6  (
            .in0(N__25863),
            .in1(N__22915),
            .in2(N__22900),
            .in3(N__22908),
            .lcout(\b2v_inst11.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36613),
            .ce(),
            .sr(N__25980));
    defparam \b2v_inst11.dutycycle_RNI1KT13_8_LC_7_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI1KT13_8_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI1KT13_8_LC_7_11_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst11.dutycycle_RNI1KT13_8_LC_7_11_7  (
            .in0(N__22881),
            .in1(N__22870),
            .in2(N__27701),
            .in3(N__25862),
            .lcout(\b2v_inst11.dutycycle_RNI1KT13Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI8JP5_0_LC_7_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI8JP5_0_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI8JP5_0_LC_7_12_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \b2v_inst11.func_state_RNI8JP5_0_LC_7_12_0  (
            .in0(N__23389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24638),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI6P011_1_LC_7_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI6P011_1_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI6P011_1_LC_7_12_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.func_state_RNI6P011_1_LC_7_12_1  (
            .in0(N__24514),
            .in1(N__24931),
            .in2(N__24400),
            .in3(N__23672),
            .lcout(\b2v_inst11.N_295 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIU8G3G_2_LC_7_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIU8G3G_2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIU8G3G_2_LC_7_12_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_RNIU8G3G_2_LC_7_12_2  (
            .in0(N__23919),
            .in1(N__27668),
            .in2(N__23947),
            .in3(N__23934),
            .lcout(dutycycle_RNIU8G3G_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIF6NL_LC_7_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIF6NL_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIF6NL_LC_7_12_4 .LUT_INIT=16'b1110111110101010;
    LogicCell40 \b2v_inst11.un1_dutycycle_94_cry_1_c_RNIF6NL_LC_7_12_4  (
            .in0(N__24370),
            .in1(N__24226),
            .in2(N__24217),
            .in3(N__24126),
            .lcout(),
            .ltout(\b2v_inst11.g1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.func_state_RNI5M9V2_1_LC_7_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.func_state_RNI5M9V2_1_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.func_state_RNI5M9V2_1_LC_7_12_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \b2v_inst11.func_state_RNI5M9V2_1_LC_7_12_5  (
            .in0(N__23876),
            .in1(_gnd_net_),
            .in2(N__23956),
            .in3(N__23953),
            .lcout(\b2v_inst11.g1 ),
            .ltout(\b2v_inst11.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_2_LC_7_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_2_LC_7_12_6 .SEQ_MODE=4'b1011;
    defparam \b2v_inst11.dutycycle_2_LC_7_12_6 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \b2v_inst11.dutycycle_2_LC_7_12_6  (
            .in0(N__23920),
            .in1(N__27669),
            .in2(N__23938),
            .in3(N__23935),
            .lcout(\b2v_inst11.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36621),
            .ce(),
            .sr(N__25945));
    defparam \b2v_inst5.RSMRSTn_fast_RNIVS8U1_LC_7_12_7 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_RNIVS8U1_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_fast_RNIVS8U1_LC_7_12_7 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_RNIVS8U1_LC_7_12_7  (
            .in0(N__23875),
            .in1(N__23671),
            .in2(N__23531),
            .in3(N__23388),
            .lcout(\b2v_inst5.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_LC_7_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_LC_7_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__32439),
            .in2(N__32400),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\b2v_inst11.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_7_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_7_13_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_1_c_RNIIIQD_LC_7_13_1  (
            .in0(N__27448),
            .in1(N__32357),
            .in2(_gnd_net_),
            .in3(N__24706),
            .lcout(\b2v_inst11.count_1_2 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_1 ),
            .carryout(\b2v_inst11.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_7_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_7_13_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_2_c_RNIJKRD_LC_7_13_2  (
            .in0(N__27452),
            .in1(N__32306),
            .in2(_gnd_net_),
            .in3(N__24703),
            .lcout(\b2v_inst11.count_1_3 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_2 ),
            .carryout(\b2v_inst11.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_7_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_7_13_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_3_c_RNIKMSD_LC_7_13_3  (
            .in0(N__27449),
            .in1(N__32940),
            .in2(_gnd_net_),
            .in3(N__24700),
            .lcout(\b2v_inst11.count_1_4 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_3 ),
            .carryout(\b2v_inst11.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_7_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_7_13_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_4_c_RNILOTD_LC_7_13_4  (
            .in0(N__27453),
            .in1(N__32901),
            .in2(_gnd_net_),
            .in3(N__24697),
            .lcout(\b2v_inst11.count_1_5 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_4 ),
            .carryout(\b2v_inst11.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_7_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_7_13_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_5_c_RNIMQUD_LC_7_13_5  (
            .in0(N__27450),
            .in1(N__32847),
            .in2(_gnd_net_),
            .in3(N__24694),
            .lcout(\b2v_inst11.count_1_6 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_5 ),
            .carryout(\b2v_inst11.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_7_13_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_7_13_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_6_c_RNINSVD_LC_7_13_6  (
            .in0(N__27454),
            .in1(N__32804),
            .in2(_gnd_net_),
            .in3(N__24679),
            .lcout(\b2v_inst11.count_1_7 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_6 ),
            .carryout(\b2v_inst11.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_7_13_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_7_13_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_7_c_RNIOU0E_LC_7_13_7  (
            .in0(N__27451),
            .in1(N__32766),
            .in2(_gnd_net_),
            .in3(N__24676),
            .lcout(\b2v_inst11.count_1_8 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_7 ),
            .carryout(\b2v_inst11.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_7_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_7_14_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_8_c_RNIP02E_LC_7_14_0  (
            .in0(N__27438),
            .in1(N__32711),
            .in2(_gnd_net_),
            .in3(N__24661),
            .lcout(\b2v_inst11.count_1_9 ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\b2v_inst11.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_7_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_7_14_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_9_c_RNIQ23E_LC_7_14_1  (
            .in0(N__27455),
            .in1(N__32657),
            .in2(_gnd_net_),
            .in3(N__24646),
            .lcout(\b2v_inst11.count_1_10 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_9 ),
            .carryout(\b2v_inst11.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_7_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_7_14_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_10_c_RNI24R6_LC_7_14_2  (
            .in0(N__27437),
            .in1(N__32615),
            .in2(_gnd_net_),
            .in3(N__24775),
            .lcout(\b2v_inst11.count_1_11 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_10 ),
            .carryout(\b2v_inst11.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_7_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_7_14_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_11_c_RNI36S6_LC_7_14_3  (
            .in0(N__27456),
            .in1(N__33120),
            .in2(_gnd_net_),
            .in3(N__24772),
            .lcout(\b2v_inst11.count_1_12 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_11 ),
            .carryout(\b2v_inst11.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_7_14_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_7_14_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_12_c_RNI48T6_LC_7_14_4  (
            .in0(N__27439),
            .in1(N__33087),
            .in2(_gnd_net_),
            .in3(N__24769),
            .lcout(\b2v_inst11.count_1_13 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_12 ),
            .carryout(\b2v_inst11.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_7_14_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_7_14_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_13_c_RNI5AU6_LC_7_14_5  (
            .in0(N__27457),
            .in1(N__33051),
            .in2(_gnd_net_),
            .in3(N__24766),
            .lcout(\b2v_inst11.count_1_14 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_count_cry_13 ),
            .carryout(\b2v_inst11.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_7_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_7_14_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst11.un1_count_cry_14_c_RNI6CV6_LC_7_14_6  (
            .in0(N__27440),
            .in1(N__33018),
            .in2(_gnd_net_),
            .in3(N__24763),
            .lcout(\b2v_inst11.un1_count_cry_14_c_RNI6CVZ0Z6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQF4M_14_LC_7_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQF4M_14_LC_7_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIQF4M_14_LC_7_14_7  (
            .in0(N__35901),
            .in1(N__24727),
            .in2(_gnd_net_),
            .in3(N__24738),
            .lcout(\b2v_inst11.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_7_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIQ0EN_5_LC_7_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIQ0EN_5_LC_7_15_0  (
            .in0(N__35886),
            .in1(N__24745),
            .in2(_gnd_net_),
            .in3(N__24756),
            .lcout(\b2v_inst11.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_5_LC_7_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_5_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_5_LC_7_15_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_5_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24760),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36637),
            .ce(N__36355),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_14_LC_7_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_14_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_14_LC_7_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_14_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24739),
            .lcout(\b2v_inst11.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36637),
            .ce(N__36355),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIS3FN_6_LC_7_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIS3FN_6_LC_7_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIS3FN_6_LC_7_15_4  (
            .in0(N__35885),
            .in1(N__24973),
            .in2(_gnd_net_),
            .in3(N__24984),
            .lcout(\b2v_inst11.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_6_LC_7_15_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_6_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_6_LC_7_15_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_6_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24988),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36637),
            .ce(N__36355),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNISI5M_15_LC_7_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNISI5M_15_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNISI5M_15_LC_7_15_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNISI5M_15_LC_7_15_6  (
            .in0(N__24955),
            .in1(N__35870),
            .in2(_gnd_net_),
            .in3(N__24963),
            .lcout(\b2v_inst11.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_15_LC_7_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_15_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_15_LC_7_15_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_15_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24967),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36637),
            .ce(N__36355),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_16_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_16_0 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_RNICRLO_LC_7_16_0  (
            .in0(N__36409),
            .in1(N__24940),
            .in2(N__32989),
            .in3(N__29877),
            .lcout(),
            .ltout(\b2v_inst11.pwm_out_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNIEV5S_LC_7_16_1 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNIEV5S_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNIEV5S_LC_7_16_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst11.pwm_out_RNIEV5S_LC_7_16_1  (
            .in0(N__29876),
            .in1(_gnd_net_),
            .in2(N__24949),
            .in3(N__27484),
            .lcout(PWRBTN_LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst20.tmp_1_rep1_LC_7_16_3 .C_ON=1'b0;
    defparam \b2v_inst20.tmp_1_rep1_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst20.tmp_1_rep1_LC_7_16_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst20.tmp_1_rep1_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__24901),
            .in2(_gnd_net_),
            .in3(N__24836),
            .lcout(SYNTHESIZED_WIRE_1keep_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36643),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_16_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_0_LC_7_16_4  (
            .in0(N__35917),
            .in1(N__29875),
            .in2(_gnd_net_),
            .in3(N__29838),
            .lcout(\b2v_inst11.pwm_out_1_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.G_146_LC_7_16_7 .C_ON=1'b0;
    defparam \b2v_inst36.G_146_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.G_146_LC_7_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \b2v_inst36.G_146_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__24900),
            .in2(_gnd_net_),
            .in3(N__24835),
            .lcout(G_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_0_LC_8_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_0_LC_8_1_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_0_LC_8_1_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst36.count_0_LC_8_1_0  (
            .in0(N__27349),
            .in1(N__30959),
            .in2(_gnd_net_),
            .in3(N__30842),
            .lcout(\b2v_inst36.count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36657),
            .ce(N__30700),
            .sr(N__30590));
    defparam \b2v_inst36.count_RNI471O_1_LC_8_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI471O_1_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI471O_1_LC_8_1_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst36.count_RNI471O_1_LC_8_1_1  (
            .in0(N__25009),
            .in1(N__25021),
            .in2(_gnd_net_),
            .in3(N__30701),
            .lcout(),
            .ltout(\b2v_inst36.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI471O_2_1_LC_8_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI471O_2_1_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI471O_2_1_LC_8_1_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst36.count_RNI471O_2_1_LC_8_1_2  (
            .in0(N__28027),
            .in1(N__27904),
            .in2(N__25045),
            .in3(N__28150),
            .lcout(),
            .ltout(\b2v_inst36.un12_clk_100khz_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNISMPL1_1_LC_8_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNISMPL1_1_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNISMPL1_1_LC_8_1_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNISMPL1_1_LC_8_1_3  (
            .in0(N__25000),
            .in1(N__25042),
            .in2(N__25033),
            .in3(N__30382),
            .lcout(\b2v_inst36.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI361O_0_LC_8_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI361O_0_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI361O_0_LC_8_1_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst36.count_RNI361O_0_LC_8_1_4  (
            .in0(N__25030),
            .in1(N__24994),
            .in2(_gnd_net_),
            .in3(N__30693),
            .lcout(\b2v_inst36.countZ0Z_0 ),
            .ltout(\b2v_inst36.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_1_LC_8_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_1_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_1_LC_8_1_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst36.count_RNI_1_LC_8_1_5  (
            .in0(N__30957),
            .in1(_gnd_net_),
            .in2(N__25024),
            .in3(N__27364),
            .lcout(\b2v_inst36.count_rst_13 ),
            .ltout(\b2v_inst36.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI471O_0_1_LC_8_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI471O_0_1_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI471O_0_1_LC_8_1_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNI471O_0_1_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(N__25008),
            .in2(N__25015),
            .in3(N__30694),
            .lcout(\b2v_inst36.un2_count_1_axb_1 ),
            .ltout(\b2v_inst36.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_1_LC_8_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_1_LC_8_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_1_LC_8_1_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \b2v_inst36.count_1_LC_8_1_7  (
            .in0(N__30958),
            .in1(_gnd_net_),
            .in2(N__25012),
            .in3(N__27348),
            .lcout(\b2v_inst36.count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36657),
            .ce(N__30700),
            .sr(N__30590));
    defparam \b2v_inst36.count_RNIOFOT_0_14_LC_8_2_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIOFOT_0_14_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIOFOT_0_14_LC_8_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst36.count_RNIOFOT_0_14_LC_8_2_0  (
            .in0(N__28060),
            .in1(N__27350),
            .in2(N__27952),
            .in3(N__28108),
            .lcout(\b2v_inst36.un12_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_0_LC_8_2_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_0_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_0_LC_8_2_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \b2v_inst36.count_RNI_0_LC_8_2_1  (
            .in0(N__27351),
            .in1(N__30912),
            .in2(_gnd_net_),
            .in3(N__30811),
            .lcout(\b2v_inst36.count_rst_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_2 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_2 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_c_RNIQ3J1_LC_8_2_2  (
            .in0(N__30813),
            .in1(N__28026),
            .in2(N__30956),
            .in3(N__28008),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIFGBV_11_LC_8_2_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIFGBV_11_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIFGBV_11_LC_8_2_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIFGBV_11_LC_8_2_3  (
            .in0(_gnd_net_),
            .in1(N__25078),
            .in2(N__25084),
            .in3(N__30661),
            .lcout(\b2v_inst36.countZ0Z_11 ),
            .ltout(\b2v_inst36.countZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_11_LC_8_2_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_11_LC_8_2_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_11_LC_8_2_4 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \b2v_inst36.count_11_LC_8_2_4  (
            .in0(N__30814),
            .in1(N__30927),
            .in2(N__25081),
            .in3(N__28009),
            .lcout(\b2v_inst36.count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36652),
            .ce(N__30730),
            .sr(N__30592));
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_8_2_5 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_8_2_5 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_RNIAQA8_LC_8_2_5  (
            .in0(N__27849),
            .in1(N__30399),
            .in2(N__30960),
            .in3(N__30812),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIF2C01_2_LC_8_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIF2C01_2_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIF2C01_2_LC_8_2_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNIF2C01_2_LC_8_2_6  (
            .in0(N__30660),
            .in1(_gnd_net_),
            .in2(N__25072),
            .in3(N__25066),
            .lcout(\b2v_inst36.countZ0Z_2 ),
            .ltout(\b2v_inst36.countZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_2_LC_8_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_2_LC_8_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_2_LC_8_2_7 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.count_2_LC_8_2_7  (
            .in0(N__27850),
            .in1(N__30916),
            .in2(N__25069),
            .in3(N__30815),
            .lcout(\b2v_inst36.count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36652),
            .ce(N__30730),
            .sr(N__30592));
    defparam \b2v_inst36.curr_state_RNI3NTL_1_LC_8_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI3NTL_1_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI3NTL_1_LC_8_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst36.curr_state_RNI3NTL_1_LC_8_3_0  (
            .in0(N__25051),
            .in1(N__25060),
            .in2(_gnd_net_),
            .in3(N__35930),
            .lcout(\b2v_inst36.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst36.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNIKEBL_1_LC_8_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNIKEBL_1_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNIKEBL_1_LC_8_3_1 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \b2v_inst36.curr_state_RNIKEBL_1_LC_8_3_1  (
            .in0(N__30536),
            .in1(N__25365),
            .in2(N__25054),
            .in3(N__36407),
            .lcout(\b2v_inst36.count_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_1_LC_8_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_1_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst36.curr_state_1_LC_8_3_2 .LUT_INIT=16'b0100000011100000;
    LogicCell40 \b2v_inst36.curr_state_1_LC_8_3_2  (
            .in0(N__25291),
            .in1(N__25336),
            .in2(N__25369),
            .in3(N__30856),
            .lcout(\b2v_inst36.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36646),
            .ce(N__36368),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI0A86_1_LC_8_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI0A86_1_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI0A86_1_LC_8_3_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \b2v_inst36.curr_state_RNI0A86_1_LC_8_3_3  (
            .in0(N__35931),
            .in1(N__25364),
            .in2(N__25351),
            .in3(N__25290),
            .lcout(\b2v_inst36.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_3_4 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_3_4 .LUT_INIT=16'b0000000001100000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_c_RNIF4G8_LC_8_3_4  (
            .in0(N__31004),
            .in1(N__30765),
            .in2(N__30980),
            .in3(N__30857),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIPHH01_7_LC_8_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIPHH01_7_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIPHH01_7_LC_8_3_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \b2v_inst36.count_RNIPHH01_7_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__30724),
            .in2(N__25264),
            .in3(N__30745),
            .lcout(\b2v_inst36.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.curr_state_RNI_1_LC_8_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.curr_state_RNI_1_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.curr_state_RNI_1_LC_8_3_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst36.curr_state_RNI_1_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30535),
            .lcout(\b2v_inst36.N_2942_i ),
            .ltout(\b2v_inst36.N_2942_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_3_7 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_c_RNIG6H8_LC_8_3_7  (
            .in0(N__30855),
            .in1(N__27903),
            .in2(N__25261),
            .in3(N__27876),
            .lcout(\b2v_inst36.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_RNIFF751_9_LC_8_4_0 .C_ON=1'b0;
    defparam \b2v_inst200.count_RNIFF751_9_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst200.count_RNIFF751_9_LC_8_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst200.count_RNIFF751_9_LC_8_4_0  (
            .in0(N__25240),
            .in1(N__25225),
            .in2(_gnd_net_),
            .in3(N__25202),
            .lcout(\b2v_inst200.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst200.count_9_LC_8_4_1 .C_ON=1'b0;
    defparam \b2v_inst200.count_9_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst200.count_9_LC_8_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst200.count_9_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25239),
            .lcout(\b2v_inst200.count_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36639),
            .ce(N__25157),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIOFOT_14_LC_8_4_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIOFOT_14_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIOFOT_14_LC_8_4_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNIOFOT_14_LC_8_4_2  (
            .in0(N__25099),
            .in1(N__30680),
            .in2(_gnd_net_),
            .in3(N__27933),
            .lcout(\b2v_inst36.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIL7E23_11_LC_8_4_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL7E23_11_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL7E23_11_LC_8_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst5.count_RNIL7E23_11_LC_8_4_3  (
            .in0(N__31443),
            .in1(N__25090),
            .in2(_gnd_net_),
            .in3(N__31911),
            .lcout(\b2v_inst5.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNINAF23_12_LC_8_4_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNINAF23_12_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNINAF23_12_LC_8_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst5.count_RNINAF23_12_LC_8_4_4  (
            .in0(N__31912),
            .in1(N__25423),
            .in2(_gnd_net_),
            .in3(N__31410),
            .lcout(\b2v_inst5.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIRGH23_14_LC_8_4_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRGH23_14_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRGH23_14_LC_8_4_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIRGH23_14_LC_8_4_5  (
            .in0(N__25414),
            .in1(N__31913),
            .in2(_gnd_net_),
            .in3(N__31323),
            .lcout(\b2v_inst5.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNITJI23_15_LC_8_4_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNITJI23_15_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNITJI23_15_LC_8_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \b2v_inst5.count_RNITJI23_15_LC_8_4_6  (
            .in0(N__31914),
            .in1(N__31285),
            .in2(_gnd_net_),
            .in3(N__31267),
            .lcout(\b2v_inst5.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_5_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__28681),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_5_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_5_1  (
            .in0(_gnd_net_),
            .in1(N__25489),
            .in2(N__25517),
            .in3(N__25408),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_5_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__25405),
            .in2(N__25519),
            .in3(N__25399),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_5_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__25396),
            .in2(N__25483),
            .in3(N__25390),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_5_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__25387),
            .in2(N__25482),
            .in3(N__25381),
            .lcout(\b2v_inst11.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_5_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_5_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_5_5  (
            .in0(N__32466),
            .in1(N__25378),
            .in2(N__25518),
            .in3(N__25372),
            .lcout(\b2v_inst11.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un138_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_5_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_5_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_5_6  (
            .in0(N__25528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25522),
            .lcout(\b2v_inst11.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_5_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25475),
            .lcout(\b2v_inst11.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_6_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_6_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_6_0  (
            .in0(N__28576),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_8_6_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_8_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28656),
            .lcout(\b2v_inst11.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_6_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25473),
            .lcout(\b2v_inst11.mult1_un131_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_6_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_6_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_6_4  (
            .in0(N__28627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_6_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_6_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_6_5  (
            .in0(N__28708),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_7_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__28575),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_7_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__25675),
            .in2(N__28506),
            .in3(N__25426),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_7_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__28502),
            .in2(N__28360),
            .in3(N__25636),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_7_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__28348),
            .in2(N__31689),
            .in3(N__25624),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_7_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__31685),
            .in2(N__28339),
            .in3(N__25615),
            .lcout(\b2v_inst11.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_7_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_7_5  (
            .in0(N__32578),
            .in1(N__28327),
            .in2(N__28507),
            .in3(N__25603),
            .lcout(\b2v_inst11.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un117_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_7_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28525),
            .in3(N__25600),
            .lcout(\b2v_inst11.mult1_un117_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un117_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25597),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_8_8_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_8_8_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst5.curr_state_7_1_0__m4_0_a2_LC_8_8_0  (
            .in0(N__31494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25576),
            .lcout(N_413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_8_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29251),
            .lcout(\b2v_inst11.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_8_8_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_8_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28830),
            .lcout(\b2v_inst11.mult1_un103_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_8_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35213),
            .lcout(\b2v_inst11.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_8_8_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_8_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28542),
            .lcout(\b2v_inst11.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI4ALGH_5_LC_8_8_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI4ALGH_5_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI4ALGH_5_LC_8_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.count_RNI4ALGH_5_LC_8_8_7  (
            .in0(N__28270),
            .in1(N__32203),
            .in2(N__31762),
            .in3(N__25669),
            .lcout(\b2v_inst5.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_8_9_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_14_LC_8_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_14_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__29705),
            .in2(_gnd_net_),
            .in3(N__25663),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_8_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_10_LC_8_9_1 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_10_LC_8_9_1  (
            .in0(N__26433),
            .in1(N__26206),
            .in2(N__29027),
            .in3(N__29219),
            .lcout(),
            .ltout(\b2v_inst11.i7_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_11_LC_8_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_11_LC_8_9_2 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_11_LC_8_9_2  (
            .in0(N__29128),
            .in1(N__26035),
            .in2(N__25657),
            .in3(N__29000),
            .lcout(\b2v_inst11.dutycycle_RNIZ0Z_11 ),
            .ltout(\b2v_inst11.dutycycle_RNIZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_8_9_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_13_LC_8_9_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_13_LC_8_9_3  (
            .in0(N__29001),
            .in1(_gnd_net_),
            .in2(N__25654),
            .in3(N__28882),
            .lcout(\b2v_inst11.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_8_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_8_LC_8_9_4 .LUT_INIT=16'b1111001010110000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_8_LC_8_9_4  (
            .in0(N__26333),
            .in1(N__25651),
            .in2(N__26843),
            .in3(N__26189),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_12_LC_8_9_5  (
            .in0(N__26434),
            .in1(N__29033),
            .in2(N__25645),
            .in3(N__26334),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_5_10_LC_8_9_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_5_10_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_5_10_LC_8_9_6 .LUT_INIT=16'b0001010100010001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_5_10_LC_8_9_6  (
            .in0(N__29218),
            .in1(N__26432),
            .in2(N__26338),
            .in3(N__26041),
            .lcout(\b2v_inst11.i6_mux_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_8_9_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_13_LC_8_9_7 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_13_LC_8_9_7  (
            .in0(N__29706),
            .in1(N__28881),
            .in2(N__29028),
            .in3(N__26029),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIC6LA7_12_LC_8_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIC6LA7_12_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIC6LA7_12_LC_8_10_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \b2v_inst11.dutycycle_RNIC6LA7_12_LC_8_10_0  (
            .in0(N__25826),
            .in1(N__25989),
            .in2(N__26008),
            .in3(N__26022),
            .lcout(\b2v_inst11.dutycycleZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_12_LC_8_10_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_12_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_12_LC_8_10_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \b2v_inst11.dutycycle_12_LC_8_10_1  (
            .in0(N__26023),
            .in1(N__26004),
            .in2(N__25993),
            .in3(N__25830),
            .lcout(\b2v_inst11.dutycycleZ1Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36614),
            .ce(),
            .sr(N__25947));
    defparam \b2v_inst11.dutycycle_15_LC_8_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_15_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.dutycycle_15_LC_8_10_2 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \b2v_inst11.dutycycle_15_LC_8_10_2  (
            .in0(N__25705),
            .in1(N__25719),
            .in2(N__25857),
            .in3(N__25873),
            .lcout(\b2v_inst11.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36614),
            .ce(),
            .sr(N__25947));
    defparam \b2v_inst11.dutycycle_RNIVV20B_15_LC_8_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIVV20B_15_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIVV20B_15_LC_8_10_3 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \b2v_inst11.dutycycle_RNIVV20B_15_LC_8_10_3  (
            .in0(N__25872),
            .in1(N__25825),
            .in2(N__25723),
            .in3(N__25704),
            .lcout(\b2v_inst11.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_10_LC_8_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_10_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_10_LC_8_10_4 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_10_LC_8_10_4  (
            .in0(N__26280),
            .in1(N__29190),
            .in2(N__26845),
            .in3(N__25693),
            .lcout(),
            .ltout(\b2v_inst11.un1_dutycycle_53_50_1_i_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_8_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_11_LC_8_10_5 .LUT_INIT=16'b0000101100000010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_11_LC_8_10_5  (
            .in0(N__29191),
            .in1(N__26356),
            .in2(N__25681),
            .in3(N__29129),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_4Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_8_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_11_LC_8_10_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_11_LC_8_10_6  (
            .in0(N__29130),
            .in1(N__29594),
            .in2(N__25678),
            .in3(N__29005),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_8_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_10_LC_8_10_7 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_10_LC_8_10_7  (
            .in0(N__29189),
            .in1(N__26437),
            .in2(N__26309),
            .in3(N__26059),
            .lcout(\b2v_inst11.un1_dutycycle_53_50_1_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_8_11_0 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_3_LC_8_11_0 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_3_LC_8_11_0  (
            .in0(N__28775),
            .in1(N__26350),
            .in2(N__28606),
            .in3(N__26167),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_8_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_1_LC_8_11_1 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__29390),
            .in2(N__29535),
            .in3(N__33361),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_1 ),
            .ltout(\b2v_inst11.dutycycle_RNI_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_8_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_0_2_LC_8_11_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_0_2_LC_8_11_2  (
            .in0(N__28774),
            .in1(N__30242),
            .in2(N__26344),
            .in3(N__26166),
            .lcout(\b2v_inst11.dutycycle_RNI_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_3_LC_8_11_3 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_3_LC_8_11_3  (
            .in0(N__29517),
            .in1(N__26835),
            .in2(_gnd_net_),
            .in3(N__28773),
            .lcout(),
            .ltout(\b2v_inst11.dutycycle_RNI_2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_8_11_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_8_LC_8_11_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_8_LC_8_11_4  (
            .in0(N__26276),
            .in1(N__29392),
            .in2(N__26341),
            .in3(N__29518),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_8_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_8_LC_8_11_5 .LUT_INIT=16'b0011001101111111;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_8_LC_8_11_5  (
            .in0(N__26164),
            .in1(N__26275),
            .in2(N__29536),
            .in3(N__26834),
            .lcout(\b2v_inst11.m6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_8_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_2_6_LC_8_11_6 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \b2v_inst11.dutycycle_RNI_2_6_LC_8_11_6  (
            .in0(N__26833),
            .in1(N__29516),
            .in2(_gnd_net_),
            .in3(N__26165),
            .lcout(\b2v_inst11.un1_dutycycle_53_50_1_i_i_a6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_fast_RNIUPHS3_0_LC_8_12_0 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_RNIUPHS3_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_fast_RNIUPHS3_0_LC_8_12_0 .LUT_INIT=16'b1100000011100011;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_RNIUPHS3_0_LC_8_12_0  (
            .in0(N__26482),
            .in1(N__27187),
            .in2(N__27181),
            .in3(N__26854),
            .lcout(N_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_8_12_1 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_12_LC_8_12_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_12_LC_8_12_1  (
            .in0(N__26886),
            .in1(N__27199),
            .in2(_gnd_net_),
            .in3(N__26645),
            .lcout(b2v_inst11_un1_dutycycle_164_0),
            .ltout(b2v_inst11_un1_dutycycle_164_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.RSMRSTn_fast_RNIUPHS3_LC_8_12_2 .C_ON=1'b0;
    defparam \b2v_inst5.RSMRSTn_fast_RNIUPHS3_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.RSMRSTn_fast_RNIUPHS3_LC_8_12_2 .LUT_INIT=16'b1010000010101101;
    LogicCell40 \b2v_inst5.RSMRSTn_fast_RNIUPHS3_LC_8_12_2  (
            .in0(N__27177),
            .in1(N__26481),
            .in2(N__27166),
            .in3(N__26853),
            .lcout(\b2v_inst5.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_8_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_3_LC_8_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_3_LC_8_12_3  (
            .in0(N__28784),
            .in1(N__26837),
            .in2(_gnd_net_),
            .in3(N__29531),
            .lcout(\b2v_inst11.dutycycle_RNI_4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_4_1_LC_8_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_4_1_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_4_1_LC_8_12_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \b2v_inst11.dutycycle_RNI_4_1_LC_8_12_4  (
            .in0(N__26646),
            .in1(N__33629),
            .in2(N__27146),
            .in3(N__33355),
            .lcout(\b2v_inst11.un1_dutycycle_96_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNIVS8U1_2_LC_8_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNIVS8U1_2_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNIVS8U1_2_LC_8_12_6 .LUT_INIT=16'b0000010010101110;
    LogicCell40 \b2v_inst11.dutycycle_RNIVS8U1_2_LC_8_12_6  (
            .in0(N__26962),
            .in1(N__26943),
            .in2(N__26887),
            .in3(N__30241),
            .lcout(N_73_mux_i_i_o3_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_3_LC_8_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_3_LC_8_12_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \b2v_inst11.dutycycle_RNI_3_LC_8_12_7  (
            .in0(N__28785),
            .in1(N__26838),
            .in2(N__26665),
            .in3(N__26644),
            .lcout(g3_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIM92M_12_LC_8_13_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIM92M_12_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIM92M_12_LC_8_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIM92M_12_LC_8_13_0  (
            .in0(N__35922),
            .in1(N__26458),
            .in2(_gnd_net_),
            .in3(N__26466),
            .lcout(\b2v_inst11.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_12_LC_8_13_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_12_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_12_LC_8_13_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_12_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26470),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36632),
            .ce(N__36362),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIMQBN_3_LC_8_13_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIMQBN_3_LC_8_13_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \b2v_inst11.count_RNIMQBN_3_LC_8_13_2  (
            .in0(N__27244),
            .in1(_gnd_net_),
            .in2(N__35934),
            .in3(N__27252),
            .lcout(\b2v_inst11.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_3_LC_8_13_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_3_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_3_LC_8_13_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27256),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36632),
            .ce(N__36362),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOC3M_13_LC_8_13_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOC3M_13_LC_8_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOC3M_13_LC_8_13_4  (
            .in0(N__35923),
            .in1(N__27226),
            .in2(_gnd_net_),
            .in3(N__27234),
            .lcout(\b2v_inst11.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_13_LC_8_13_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_13_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_13_LC_8_13_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_13_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27238),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36632),
            .ce(N__36362),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNIOTCN_4_LC_8_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNIOTCN_4_LC_8_13_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst11.count_RNIOTCN_4_LC_8_13_6  (
            .in0(N__35918),
            .in1(N__27208),
            .in2(_gnd_net_),
            .in3(N__27216),
            .lcout(\b2v_inst11.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_4_LC_8_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_4_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_4_LC_8_13_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \b2v_inst11.count_4_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27220),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36632),
            .ce(N__36362),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNO_0_LC_8_14_0 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNO_0_LC_8_14_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \b2v_inst11.pwm_out_RNO_0_LC_8_14_0  (
            .in0(N__35924),
            .in1(N__29878),
            .in2(_gnd_net_),
            .in3(N__29832),
            .lcout(\b2v_inst11.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_9_LC_8_14_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_9_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_9_LC_8_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst11.count_RNI_9_LC_8_14_1  (
            .in0(N__33119),
            .in1(N__32625),
            .in2(N__32673),
            .in3(N__32718),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_5_LC_8_14_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_5_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_5_LC_8_14_2 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \b2v_inst11.count_RNI_5_LC_8_14_2  (
            .in0(N__32840),
            .in1(N__32894),
            .in2(N__27202),
            .in3(N__27325),
            .lcout(\b2v_inst11.un79_clk_100khzlto15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_2_LC_8_14_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_2_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_2_LC_8_14_3 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.count_RNI_2_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__32939),
            .in2(N__32310),
            .in3(N__32361),
            .lcout(\b2v_inst11.un79_clk_100khzlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_15_LC_8_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_15_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_15_LC_8_14_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst11.count_RNI_15_LC_8_14_4  (
            .in0(N__32811),
            .in1(N__32759),
            .in2(_gnd_net_),
            .in3(N__33017),
            .lcout(),
            .ltout(\b2v_inst11.un79_clk_100khzlto15_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_13_LC_8_14_5 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_13_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_13_LC_8_14_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \b2v_inst11.count_RNI_13_LC_8_14_5  (
            .in0(N__33050),
            .in1(N__33086),
            .in2(N__27319),
            .in3(N__27316),
            .lcout(\b2v_inst11.count_RNIZ0Z_13 ),
            .ltout(\b2v_inst11.count_RNIZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_RNO_1_LC_8_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_RNO_1_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.pwm_out_RNO_1_LC_8_14_6 .LUT_INIT=16'b0011001101111111;
    LogicCell40 \b2v_inst11.pwm_out_RNO_1_LC_8_14_6  (
            .in0(N__35925),
            .in1(N__36408),
            .in2(N__27310),
            .in3(N__29879),
            .lcout(\b2v_inst11.g0_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI03G9_0_LC_8_15_0 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI03G9_0_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI03G9_0_LC_8_15_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst11.count_RNI03G9_0_LC_8_15_0  (
            .in0(N__27292),
            .in1(N__35859),
            .in2(_gnd_net_),
            .in3(N__27370),
            .lcout(\b2v_inst11.countZ0Z_0 ),
            .ltout(\b2v_inst11.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_1_LC_8_15_1 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_1_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_1_LC_8_15_1 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \b2v_inst11.count_RNI_1_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__27420),
            .in2(N__27307),
            .in3(N__32393),
            .lcout(),
            .ltout(\b2v_inst11.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI14G9_1_LC_8_15_2 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI14G9_1_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI14G9_1_LC_8_15_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.count_RNI14G9_1_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__27298),
            .in2(N__27304),
            .in3(N__35860),
            .lcout(\b2v_inst11.countZ0Z_1 ),
            .ltout(\b2v_inst11.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_1_LC_8_15_3 .C_ON=1'b0;
    defparam \b2v_inst11.count_1_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_1_LC_8_15_3 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \b2v_inst11.count_1_LC_8_15_3  (
            .in0(N__32437),
            .in1(_gnd_net_),
            .in2(N__27301),
            .in3(N__27419),
            .lcout(\b2v_inst11.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36645),
            .ce(N__36359),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_0_LC_8_15_4 .C_ON=1'b0;
    defparam \b2v_inst11.count_0_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_0_LC_8_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \b2v_inst11.count_0_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__32436),
            .in2(_gnd_net_),
            .in3(N__27418),
            .lcout(\b2v_inst11.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36645),
            .ce(N__36359),
            .sr(_gnd_net_));
    defparam SLP_S3n_ibuf_RNIHESTE_LC_8_15_5.C_ON=1'b0;
    defparam SLP_S3n_ibuf_RNIHESTE_LC_8_15_5.SEQ_MODE=4'b0000;
    defparam SLP_S3n_ibuf_RNIHESTE_LC_8_15_5.LUT_INIT=16'b0100010000000000;
    LogicCell40 SLP_S3n_ibuf_RNIHESTE_LC_8_15_5 (
            .in0(N__27286),
            .in1(N__27595),
            .in2(_gnd_net_),
            .in3(N__27553),
            .lcout(N_73_mux_i_i_a7_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI0AHN_8_LC_8_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI0AHN_8_LC_8_15_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst11.count_RNI0AHN_8_LC_8_15_6  (
            .in0(N__27511),
            .in1(N__27499),
            .in2(_gnd_net_),
            .in3(N__35861),
            .lcout(\b2v_inst11.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_8_LC_8_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_8_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.count_8_LC_8_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.count_8_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27510),
            .lcout(\b2v_inst11.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36645),
            .ce(N__36359),
            .sr(_gnd_net_));
    defparam \b2v_inst11.pwm_out_LC_8_16_2 .C_ON=1'b0;
    defparam \b2v_inst11.pwm_out_LC_8_16_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst11.pwm_out_LC_8_16_2 .LUT_INIT=16'b1010101011100000;
    LogicCell40 \b2v_inst11.pwm_out_LC_8_16_2  (
            .in0(N__27483),
            .in1(N__32988),
            .in2(N__29883),
            .in3(N__27493),
            .lcout(\b2v_inst11.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36651),
            .ce(),
            .sr(N__27472));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_8_16_4 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_8_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_RNI_LC_8_16_4  (
            .in0(N__29874),
            .in1(N__29837),
            .in2(_gnd_net_),
            .in3(N__32987),
            .lcout(),
            .ltout(\b2v_inst11.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_8_16_5 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIJK34_0_LC_8_16_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst11.curr_state_RNIJK34_0_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(N__29806),
            .in2(N__27463),
            .in3(N__35915),
            .lcout(\b2v_inst11.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst11.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_8_16_6 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.curr_state_RNIOCA3_0_LC_8_16_6 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \b2v_inst11.curr_state_RNIOCA3_0_LC_8_16_6  (
            .in0(N__35916),
            .in1(_gnd_net_),
            .in2(N__27460),
            .in3(N__29836),
            .lcout(\b2v_inst11.count_0_sqmuxa_i ),
            .ltout(\b2v_inst11.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.count_RNI_0_LC_8_16_7 .C_ON=1'b0;
    defparam \b2v_inst11.count_RNI_0_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.count_RNI_0_LC_8_16_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst11.count_RNI_0_LC_8_16_7  (
            .in0(N__32438),
            .in1(_gnd_net_),
            .in2(N__27373),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_c_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(N__27363),
            .in2(N__27352),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_1_THRU_LUT4_0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__30398),
            .in2(_gnd_net_),
            .in3(N__27841),
            .lcout(\b2v_inst36.un2_count_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_1 ),
            .carryout(\b2v_inst36.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_THRU_LUT4_0_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(N__30365),
            .in2(_gnd_net_),
            .in3(N__27838),
            .lcout(\b2v_inst36.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_2 ),
            .carryout(\b2v_inst36.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_3_c_RNICUC8_LC_9_1_3  (
            .in0(N__30978),
            .in1(N__27835),
            .in2(_gnd_net_),
            .in3(N__27808),
            .lcout(\b2v_inst36.count_rst_10 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_3 ),
            .carryout(\b2v_inst36.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_THRU_LUT4_0_LC_9_1_4  (
            .in0(_gnd_net_),
            .in1(N__30321),
            .in2(_gnd_net_),
            .in3(N__27805),
            .lcout(\b2v_inst36.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_4 ),
            .carryout(\b2v_inst36.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_9_1_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_9_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_9_1_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_5_c_RNIE2F8_LC_9_1_5  (
            .in0(N__30979),
            .in1(N__27801),
            .in2(_gnd_net_),
            .in3(N__27775),
            .lcout(\b2v_inst36.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_5 ),
            .carryout(\b2v_inst36.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_6_THRU_LUT4_0_LC_9_1_6  (
            .in0(_gnd_net_),
            .in1(N__31015),
            .in2(_gnd_net_),
            .in3(N__27772),
            .lcout(\b2v_inst36.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_6 ),
            .carryout(\b2v_inst36.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_7_THRU_LUT4_0_LC_9_1_7  (
            .in0(_gnd_net_),
            .in1(N__27902),
            .in2(_gnd_net_),
            .in3(N__27769),
            .lcout(\b2v_inst36.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_7 ),
            .carryout(\b2v_inst36.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_8_c_RNIH8I8_LC_9_2_0  (
            .in0(N__30973),
            .in1(N__27766),
            .in2(_gnd_net_),
            .in3(N__27730),
            .lcout(\b2v_inst36.count_rst_5 ),
            .ltout(),
            .carryin(bfn_9_2_0_),
            .carryout(\b2v_inst36.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_THRU_LUT4_0_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__28142),
            .in2(_gnd_net_),
            .in3(N__27727),
            .lcout(\b2v_inst36.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_9 ),
            .carryout(\b2v_inst36.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_10_THRU_LUT4_0_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(N__28025),
            .in2(_gnd_net_),
            .in3(N__28000),
            .lcout(\b2v_inst36.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_10 ),
            .carryout(\b2v_inst36.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_11_c_RNIR5K1_LC_9_2_3  (
            .in0(N__30950),
            .in1(N__27997),
            .in2(_gnd_net_),
            .in3(N__27958),
            .lcout(\b2v_inst36.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_11 ),
            .carryout(\b2v_inst36.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_12_c_RNIS7L1_LC_9_2_4  (
            .in0(N__30974),
            .in1(N__28107),
            .in2(_gnd_net_),
            .in3(N__27955),
            .lcout(\b2v_inst36.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_12 ),
            .carryout(\b2v_inst36.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNILPEV_LC_9_2_5 .C_ON=1'b1;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNILPEV_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_13_c_RNILPEV_LC_9_2_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_13_c_RNILPEV_LC_9_2_5  (
            .in0(N__30951),
            .in1(N__27948),
            .in2(_gnd_net_),
            .in3(N__27916),
            .lcout(\b2v_inst36.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst36.un2_count_1_cry_13 ),
            .carryout(\b2v_inst36.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_14_c_RNIUBN1_LC_9_2_6  (
            .in0(N__28059),
            .in1(N__30952),
            .in2(_gnd_net_),
            .in3(N__27913),
            .lcout(\b2v_inst36.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_15_LC_9_2_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_15_LC_9_2_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_15_LC_9_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst36.count_15_LC_9_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28071),
            .lcout(\b2v_inst36.count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36659),
            .ce(N__30733),
            .sr(N__30588));
    defparam \b2v_inst36.count_RNIRKI01_8_LC_9_3_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIRKI01_8_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIRKI01_8_LC_9_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst36.count_RNIRKI01_8_LC_9_3_0  (
            .in0(N__27910),
            .in1(N__27856),
            .in2(_gnd_net_),
            .in3(N__30707),
            .lcout(\b2v_inst36.countZ0Z_8 ),
            .ltout(\b2v_inst36.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_8_LC_9_3_1 .C_ON=1'b0;
    defparam \b2v_inst36.count_8_LC_9_3_1 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_8_LC_9_3_1 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst36.count_8_LC_9_3_1  (
            .in0(N__30859),
            .in1(N__27877),
            .in2(N__27859),
            .in3(N__30977),
            .lcout(\b2v_inst36.count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36653),
            .ce(N__30710),
            .sr(N__30580));
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_9_3_2 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_9_3_2 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_9_c_RNIIAJ8_LC_9_3_2  (
            .in0(N__30975),
            .in1(N__28125),
            .in2(N__28149),
            .in3(N__30858),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI6MB61_10_LC_9_3_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI6MB61_10_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI6MB61_10_LC_9_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNI6MB61_10_LC_9_3_3  (
            .in0(N__30708),
            .in1(_gnd_net_),
            .in2(N__28153),
            .in3(N__28114),
            .lcout(\b2v_inst36.countZ0Z_10 ),
            .ltout(\b2v_inst36.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_10_LC_9_3_4 .C_ON=1'b0;
    defparam \b2v_inst36.count_10_LC_9_3_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_10_LC_9_3_4 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \b2v_inst36.count_10_LC_9_3_4  (
            .in0(N__30976),
            .in1(N__28126),
            .in2(N__28117),
            .in3(N__30860),
            .lcout(\b2v_inst36.count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36653),
            .ce(N__30710),
            .sr(N__30580));
    defparam \b2v_inst36.count_RNIJMDV_13_LC_9_3_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIJMDV_13_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIJMDV_13_LC_9_3_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \b2v_inst36.count_RNIJMDV_13_LC_9_3_5  (
            .in0(N__30709),
            .in1(N__28087),
            .in2(_gnd_net_),
            .in3(N__28095),
            .lcout(\b2v_inst36.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_13_LC_9_3_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_13_LC_9_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_13_LC_9_3_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst36.count_13_LC_9_3_6  (
            .in0(N__28096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst36.count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36653),
            .ce(N__30710),
            .sr(N__30580));
    defparam \b2v_inst36.count_RNINSFV_15_LC_9_3_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNINSFV_15_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNINSFV_15_LC_9_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst36.count_RNINSFV_15_LC_9_3_7  (
            .in0(N__28081),
            .in1(N__30711),
            .in2(_gnd_net_),
            .in3(N__28072),
            .lcout(\b2v_inst36.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIL1AS2_0_2_LC_9_4_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL1AS2_0_2_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL1AS2_0_2_LC_9_4_0 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \b2v_inst5.count_RNIL1AS2_0_2_LC_9_4_0  (
            .in0(N__31940),
            .in1(N__28036),
            .in2(N__31219),
            .in3(N__31191),
            .lcout(\b2v_inst5.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIL1AS2_2_LC_9_4_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIL1AS2_2_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIL1AS2_2_LC_9_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIL1AS2_2_LC_9_4_1  (
            .in0(N__28035),
            .in1(N__31873),
            .in2(_gnd_net_),
            .in3(N__31214),
            .lcout(\b2v_inst5.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_2_LC_9_4_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_2_LC_9_4_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_2_LC_9_4_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_2_LC_9_4_2  (
            .in0(N__31215),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36647),
            .ce(N__31939),
            .sr(N__32092));
    defparam \b2v_inst5.count_RNIN4BS2_3_LC_9_4_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIN4BS2_3_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIN4BS2_3_LC_9_4_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \b2v_inst5.count_RNIN4BS2_3_LC_9_4_3  (
            .in0(N__28177),
            .in1(N__32090),
            .in2(N__31177),
            .in3(N__31874),
            .lcout(\b2v_inst5.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI_1_LC_9_4_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI_1_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI_1_LC_9_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst5.count_RNI_1_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(N__31548),
            .in2(_gnd_net_),
            .in3(N__31250),
            .lcout(\b2v_inst5.count_RNIZ0Z_1 ),
            .ltout(\b2v_inst5.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIUHFI2_1_LC_9_4_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIUHFI2_1_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIUHFI2_1_LC_9_4_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \b2v_inst5.count_RNIUHFI2_1_LC_9_4_5  (
            .in0(N__28165),
            .in1(N__31872),
            .in2(N__28180),
            .in3(N__32089),
            .lcout(\b2v_inst5.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_3_LC_9_4_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_3_LC_9_4_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_3_LC_9_4_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \b2v_inst5.count_3_LC_9_4_6  (
            .in0(N__32091),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31176),
            .lcout(\b2v_inst5.count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36647),
            .ce(N__31939),
            .sr(N__32092));
    defparam \b2v_inst5.count_1_LC_9_4_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_1_LC_9_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_1_LC_9_4_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst5.count_1_LC_9_4_7  (
            .in0(_gnd_net_),
            .in1(N__28171),
            .in2(_gnd_net_),
            .in3(N__32093),
            .lcout(\b2v_inst5.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36647),
            .ce(N__31939),
            .sr(N__32092));
    defparam \b2v_inst5.count_RNIJJOV_0_LC_9_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIJJOV_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIJJOV_0_LC_9_5_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst5.count_RNIJJOV_0_LC_9_5_0  (
            .in0(N__31555),
            .in1(N__31517),
            .in2(_gnd_net_),
            .in3(N__32085),
            .lcout(),
            .ltout(\b2v_inst5.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNITGFI2_0_LC_9_5_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNITGFI2_0_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNITGFI2_0_LC_9_5_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.count_RNITGFI2_0_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__31459),
            .in2(N__28159),
            .in3(N__31870),
            .lcout(\b2v_inst5.un2_count_1_cry_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNIRRH21_LC_9_5_2 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNIRRH21_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_c_RNIRRH21_LC_9_5_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_c_RNIRRH21_LC_9_5_2  (
            .in0(N__31386),
            .in1(N__31519),
            .in2(N__31372),
            .in3(N__32087),
            .lcout(\b2v_inst5.count_rst_1 ),
            .ltout(\b2v_inst5.count_rst_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIPDG23_13_LC_9_5_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIPDG23_13_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIPDG23_13_LC_9_5_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.count_RNIPDG23_13_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__28305),
            .in2(N__28156),
            .in3(N__31871),
            .lcout(\b2v_inst5.un2_count_1_axb_13 ),
            .ltout(\b2v_inst5.un2_count_1_axb_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_13_LC_9_5_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_13_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_13_LC_9_5_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst5.count_13_LC_9_5_4  (
            .in0(N__31525),
            .in1(N__32088),
            .in2(N__28318),
            .in3(N__31371),
            .lcout(\b2v_inst5.count_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36640),
            .ce(N__31909),
            .sr(N__32172));
    defparam \b2v_inst5.count_RNIPDG23_0_13_LC_9_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIPDG23_0_13_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIPDG23_0_13_LC_9_5_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \b2v_inst5.count_RNIPDG23_0_13_LC_9_5_5  (
            .in0(N__31251),
            .in1(N__28315),
            .in2(N__28309),
            .in3(N__31910),
            .lcout(\b2v_inst5.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIFEP91_LC_9_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIFEP91_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_c_RNIFEP91_LC_9_5_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_c_RNIFEP91_LC_9_5_6  (
            .in0(N__31059),
            .in1(N__31518),
            .in2(N__31102),
            .in3(N__32086),
            .lcout(\b2v_inst5.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI_15_LC_9_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI_15_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI_15_LC_9_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst5.count_RNI_15_LC_9_5_7  (
            .in0(N__31425),
            .in1(N__31299),
            .in2(N__31345),
            .in3(N__31556),
            .lcout(\b2v_inst5.un12_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__28707),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__28261),
            .in2(N__28386),
            .in3(N__28240),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__28237),
            .in2(N__28387),
            .in3(N__28222),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__32468),
            .in2(N__28219),
            .in3(N__28201),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__28198),
            .in2(N__32475),
            .in3(N__28183),
            .lcout(\b2v_inst11.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5  (
            .in0(N__32497),
            .in1(N__28385),
            .in2(N__28417),
            .in3(N__28399),
            .lcout(\b2v_inst11.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un145_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6  (
            .in0(N__28396),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28390),
            .lcout(\b2v_inst11.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32467),
            .lcout(\b2v_inst11.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_9_7_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_9_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__28543),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_9_7_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__28366),
            .in2(N__28803),
            .in3(N__28351),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_9_7_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__28799),
            .in2(N__28489),
            .in3(N__28342),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_9_7_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__28477),
            .in2(N__28831),
            .in3(N__28330),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_9_7_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__28829),
            .in2(N__28468),
            .in3(N__28321),
            .lcout(\b2v_inst11.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_9_7_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_9_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_9_7_5  (
            .in0(N__31681),
            .in1(N__28456),
            .in2(N__28804),
            .in3(N__28516),
            .lcout(\b2v_inst11.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un110_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_9_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_9_7_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28429),
            .in3(N__28513),
            .lcout(\b2v_inst11.mult1_un110_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un110_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_9_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_9_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28510),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_8_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__29250),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_8_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__35077),
            .in2(N__28446),
            .in3(N__28480),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_8_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__28442),
            .in2(N__34837),
            .in3(N__28471),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_8_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__34810),
            .in2(N__35218),
            .in3(N__28459),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_8_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__35217),
            .in2(N__34786),
            .in3(N__28450),
            .lcout(\b2v_inst11.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_8_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_8_5  (
            .in0(N__28825),
            .in1(N__35269),
            .in2(N__28447),
            .in3(N__28420),
            .lcout(\b2v_inst11.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un103_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_8_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35248),
            .in3(N__28834),
            .lcout(\b2v_inst11.mult1_un103_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un103_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_9_8_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_9_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28807),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_9_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_6_3_LC_9_9_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_6_3_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__28786),
            .in2(N__33634),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_dutycycle_53_axb_0 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_9_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_0_c_RNI5VFB_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__28693),
            .in2(N__33633),
            .in3(N__28660),
            .lcout(\b2v_inst11.mult1_un138_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_0 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_9_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_1_c_RNI61HB_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__30283),
            .in2(N__29272),
            .in3(N__28639),
            .lcout(\b2v_inst11.mult1_un131_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_1 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_9_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_2_c_RNI73IB_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__28636),
            .in2(N__30296),
            .in3(N__28609),
            .lcout(\b2v_inst11.mult1_un124_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_2 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_9_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_3_c_RNI85JB_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__28605),
            .in2(N__28588),
            .in3(N__28561),
            .lcout(\b2v_inst11.mult1_un117_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_3 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_9_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_4_c_RNI97KB_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__29393),
            .in2(N__28558),
            .in3(N__28528),
            .lcout(\b2v_inst11.mult1_un110_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_4 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_9_9_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_5_c_RNIA9LB_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__29260),
            .in2(N__29401),
            .in3(N__29239),
            .lcout(\b2v_inst11.mult1_un103_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_5 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_9_9_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_6_c_RNIBBMB_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__29236),
            .in2(N__29224),
            .in3(N__29134),
            .lcout(\b2v_inst11.mult1_un96_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_6 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_9_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_9_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_7_c_RNICDNB_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__29131),
            .in2(N__29074),
            .in3(N__29059),
            .lcout(\b2v_inst11.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_9_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_8_c_RNIDFOB_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__29056),
            .in2(N__29029),
            .in3(N__28945),
            .lcout(\b2v_inst11.mult1_un82_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_8 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_9_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_9_c_RNIEHPB_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__28897),
            .in2(N__28942),
            .in3(N__28927),
            .lcout(\b2v_inst11.mult1_un75_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_9 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_9_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_10_c_RNIM60B_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__29736),
            .in2(N__28924),
            .in3(N__28915),
            .lcout(\b2v_inst11.mult1_un68_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_10 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_9_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_11_c_RNIN81B_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__29589),
            .in2(N__28912),
            .in3(N__28903),
            .lcout(\b2v_inst11.mult1_un61_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_11 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_9_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_9_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_12_c_RNIOA2B_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__28898),
            .in2(N__28846),
            .in3(N__28837),
            .lcout(\b2v_inst11.mult1_un54_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_12 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_9_10_6 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_9_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_13_c_RNIPC3B_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__29732),
            .in2(N__29659),
            .in3(N__29650),
            .lcout(\b2v_inst11.mult1_un47_sum ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_13 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_9_10_7 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_9_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__29590),
            .in2(N__29647),
            .in3(N__29629),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4BZ0 ),
            .ltout(),
            .carryin(\b2v_inst11.un1_dutycycle_53_cry_14 ),
            .carryout(\b2v_inst11.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_9_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_9_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5B_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(N__29626),
            .in2(N__29607),
            .in3(N__29545),
            .lcout(\b2v_inst11.un1_dutycycle_53_cry_15_c_RNIRG5BZ0 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\b2v_inst11.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_9_11_1 .C_ON=1'b0;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.CO2_THRU_LUT4_0_LC_9_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.CO2_THRU_LUT4_0_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29542),
            .lcout(\b2v_inst11.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_11_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_11_2 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29923),
            .in3(N__29774),
            .lcout(\b2v_inst11.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_11_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30024),
            .lcout(\b2v_inst11.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.dutycycle_RNI_1_1_LC_9_11_5 .C_ON=1'b0;
    defparam \b2v_inst11.dutycycle_RNI_1_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.dutycycle_RNI_1_1_LC_9_11_5 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \b2v_inst11.dutycycle_RNI_1_1_LC_9_11_5  (
            .in0(N__29524),
            .in1(N__29391),
            .in2(N__30297),
            .in3(N__33362),
            .lcout(\b2v_inst11.dutycycle_RNI_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_7 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__29920),
            .in2(N__29779),
            .in3(N__29793),
            .lcout(\b2v_inst11.mult1_un40_sum_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.curr_state_0_LC_9_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.curr_state_0_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst11.curr_state_0_LC_9_12_0 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \b2v_inst11.curr_state_0_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__32983),
            .in2(N__29887),
            .in3(N__29839),
            .lcout(\b2v_inst11.curr_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36633),
            .ce(N__36365),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_12_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_12_2 .LUT_INIT=16'b1111000011000011;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__29922),
            .in2(N__29794),
            .in3(N__29778),
            .lcout(\b2v_inst11.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_12_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30054),
            .in3(N__29938),
            .lcout(\b2v_inst11.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_12_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_12_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_12_5  (
            .in0(N__30086),
            .in1(N__30087),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33261),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29761),
            .in3(N__29749),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__30034),
            .in2(N__30010),
            .in3(N__29746),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__30437),
            .in2(N__29977),
            .in3(N__29743),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__30438),
            .in2(N__29953),
            .in3(N__29740),
            .lcout(\b2v_inst11.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_13_5  (
            .in0(N__36187),
            .in1(N__30088),
            .in2(N__30070),
            .in3(N__30061),
            .lcout(\b2v_inst11.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un54_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_13_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__29937),
            .in2(N__30058),
            .in3(N__30037),
            .lcout(\b2v_inst11.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_13_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_13_7  (
            .in0(N__30005),
            .in1(N__30006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_14_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30028),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_14_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29896),
            .in3(N__29992),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_14_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29989),
            .in3(N__29968),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_14_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__30436),
            .in2(N__29965),
            .in3(N__29944),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un47_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_9_14_4 .C_ON=1'b0;
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_9_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29941),
            .lcout(\b2v_inst11.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_9_14_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_9_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_dutycycle_53_cry_14_c_RNIQE4B_0_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29921),
            .lcout(\b2v_inst11.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_9_14_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_9_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_9_14_7  (
            .in0(N__30291),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_9_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_9_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__33363),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__30190),
            .in2(N__30488),
            .in3(N__30184),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__30181),
            .in2(N__30490),
            .in3(N__30169),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__30166),
            .in2(N__31747),
            .in3(N__30148),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__30145),
            .in2(N__31746),
            .in3(N__30127),
            .lcout(\b2v_inst11.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_15_5  (
            .in0(N__33954),
            .in1(N__30124),
            .in2(N__30489),
            .in3(N__30106),
            .lcout(\b2v_inst11.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un159_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_15_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__30103),
            .in2(_gnd_net_),
            .in3(N__30091),
            .lcout(\b2v_inst11.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_15_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31739),
            .lcout(\b2v_inst11.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.curr_state_1_LC_9_16_0 .C_ON=1'b0;
    defparam \b2v_inst5.curr_state_1_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \b2v_inst5.curr_state_1_LC_9_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst5.curr_state_1_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30466),
            .lcout(\b2v_inst5.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36658),
            .ce(N__36360),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_16_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_16_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_16_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNI_2_LC_11_1_0 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNI_2_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNI_2_LC_11_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst36.count_RNI_2_LC_11_1_0  (
            .in0(N__30366),
            .in1(N__31013),
            .in2(N__30325),
            .in3(N__30406),
            .lcout(\b2v_inst36.un12_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_11_1_1 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_11_1_1 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_2_c_RNIBSB8_LC_11_1_1  (
            .in0(N__30348),
            .in1(N__30981),
            .in2(N__30861),
            .in3(N__30367),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNIH5D01_3_LC_11_1_2 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNIH5D01_3_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNIH5D01_3_LC_11_1_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst36.count_RNIH5D01_3_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(N__30334),
            .in2(N__30370),
            .in3(N__30725),
            .lcout(\b2v_inst36.countZ0Z_3 ),
            .ltout(\b2v_inst36.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_3_LC_11_1_3 .C_ON=1'b0;
    defparam \b2v_inst36.count_3_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_3_LC_11_1_3 .LUT_INIT=16'b0000000001001000;
    LogicCell40 \b2v_inst36.count_3_LC_11_1_3  (
            .in0(N__30349),
            .in1(N__30985),
            .in2(N__30337),
            .in3(N__30854),
            .lcout(\b2v_inst36.count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36664),
            .ce(N__30731),
            .sr(N__30589));
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_11_1_4 .C_ON=1'b0;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_11_1_4 .LUT_INIT=16'b0001000001000000;
    LogicCell40 \b2v_inst36.un2_count_1_cry_4_c_RNID0E8_LC_11_1_4  (
            .in0(N__30852),
            .in1(N__31038),
            .in2(N__30988),
            .in3(N__30320),
            .lcout(),
            .ltout(\b2v_inst36.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_RNILBF01_5_LC_11_1_5 .C_ON=1'b0;
    defparam \b2v_inst36.count_RNILBF01_5_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst36.count_RNILBF01_5_LC_11_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst36.count_RNILBF01_5_LC_11_1_5  (
            .in0(N__30726),
            .in1(_gnd_net_),
            .in2(N__30328),
            .in3(N__31021),
            .lcout(\b2v_inst36.countZ0Z_5 ),
            .ltout(\b2v_inst36.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst36.count_5_LC_11_1_6 .C_ON=1'b0;
    defparam \b2v_inst36.count_5_LC_11_1_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_5_LC_11_1_6 .LUT_INIT=16'b0001010000000000;
    LogicCell40 \b2v_inst36.count_5_LC_11_1_6  (
            .in0(N__30853),
            .in1(N__31039),
            .in2(N__31024),
            .in3(N__30987),
            .lcout(\b2v_inst36.count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36664),
            .ce(N__30731),
            .sr(N__30589));
    defparam \b2v_inst36.count_7_LC_11_1_7 .C_ON=1'b0;
    defparam \b2v_inst36.count_7_LC_11_1_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst36.count_7_LC_11_1_7 .LUT_INIT=16'b0000010000001000;
    LogicCell40 \b2v_inst36.count_7_LC_11_1_7  (
            .in0(N__31014),
            .in1(N__30986),
            .in2(N__30862),
            .in3(N__30766),
            .lcout(\b2v_inst36.count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36664),
            .ce(N__30731),
            .sr(N__30589));
    defparam \b2v_inst6.count_14_LC_11_2_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_14_LC_11_2_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_14_LC_11_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_14_LC_11_2_0  (
            .in0(N__33991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36662),
            .ce(N__35058),
            .sr(N__36129));
    defparam \b2v_inst6.count_RNIPG489_14_LC_11_2_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIPG489_14_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIPG489_14_LC_11_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIPG489_14_LC_11_2_1  (
            .in0(N__30505),
            .in1(N__33990),
            .in2(_gnd_net_),
            .in3(N__35040),
            .lcout(\b2v_inst6.countZ0Z_14 ),
            .ltout(\b2v_inst6.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_2_LC_11_2_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_2_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_2_LC_11_2_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \b2v_inst6.count_RNI_2_LC_11_2_2  (
            .in0(N__34147),
            .in1(N__34044),
            .in2(N__30499),
            .in3(N__33871),
            .lcout(\b2v_inst6.count_1_i_a3_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_13_LC_11_2_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_13_LC_11_2_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_13_LC_11_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_13_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34159),
            .lcout(\b2v_inst6.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36662),
            .ce(N__35058),
            .sr(N__36129));
    defparam \b2v_inst6.count_RNIRB4V8_6_LC_11_2_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRB4V8_6_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRB4V8_6_LC_11_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst6.count_RNIRB4V8_6_LC_11_2_5  (
            .in0(N__34029),
            .in1(N__30496),
            .in2(_gnd_net_),
            .in3(N__35039),
            .lcout(\b2v_inst6.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_6_LC_11_2_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_6_LC_11_2_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_6_LC_11_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_6_LC_11_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34030),
            .lcout(\b2v_inst6.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36662),
            .ce(N__35058),
            .sr(N__36129));
    defparam \b2v_inst6.count_RNIJVVU8_2_LC_11_2_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIJVVU8_2_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIJVVU8_2_LC_11_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIJVVU8_2_LC_11_2_7  (
            .in0(N__34351),
            .in1(N__34362),
            .in2(_gnd_net_),
            .in3(N__35038),
            .lcout(\b2v_inst6.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_1_c_LC_11_3_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_1_c_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_1_c_LC_11_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_1_c_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__31255),
            .in2(N__31564),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNI92J91_LC_11_3_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNI92J91_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_1_c_RNI92J91_LC_11_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_1_c_RNI92J91_LC_11_3_1  (
            .in0(N__32175),
            .in1(N__31231),
            .in2(_gnd_net_),
            .in3(N__31198),
            .lcout(\b2v_inst5.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_1 ),
            .carryout(\b2v_inst5.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_3_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \b2v_inst5.un2_count_1_cry_2_c_RNINGR9_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__31195),
            .in2(_gnd_net_),
            .in3(N__31159),
            .lcout(\b2v_inst5.un2_count_1_cry_2_c_RNINGRZ0Z9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_2 ),
            .carryout(\b2v_inst5.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_3_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_3_THRU_LUT4_0_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__31156),
            .in2(_gnd_net_),
            .in3(N__31114),
            .lcout(\b2v_inst5.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_3 ),
            .carryout(\b2v_inst5.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIC8M91_LC_11_3_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIC8M91_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_4_c_RNIC8M91_LC_11_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_4_c_RNIC8M91_LC_11_3_4  (
            .in0(N__32177),
            .in1(N__32269),
            .in2(_gnd_net_),
            .in3(N__31111),
            .lcout(\b2v_inst5.count_rst_9 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_4 ),
            .carryout(\b2v_inst5.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIDAN91_LC_11_3_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIDAN91_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_5_c_RNIDAN91_LC_11_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_5_c_RNIDAN91_LC_11_3_5  (
            .in0(N__32176),
            .in1(N__32242),
            .in2(_gnd_net_),
            .in3(N__31108),
            .lcout(\b2v_inst5.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_5 ),
            .carryout(\b2v_inst5.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIECO91_LC_11_3_6 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIECO91_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_6_c_RNIECO91_LC_11_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_6_c_RNIECO91_LC_11_3_6  (
            .in0(N__32178),
            .in1(N__32191),
            .in2(_gnd_net_),
            .in3(N__31105),
            .lcout(\b2v_inst5.count_rst_7 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_6 ),
            .carryout(\b2v_inst5.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_7 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(N__31101),
            .in2(_gnd_net_),
            .in3(N__31042),
            .lcout(\b2v_inst5.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_7 ),
            .carryout(\b2v_inst5.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_4_0 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_THRU_LUT4_0_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__31659),
            .in2(_gnd_net_),
            .in3(N__31450),
            .lcout(\b2v_inst5.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\b2v_inst5.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_4_1 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_THRU_LUT4_0_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__31599),
            .in2(_gnd_net_),
            .in3(N__31447),
            .lcout(\b2v_inst5.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_9 ),
            .carryout(\b2v_inst5.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNIPNF21_LC_11_4_2 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNIPNF21_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_10_c_RNIPNF21_LC_11_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_10_c_RNIPNF21_LC_11_4_2  (
            .in0(N__32179),
            .in1(N__31956),
            .in2(_gnd_net_),
            .in3(N__31429),
            .lcout(\b2v_inst5.count_rst_3 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_10 ),
            .carryout(\b2v_inst5.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNIQPG21_LC_11_4_3 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNIQPG21_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_11_c_RNIQPG21_LC_11_4_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_11_c_RNIQPG21_LC_11_4_3  (
            .in0(N__32180),
            .in1(N__31426),
            .in2(_gnd_net_),
            .in3(N__31393),
            .lcout(\b2v_inst5.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_11 ),
            .carryout(\b2v_inst5.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_4_4 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.un2_count_1_cry_12_THRU_LUT4_0_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__31390),
            .in2(_gnd_net_),
            .in3(N__31348),
            .lcout(\b2v_inst5.un2_count_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_12 ),
            .carryout(\b2v_inst5.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNISTI21_LC_11_4_5 .C_ON=1'b1;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNISTI21_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_13_c_RNISTI21_LC_11_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst5.un2_count_1_cry_13_c_RNISTI21_LC_11_4_5  (
            .in0(N__32181),
            .in1(N__31341),
            .in2(_gnd_net_),
            .in3(N__31306),
            .lcout(\b2v_inst5.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst5.un2_count_1_cry_13 ),
            .carryout(\b2v_inst5.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNITVJ21_LC_11_4_6 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNITVJ21_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_14_c_RNITVJ21_LC_11_4_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_14_c_RNITVJ21_LC_11_4_6  (
            .in0(N__31303),
            .in1(N__32182),
            .in2(_gnd_net_),
            .in3(N__31288),
            .lcout(\b2v_inst5.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_15_LC_11_4_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_15_LC_11_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_15_LC_11_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst5.count_15_LC_11_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31278),
            .lcout(\b2v_inst5.count_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36655),
            .ce(N__31927),
            .sr(N__32174));
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNIGGQ91_LC_11_5_0 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNIGGQ91_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_8_c_RNIGGQ91_LC_11_5_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_8_c_RNIGGQ91_LC_11_5_0  (
            .in0(N__31660),
            .in1(N__31520),
            .in2(N__31648),
            .in3(N__32140),
            .lcout(\b2v_inst5.count_rst_5 ),
            .ltout(\b2v_inst5.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNI3NHS2_9_LC_11_5_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI3NHS2_9_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI3NHS2_9_LC_11_5_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \b2v_inst5.count_RNI3NHS2_9_LC_11_5_1  (
            .in0(N__31633),
            .in1(_gnd_net_),
            .in2(N__31663),
            .in3(N__31882),
            .lcout(\b2v_inst5.un2_count_1_axb_9 ),
            .ltout(\b2v_inst5.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_9_LC_11_5_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_9_LC_11_5_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_9_LC_11_5_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_9_LC_11_5_2  (
            .in0(N__31647),
            .in1(N__31522),
            .in2(N__31636),
            .in3(N__32143),
            .lcout(\b2v_inst5.count_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36648),
            .ce(N__31883),
            .sr(N__32170));
    defparam \b2v_inst5.count_RNI3NHS2_0_9_LC_11_5_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNI3NHS2_0_9_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNI3NHS2_0_9_LC_11_5_3 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \b2v_inst5.count_RNI3NHS2_0_9_LC_11_5_3  (
            .in0(N__31632),
            .in1(N__31881),
            .in2(N__31624),
            .in3(N__31595),
            .lcout(\b2v_inst5.un12_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNIHIR91_LC_11_5_4 .C_ON=1'b0;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNIHIR91_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un2_count_1_cry_9_c_RNIHIR91_LC_11_5_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.un2_count_1_cry_9_c_RNIHIR91_LC_11_5_4  (
            .in0(N__31582),
            .in1(N__31523),
            .in2(N__31600),
            .in3(N__32139),
            .lcout(),
            .ltout(\b2v_inst5.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIC1Q93_10_LC_11_5_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIC1Q93_10_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIC1Q93_10_LC_11_5_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst5.count_RNIC1Q93_10_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__31570),
            .in2(N__31603),
            .in3(N__31880),
            .lcout(\b2v_inst5.countZ0Z_10 ),
            .ltout(\b2v_inst5.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_10_LC_11_5_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_10_LC_11_5_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_10_LC_11_5_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst5.count_10_LC_11_5_6  (
            .in0(N__31581),
            .in1(N__31521),
            .in2(N__31573),
            .in3(N__32142),
            .lcout(\b2v_inst5.count_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36648),
            .ce(N__31883),
            .sr(N__32170));
    defparam \b2v_inst5.count_0_LC_11_5_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_0_LC_11_5_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_0_LC_11_5_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \b2v_inst5.count_0_LC_11_5_7  (
            .in0(N__32141),
            .in1(N__31560),
            .in2(_gnd_net_),
            .in3(N__31524),
            .lcout(\b2v_inst5.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36648),
            .ce(N__31883),
            .sr(N__32170));
    defparam \b2v_inst5.count_6_LC_11_6_0 .C_ON=1'b0;
    defparam \b2v_inst5.count_6_LC_11_6_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_6_LC_11_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_6_LC_11_6_0  (
            .in0(N__32254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36641),
            .ce(N__31907),
            .sr(N__32171));
    defparam \b2v_inst5.count_RNIRADS2_5_LC_11_6_1 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRADS2_5_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRADS2_5_LC_11_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIRADS2_5_LC_11_6_1  (
            .in0(N__32211),
            .in1(N__31884),
            .in2(_gnd_net_),
            .in3(N__32231),
            .lcout(\b2v_inst5.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_5_LC_11_6_2 .C_ON=1'b0;
    defparam \b2v_inst5.count_5_LC_11_6_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_5_LC_11_6_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_5_LC_11_6_2  (
            .in0(N__32232),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36641),
            .ce(N__31907),
            .sr(N__32171));
    defparam \b2v_inst5.count_RNITDES2_6_LC_11_6_3 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNITDES2_6_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNITDES2_6_LC_11_6_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNITDES2_6_LC_11_6_3  (
            .in0(N__32260),
            .in1(N__31885),
            .in2(_gnd_net_),
            .in3(N__32253),
            .lcout(\b2v_inst5.countZ0Z_6 ),
            .ltout(\b2v_inst5.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIRADS2_0_5_LC_11_6_4 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIRADS2_0_5_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIRADS2_0_5_LC_11_6_4 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \b2v_inst5.count_RNIRADS2_0_5_LC_11_6_4  (
            .in0(N__31887),
            .in1(N__32233),
            .in2(N__32215),
            .in3(N__32212),
            .lcout(\b2v_inst5.un12_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_RNIVGFS2_7_LC_11_6_5 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIVGFS2_7_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIVGFS2_7_LC_11_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst5.count_RNIVGFS2_7_LC_11_6_5  (
            .in0(N__31986),
            .in1(N__31886),
            .in2(_gnd_net_),
            .in3(N__31976),
            .lcout(\b2v_inst5.un2_count_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.count_7_LC_11_6_6 .C_ON=1'b0;
    defparam \b2v_inst5.count_7_LC_11_6_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst5.count_7_LC_11_6_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst5.count_7_LC_11_6_6  (
            .in0(N__31977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst5.count_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36641),
            .ce(N__31907),
            .sr(N__32171));
    defparam \b2v_inst5.count_RNIVGFS2_0_7_LC_11_6_7 .C_ON=1'b0;
    defparam \b2v_inst5.count_RNIVGFS2_0_7_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.count_RNIVGFS2_0_7_LC_11_6_7 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \b2v_inst5.count_RNIVGFS2_0_7_LC_11_6_7  (
            .in0(N__31987),
            .in1(N__31978),
            .in2(N__31963),
            .in3(N__31908),
            .lcout(\b2v_inst5.un12_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_7_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31730),
            .lcout(\b2v_inst11.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_11_7_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_11_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31690),
            .lcout(\b2v_inst11.mult1_un110_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_11_7_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_11_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32587),
            .lcout(\b2v_inst11.mult1_un117_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_7_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32560),
            .lcout(\b2v_inst11.mult1_un124_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_11_7_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_11_7_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_11_7_6  (
            .in0(N__32521),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un145_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_7_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32479),
            .lcout(\b2v_inst11.mult1_un138_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_11_8_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_11_8_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_0_c_inv_LC_11_8_0  (
            .in0(N__32446),
            .in1(N__32410),
            .in2(N__33889),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_11_8_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_11_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_1_c_inv_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__32374),
            .in2(N__33190),
            .in3(N__32404),
            .lcout(\b2v_inst11.N_5530_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_0 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_11_8_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_11_8_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_2_c_inv_LC_11_8_2  (
            .in0(N__32368),
            .in1(N__32323),
            .in2(N__32332),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5531_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_1 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_11_8_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_11_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_3_c_inv_LC_11_8_3  (
            .in0(N__32317),
            .in1(N__32275),
            .in2(N__32287),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5532_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_2 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_11_8_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_11_8_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_4_c_inv_LC_11_8_4  (
            .in0(N__32950),
            .in1(N__32914),
            .in2(N__32923),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5533_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_3 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_11_8_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_11_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_5_c_inv_LC_11_8_5  (
            .in0(N__32908),
            .in1(N__32866),
            .in2(N__32881),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5534_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_4 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_11_8_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_11_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_6_c_inv_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__32824),
            .in2(N__32860),
            .in3(N__32851),
            .lcout(\b2v_inst11.N_5535_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_5 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_11_8_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_11_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_7_c_inv_LC_11_8_7  (
            .in0(N__32818),
            .in1(N__32776),
            .in2(N__32785),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5536_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_6 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_11_9_0 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_11_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_8_c_inv_LC_11_9_0  (
            .in0(N__32770),
            .in1(N__32743),
            .in2(N__32734),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5537_i ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_11_9_1 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_11_9_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_9_c_inv_LC_11_9_1  (
            .in0(N__32725),
            .in1(N__32680),
            .in2(N__32695),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5538_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_8 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_11_9_2 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_11_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_10_c_inv_LC_11_9_2  (
            .in0(N__32674),
            .in1(N__34546),
            .in2(N__32638),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5539_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_9 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_11_9_3 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_11_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_11_c_inv_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__33196),
            .in2(N__32596),
            .in3(N__32629),
            .lcout(\b2v_inst11.N_5540_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_10 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_11_9_4 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_11_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_12_c_inv_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__33175),
            .in2(N__33103),
            .in3(N__33127),
            .lcout(\b2v_inst11.N_5541_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_11 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_11_9_5 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_11_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_13_c_inv_LC_11_9_5  (
            .in0(N__33094),
            .in1(N__34552),
            .in2(N__33070),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5542_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_12 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_11_9_6 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_11_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_14_c_inv_LC_11_9_6  (
            .in0(N__33061),
            .in1(N__35065),
            .in2(N__33034),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5543_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_13 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_11_9_7 .C_ON=1'b1;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_11_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_c_inv_LC_11_9_7  (
            .in0(N__33025),
            .in1(N__33238),
            .in2(N__33001),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.N_5544_i ),
            .ltout(),
            .carryin(\b2v_inst11.un85_clk_100khz_cry_14 ),
            .carryout(\b2v_inst11.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_11_10_0 .C_ON=1'b0;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32992),
            .lcout(\b2v_inst11.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_10_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33168),
            .lcout(\b2v_inst11.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_11_10_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_11_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35337),
            .lcout(\b2v_inst11.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_10_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35136),
            .lcout(\b2v_inst11.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_11_10_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_11_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35181),
            .lcout(\b2v_inst11.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33970),
            .lcout(\b2v_inst11.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_11_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_11_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35382),
            .lcout(\b2v_inst11.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__33169),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__33148),
            .in2(N__35355),
            .in3(N__33142),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__35351),
            .in2(N__35110),
            .in3(N__33139),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__35098),
            .in2(N__35383),
            .in3(N__33136),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__35381),
            .in2(N__35089),
            .in3(N__33133),
            .lcout(\b2v_inst11.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_11_5  (
            .in0(N__35180),
            .in1(N__35410),
            .in2(N__35356),
            .in3(N__33130),
            .lcout(\b2v_inst11.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un89_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35398),
            .in3(N__33367),
            .lcout(\b2v_inst11.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_11_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_11_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36230),
            .lcout(\b2v_inst11.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_11_12_0 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_11_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33364),
            .lcout(\b2v_inst11.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_11_12_3 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_11_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33262),
            .lcout(\b2v_inst11.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_11_12_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_11_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33229),
            .lcout(\b2v_inst11.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_11_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_11_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35527),
            .lcout(\b2v_inst11.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_11_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_11_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35448),
            .lcout(\b2v_inst11.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__33228),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__33205),
            .in2(N__36165),
            .in3(N__33199),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__36161),
            .in2(N__33499),
            .in3(N__33484),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__33481),
            .in2(N__36196),
            .in3(N__33472),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__36194),
            .in2(N__33469),
            .in3(N__33457),
            .lcout(\b2v_inst11.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_13_5  (
            .in0(N__35443),
            .in1(N__33454),
            .in2(N__36166),
            .in3(N__33445),
            .lcout(\b2v_inst11.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un61_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33442),
            .in3(N__33430),
            .lcout(\b2v_inst11.mult1_un61_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un61_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33427),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_14_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_14_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_i_o3_0_LC_11_14_0  (
            .in0(N__35654),
            .in1(N__36148),
            .in2(_gnd_net_),
            .in3(N__36819),
            .lcout(\b2v_inst6.N_241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst31.un6_output_LC_11_14_1 .C_ON=1'b0;
    defparam \b2v_inst31.un6_output_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst31.un6_output_LC_11_14_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \b2v_inst31.un6_output_LC_11_14_1  (
            .in0(N__34711),
            .in1(N__33424),
            .in2(N__33802),
            .in3(N__33412),
            .lcout(VCCIN_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIUL1J2_0_0_LC_11_14_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIUL1J2_0_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIUL1J2_0_0_LC_11_14_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIUL1J2_0_0_LC_11_14_2  (
            .in0(N__35652),
            .in1(N__36147),
            .in2(_gnd_net_),
            .in3(N__36817),
            .lcout(\b2v_inst6.N_276_0 ),
            .ltout(\b2v_inst6.N_276_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_14_3 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_14_3 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_LC_11_14_3  (
            .in0(N__36402),
            .in1(N__33820),
            .in2(N__33847),
            .in3(N__35632),
            .lcout(\b2v_inst6.delayed_vccin_vccinaux_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36654),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_11_14_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_11_14_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \b2v_inst6.count_0_sqmuxa_0_o2_4_LC_11_14_4  (
            .in0(N__33844),
            .in1(N__33832),
            .in2(_gnd_net_),
            .in3(N__33796),
            .lcout(\b2v_inst6.N_192 ),
            .ltout(\b2v_inst6.N_192_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIUL1J2_0_LC_11_14_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIUL1J2_0_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIUL1J2_0_LC_11_14_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIUL1J2_0_LC_11_14_5  (
            .in0(N__36818),
            .in1(_gnd_net_),
            .in2(N__33823),
            .in3(N__35653),
            .lcout(\b2v_inst6.curr_state_RNIUL1J2Z0Z_0 ),
            .ltout(\b2v_inst6.curr_state_RNIUL1J2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU0GV5_LC_11_14_6 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU0GV5_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU0GV5_LC_11_14_6 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNIU0GV5_LC_11_14_6  (
            .in0(N__33819),
            .in1(N__36401),
            .in2(N__33811),
            .in3(N__33808),
            .lcout(),
            .ltout(\b2v_inst6.delayed_vccin_vccinaux_okZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_LC_11_14_7 .C_ON=1'b0;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_LC_11_14_7 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \b2v_inst6.delayed_vccin_vccinaux_ok_RNI8L1J7_LC_11_14_7  (
            .in0(N__33797),
            .in1(_gnd_net_),
            .in2(N__33691),
            .in3(_gnd_net_),
            .lcout(N_222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_11_15_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_11_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__33628),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_11_15_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_11_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__33529),
            .in2(N__33918),
            .in3(N__33955),
            .lcout(G_2836),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_0 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_11_15_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_11_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__33914),
            .in2(N__33520),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_1 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_11_15_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_11_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__33508),
            .in2(N__33966),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_11_15_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_11_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__33979),
            .in2(N__33965),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_11_15_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_11_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__33928),
            .in2(N__33919),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un166_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_11_15_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_11_15_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_11_15_6  (
            .in0(N__33901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33892),
            .lcout(\b2v_inst11.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_12_1_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_LC_12_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_LC_12_1_0  (
            .in0(_gnd_net_),
            .in1(N__34900),
            .in2(N__34459),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_1_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNID55Q2_LC_12_1_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNID55Q2_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_1_c_RNID55Q2_LC_12_1_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_1_c_RNID55Q2_LC_12_1_1  (
            .in0(N__36112),
            .in1(N__33870),
            .in2(_gnd_net_),
            .in3(N__33859),
            .lcout(\b2v_inst6.count_rst_12 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_1 ),
            .carryout(\b2v_inst6.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_12_1_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_12_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_THRU_LUT4_0_LC_12_1_2  (
            .in0(_gnd_net_),
            .in1(N__34535),
            .in2(_gnd_net_),
            .in3(N__33856),
            .lcout(\b2v_inst6.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_2 ),
            .carryout(\b2v_inst6.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_12_1_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_12_1_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_12_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_THRU_LUT4_0_LC_12_1_3  (
            .in0(_gnd_net_),
            .in1(N__34227),
            .in2(_gnd_net_),
            .in3(N__33853),
            .lcout(\b2v_inst6.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_3 ),
            .carryout(\b2v_inst6.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_12_1_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_12_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_THRU_LUT4_0_LC_12_1_4  (
            .in0(_gnd_net_),
            .in1(N__34096),
            .in2(_gnd_net_),
            .in3(N__33850),
            .lcout(\b2v_inst6.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_4 ),
            .carryout(\b2v_inst6.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIHD9Q2_LC_12_1_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIHD9Q2_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_5_c_RNIHD9Q2_LC_12_1_5 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_5_c_RNIHD9Q2_LC_12_1_5  (
            .in0(N__36113),
            .in1(_gnd_net_),
            .in2(N__34045),
            .in3(N__34021),
            .lcout(\b2v_inst6.count_rst_8 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_5 ),
            .carryout(\b2v_inst6.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_12_1_6 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_12_1_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_12_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_THRU_LUT4_0_LC_12_1_6  (
            .in0(_gnd_net_),
            .in1(N__34409),
            .in2(_gnd_net_),
            .in3(N__34018),
            .lcout(\b2v_inst6.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_6 ),
            .carryout(\b2v_inst6.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_12_1_7 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_12_1_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_12_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_THRU_LUT4_0_LC_12_1_7  (
            .in0(_gnd_net_),
            .in1(N__34333),
            .in2(_gnd_net_),
            .in3(N__34015),
            .lcout(\b2v_inst6.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_7 ),
            .carryout(\b2v_inst6.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_12_2_0 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_12_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_THRU_LUT4_0_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__34073),
            .in2(_gnd_net_),
            .in3(N__34012),
            .lcout(\b2v_inst6.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\b2v_inst6.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNILLDQ2_LC_12_2_1 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNILLDQ2_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_9_c_RNILLDQ2_LC_12_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_9_c_RNILLDQ2_LC_12_2_1  (
            .in0(N__36085),
            .in1(N__34279),
            .in2(_gnd_net_),
            .in3(N__34009),
            .lcout(\b2v_inst6.count_rst_4 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_9 ),
            .carryout(\b2v_inst6.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_12_2_2 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_12_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_THRU_LUT4_0_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__34626),
            .in2(_gnd_net_),
            .in3(N__34006),
            .lcout(\b2v_inst6.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_10 ),
            .carryout(\b2v_inst6.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIUTM13_LC_12_2_3 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIUTM13_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_11_c_RNIUTM13_LC_12_2_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \b2v_inst6.un2_count_1_cry_11_c_RNIUTM13_LC_12_2_3  (
            .in0(N__36086),
            .in1(_gnd_net_),
            .in2(N__34249),
            .in3(N__34003),
            .lcout(\b2v_inst6.count_rst_2 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_11 ),
            .carryout(\b2v_inst6.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNIVVN13_LC_12_2_4 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNIVVN13_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_12_c_RNIVVN13_LC_12_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_12_c_RNIVVN13_LC_12_2_4  (
            .in0(N__36088),
            .in1(N__34143),
            .in2(_gnd_net_),
            .in3(N__34000),
            .lcout(\b2v_inst6.count_rst_1 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_12 ),
            .carryout(\b2v_inst6.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI02P13_LC_12_2_5 .C_ON=1'b1;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI02P13_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_13_c_RNI02P13_LC_12_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_13_c_RNI02P13_LC_12_2_5  (
            .in0(N__36087),
            .in1(N__33997),
            .in2(_gnd_net_),
            .in3(N__33982),
            .lcout(\b2v_inst6.count_rst_0 ),
            .ltout(),
            .carryin(\b2v_inst6.un2_count_1_cry_13 ),
            .carryout(\b2v_inst6.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNI14Q13_LC_12_2_6 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNI14Q13_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_14_c_RNI14Q13_LC_12_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \b2v_inst6.un2_count_1_cry_14_c_RNI14Q13_LC_12_2_6  (
            .in0(N__36089),
            .in1(N__34651),
            .in2(_gnd_net_),
            .in3(N__34171),
            .lcout(\b2v_inst6.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIND389_13_LC_12_2_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIND389_13_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIND389_13_LC_12_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIND389_13_LC_12_2_7  (
            .in0(N__34168),
            .in1(N__34158),
            .in2(_gnd_net_),
            .in3(N__35043),
            .lcout(\b2v_inst6.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_5_LC_12_3_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_5_LC_12_3_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_5_LC_12_3_0 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst6.count_5_LC_12_3_0  (
            .in0(N__34095),
            .in1(N__36124),
            .in2(N__36788),
            .in3(N__34126),
            .lcout(\b2v_inst6.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36663),
            .ce(N__35059),
            .sr(N__36114));
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIKJCQ2_LC_12_3_1 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIKJCQ2_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_8_c_RNIKJCQ2_LC_12_3_1 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_8_c_RNIKJCQ2_LC_12_3_1  (
            .in0(N__34059),
            .in1(N__36773),
            .in2(N__34078),
            .in3(N__36083),
            .lcout(\b2v_inst6.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIP83V8_5_LC_12_3_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIP83V8_5_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIP83V8_5_LC_12_3_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst6.count_RNIP83V8_5_LC_12_3_2  (
            .in0(N__34132),
            .in1(N__35041),
            .in2(_gnd_net_),
            .in3(N__34111),
            .lcout(\b2v_inst6.countZ0Z_5 ),
            .ltout(\b2v_inst6.countZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIGB8Q2_LC_12_3_3 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIGB8Q2_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_4_c_RNIGB8Q2_LC_12_3_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_4_c_RNIGB8Q2_LC_12_3_3  (
            .in0(N__34125),
            .in1(N__36772),
            .in2(N__34114),
            .in3(N__36082),
            .lcout(\b2v_inst6.count_rst_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI1L7V8_9_LC_12_3_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI1L7V8_9_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI1L7V8_9_LC_12_3_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst6.count_RNI1L7V8_9_LC_12_3_4  (
            .in0(N__34051),
            .in1(N__35042),
            .in2(_gnd_net_),
            .in3(N__34105),
            .lcout(\b2v_inst6.countZ0Z_9 ),
            .ltout(\b2v_inst6.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_5_LC_12_3_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_5_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_5_LC_12_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNI_5_LC_12_3_5  (
            .in0(N__34410),
            .in1(N__34331),
            .in2(N__34099),
            .in3(N__34094),
            .lcout(\b2v_inst6.count_1_i_a3_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_9_LC_12_3_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_9_LC_12_3_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_9_LC_12_3_6 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \b2v_inst6.count_9_LC_12_3_6  (
            .in0(N__36084),
            .in1(N__34074),
            .in2(N__36789),
            .in3(N__34060),
            .lcout(\b2v_inst6.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36663),
            .ce(N__35059),
            .sr(N__36114));
    defparam \b2v_inst6.count_7_LC_12_3_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_7_LC_12_3_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_7_LC_12_3_7 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst6.count_7_LC_12_3_7  (
            .in0(N__34411),
            .in1(N__36774),
            .in2(N__36130),
            .in3(N__34438),
            .lcout(\b2v_inst6.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36663),
            .ce(N__35059),
            .sr(N__36114));
    defparam \b2v_inst6.count_12_LC_12_4_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_12_LC_12_4_0 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_12_LC_12_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \b2v_inst6.count_12_LC_12_4_0  (
            .in0(N__34261),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36661),
            .ce(N__35053),
            .sr(N__36118));
    defparam \b2v_inst6.count_RNIA0P09_10_LC_12_4_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIA0P09_10_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIA0P09_10_LC_12_4_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \b2v_inst6.count_RNIA0P09_10_LC_12_4_1  (
            .in0(N__34444),
            .in1(N__35020),
            .in2(_gnd_net_),
            .in3(N__34182),
            .lcout(\b2v_inst6.countZ0Z_10 ),
            .ltout(\b2v_inst6.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_3_LC_12_4_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_3_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_3_LC_12_4_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \b2v_inst6.count_RNI_3_LC_12_4_2  (
            .in0(N__34245),
            .in1(N__34223),
            .in2(N__34270),
            .in3(N__34536),
            .lcout(\b2v_inst6.count_1_i_a3_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNILA289_12_LC_12_4_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNILA289_12_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNILA289_12_LC_12_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNILA289_12_LC_12_4_3  (
            .in0(N__34267),
            .in1(N__34260),
            .in2(_gnd_net_),
            .in3(N__35021),
            .lcout(\b2v_inst6.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIF97Q2_LC_12_4_4 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIF97Q2_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_3_c_RNIF97Q2_LC_12_4_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_3_c_RNIF97Q2_LC_12_4_4  (
            .in0(N__34203),
            .in1(N__36770),
            .in2(N__34228),
            .in3(N__36031),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIN52V8_4_LC_12_4_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIN52V8_4_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIN52V8_4_LC_12_4_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNIN52V8_4_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(N__34189),
            .in2(N__34231),
            .in3(N__35019),
            .lcout(\b2v_inst6.countZ0Z_4 ),
            .ltout(\b2v_inst6.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_4_LC_12_4_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_4_LC_12_4_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_4_LC_12_4_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.count_4_LC_12_4_6  (
            .in0(N__34204),
            .in1(N__36771),
            .in2(N__34192),
            .in3(N__36032),
            .lcout(\b2v_inst6.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36661),
            .ce(N__35053),
            .sr(N__36118));
    defparam \b2v_inst6.count_10_LC_12_4_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_10_LC_12_4_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_10_LC_12_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_10_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34183),
            .lcout(\b2v_inst6.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36661),
            .ce(N__35053),
            .sr(N__36118));
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIIFAQ2_LC_12_5_0 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIIFAQ2_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_6_c_RNIIFAQ2_LC_12_5_0 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_6_c_RNIIFAQ2_LC_12_5_0  (
            .in0(N__34408),
            .in1(N__36781),
            .in2(N__36076),
            .in3(N__34437),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNITE5V8_7_LC_12_5_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNITE5V8_7_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNITE5V8_7_LC_12_5_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNITE5V8_7_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__34423),
            .in2(N__34414),
            .in3(N__35022),
            .lcout(\b2v_inst6.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNIJHBQ2_LC_12_5_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNIJHBQ2_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_7_c_RNIJHBQ2_LC_12_5_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_7_c_RNIJHBQ2_LC_12_5_2  (
            .in0(N__34302),
            .in1(N__36782),
            .in2(N__34332),
            .in3(N__36037),
            .lcout(\b2v_inst6.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_15_LC_12_5_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_15_LC_12_5_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_15_LC_12_5_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \b2v_inst6.count_15_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__34386),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36656),
            .ce(N__35044),
            .sr(N__36036));
    defparam \b2v_inst6.count_RNIRJ589_15_LC_12_5_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRJ589_15_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRJ589_15_LC_12_5_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \b2v_inst6.count_RNIRJ589_15_LC_12_5_5  (
            .in0(N__34387),
            .in1(N__34375),
            .in2(_gnd_net_),
            .in3(N__35045),
            .lcout(\b2v_inst6.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_2_LC_12_5_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_2_LC_12_5_6 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_2_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \b2v_inst6.count_2_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34369),
            .lcout(\b2v_inst6.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36656),
            .ce(N__35044),
            .sr(N__36036));
    defparam \b2v_inst6.count_RNIVH6V8_8_LC_12_6_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIVH6V8_8_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIVH6V8_8_LC_12_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.count_RNIVH6V8_8_LC_12_6_1  (
            .in0(N__34285),
            .in1(N__34339),
            .in2(_gnd_net_),
            .in3(N__35017),
            .lcout(\b2v_inst6.countZ0Z_8 ),
            .ltout(\b2v_inst6.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_8_LC_12_6_2 .C_ON=1'b0;
    defparam \b2v_inst6.count_8_LC_12_6_2 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_8_LC_12_6_2 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.count_8_LC_12_6_2  (
            .in0(N__36030),
            .in1(N__36761),
            .in2(N__34306),
            .in3(N__34303),
            .lcout(\b2v_inst6.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36649),
            .ce(N__35018),
            .sr(N__36119));
    defparam \b2v_inst6.count_11_LC_12_6_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_11_LC_12_6_4 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_11_LC_12_6_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \b2v_inst6.count_11_LC_12_6_4  (
            .in0(N__36029),
            .in1(N__36760),
            .in2(N__34492),
            .in3(N__34624),
            .lcout(\b2v_inst6.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36649),
            .ce(N__35018),
            .sr(N__36119));
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIE76Q2_LC_12_6_5 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIE76Q2_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_2_c_RNIE76Q2_LC_12_6_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.un2_count_1_cry_2_c_RNIE76Q2_LC_12_6_5  (
            .in0(N__34512),
            .in1(N__36758),
            .in2(N__34537),
            .in3(N__36028),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIL21V8_3_LC_12_6_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIL21V8_3_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIL21V8_3_LC_12_6_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \b2v_inst6.count_RNIL21V8_3_LC_12_6_6  (
            .in0(N__35016),
            .in1(_gnd_net_),
            .in2(N__34540),
            .in3(N__34498),
            .lcout(\b2v_inst6.countZ0Z_3 ),
            .ltout(\b2v_inst6.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_3_LC_12_6_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_3_LC_12_6_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_3_LC_12_6_7 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \b2v_inst6.count_3_LC_12_6_7  (
            .in0(N__34513),
            .in1(N__36759),
            .in2(N__34501),
            .in3(N__36120),
            .lcout(\b2v_inst6.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36649),
            .ce(N__35018),
            .sr(N__36119));
    defparam \b2v_inst6.count_RNIM2CM2_0_LC_12_7_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIM2CM2_0_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIM2CM2_0_LC_12_7_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \b2v_inst6.count_RNIM2CM2_0_LC_12_7_0  (
            .in0(N__34564),
            .in1(_gnd_net_),
            .in2(N__34899),
            .in3(N__36039),
            .lcout(\b2v_inst6.count_RNIM2CM2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_0_LC_12_7_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_0_LC_12_7_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \b2v_inst6.count_RNI_0_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(N__34563),
            .in2(_gnd_net_),
            .in3(N__34892),
            .lcout(\b2v_inst6.N_394 ),
            .ltout(\b2v_inst6.N_394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNITRL13_LC_12_7_2 .C_ON=1'b0;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNITRL13_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.un2_count_1_cry_10_c_RNITRL13_LC_12_7_2 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \b2v_inst6.un2_count_1_cry_10_c_RNITRL13_LC_12_7_2  (
            .in0(N__34488),
            .in1(N__34625),
            .in2(N__34471),
            .in3(N__36038),
            .lcout(),
            .ltout(\b2v_inst6.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIJ7189_11_LC_12_7_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIJ7189_11_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIJ7189_11_LC_12_7_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \b2v_inst6.count_RNIJ7189_11_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(N__34468),
            .in2(N__34462),
            .in3(N__35023),
            .lcout(\b2v_inst6.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRR6R8_0_1_LC_12_8_0 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRR6R8_0_1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRR6R8_0_1_LC_12_8_0 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst6.count_RNIRR6R8_0_1_LC_12_8_0  (
            .in0(N__34675),
            .in1(N__34662),
            .in2(N__34995),
            .in3(N__36025),
            .lcout(\b2v_inst6.un2_count_1_axb_1 ),
            .ltout(\b2v_inst6.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNI_1_LC_12_8_1 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNI_1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNI_1_LC_12_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst6.count_RNI_1_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34768),
            .in3(N__34882),
            .lcout(\b2v_inst6.count_RNI_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_8_2 .C_ON=1'b0;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst5.un8_rsmrst_pwrgd_4_LC_12_8_2  (
            .in0(N__34765),
            .in1(N__34753),
            .in2(N__34738),
            .in3(N__34729),
            .lcout(N_1661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_1_LC_12_8_3 .C_ON=1'b0;
    defparam \b2v_inst6.count_1_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_1_LC_12_8_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \b2v_inst6.count_1_LC_12_8_3  (
            .in0(N__36027),
            .in1(_gnd_net_),
            .in2(N__34666),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36634),
            .ce(N__35046),
            .sr(N__36128));
    defparam \b2v_inst6.count_RNIRR6R8_1_LC_12_8_4 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRR6R8_1_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRR6R8_1_LC_12_8_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \b2v_inst6.count_RNIRR6R8_1_LC_12_8_4  (
            .in0(N__34674),
            .in1(N__34661),
            .in2(N__35057),
            .in3(N__36024),
            .lcout(),
            .ltout(\b2v_inst6.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRR6R8_2_1_LC_12_8_5 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRR6R8_2_1_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRR6R8_2_1_LC_12_8_5 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \b2v_inst6.count_RNIRR6R8_2_1_LC_12_8_5  (
            .in0(N__34644),
            .in1(_gnd_net_),
            .in2(N__34630),
            .in3(N__34627),
            .lcout(),
            .ltout(\b2v_inst6.count_1_i_a3_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIRR6R8_3_1_LC_12_8_6 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIRR6R8_3_1_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIRR6R8_3_1_LC_12_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \b2v_inst6.count_RNIRR6R8_3_1_LC_12_8_6  (
            .in0(N__34600),
            .in1(N__34588),
            .in2(N__34579),
            .in3(N__34576),
            .lcout(\b2v_inst6.N_389 ),
            .ltout(\b2v_inst6.N_389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_0_LC_12_8_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_0_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \b2v_inst6.count_0_LC_12_8_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \b2v_inst6.count_0_LC_12_8_7  (
            .in0(N__36026),
            .in1(_gnd_net_),
            .in2(N__34555),
            .in3(N__34883),
            .lcout(\b2v_inst6.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36634),
            .ce(N__35046),
            .sr(N__36128));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_12_9_1 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_12_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35575),
            .lcout(\b2v_inst11.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_12_9_2 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_12_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35204),
            .lcout(\b2v_inst11.mult1_un96_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_12_9_4 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_12_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34863),
            .lcout(\b2v_inst11.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_9_5 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36232),
            .lcout(\b2v_inst11.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI87PU5_0_LC_12_9_6 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI87PU5_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI87PU5_0_LC_12_9_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \b2v_inst6.curr_state_RNI87PU5_0_LC_12_9_6  (
            .in0(N__36699),
            .in1(N__36400),
            .in2(_gnd_net_),
            .in3(N__36023),
            .lcout(\b2v_inst6.count_en ),
            .ltout(\b2v_inst6.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.count_RNIQQ6R8_0_LC_12_9_7 .C_ON=1'b0;
    defparam \b2v_inst6.count_RNIQQ6R8_0_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.count_RNIQQ6R8_0_LC_12_9_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \b2v_inst6.count_RNIQQ6R8_0_LC_12_9_7  (
            .in0(N__34921),
            .in1(_gnd_net_),
            .in2(N__34909),
            .in3(N__34906),
            .lcout(\b2v_inst6.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_12_10_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__34864),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_12_10_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_12_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__34843),
            .in2(N__35154),
            .in3(N__34822),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_12_10_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_12_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__35150),
            .in2(N__34819),
            .in3(N__34798),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_12_10_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_12_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__35176),
            .in2(N__34795),
            .in3(N__34771),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_12_10_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_12_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__35275),
            .in2(N__35182),
            .in3(N__35257),
            .lcout(\b2v_inst11.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_12_10_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_12_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_12_10_5  (
            .in0(N__35203),
            .in1(N__35254),
            .in2(N__35155),
            .in3(N__35233),
            .lcout(\b2v_inst11.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un96_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_12_10_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_12_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35230),
            .in3(N__35221),
            .lcout(\b2v_inst11.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_12_10_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_12_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35175),
            .lcout(\b2v_inst11.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_11_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__35137),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_11_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__35116),
            .in2(N__35544),
            .in3(N__35101),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_11_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__35540),
            .in2(N__35314),
            .in3(N__35092),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_11_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__35302),
            .in2(N__35574),
            .in3(N__35080),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_11_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__35570),
            .in2(N__35293),
            .in3(N__35401),
            .lcout(\b2v_inst11.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_11_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_11_5  (
            .in0(N__35377),
            .in1(N__35281),
            .in2(N__35545),
            .in3(N__35389),
            .lcout(\b2v_inst11.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un82_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_11_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35590),
            .in3(N__35386),
            .lcout(\b2v_inst11.mult1_un82_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un82_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_12_11_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_12_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35359),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_12_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__35338),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_12_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__35320),
            .in2(N__35607),
            .in3(N__35305),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_12_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__35603),
            .in2(N__35497),
            .in3(N__35296),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_12_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__35476),
            .in2(N__36231),
            .in3(N__35284),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_12_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__36226),
            .in2(N__35461),
            .in3(N__35611),
            .lcout(\b2v_inst11.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_12_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_12_5  (
            .in0(N__35566),
            .in1(N__35416),
            .in2(N__35608),
            .in3(N__35581),
            .lcout(\b2v_inst11.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un75_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_12_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36256),
            .in3(N__35578),
            .lcout(\b2v_inst11.mult1_un75_sum_s_8 ),
            .ltout(\b2v_inst11.mult1_un75_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_12_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35548),
            .in3(_gnd_net_),
            .lcout(\b2v_inst11.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_13_0 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__35526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_13_1 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__35503),
            .in2(N__36273),
            .in3(N__35488),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_2 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_13_2 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__36269),
            .in2(N__35485),
            .in3(N__35470),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_3 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_13_3 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__35467),
            .in2(N__35449),
            .in3(N__35452),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_4 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_13_4 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__35447),
            .in2(N__35425),
            .in3(N__36286),
            .lcout(\b2v_inst11.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_5 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_13_5 .C_ON=1'b1;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_13_5  (
            .in0(N__36222),
            .in1(N__36283),
            .in2(N__36274),
            .in3(N__36247),
            .lcout(\b2v_inst11.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\b2v_inst11.mult1_un68_sum_cry_6 ),
            .carryout(\b2v_inst11.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_13_6 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36244),
            .in3(N__36235),
            .lcout(\b2v_inst11.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_12_13_7 .C_ON=1'b0;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_12_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst11.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36195),
            .lcout(\b2v_inst11.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI59E43_0_LC_12_14_0 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI59E43_0_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI59E43_0_LC_12_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \b2v_inst6.curr_state_RNI59E43_0_LC_12_14_0  (
            .in0(N__35944),
            .in1(N__35617),
            .in2(_gnd_net_),
            .in3(N__35898),
            .lcout(\b2v_inst6.curr_stateZ0Z_0 ),
            .ltout(\b2v_inst6.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNIM2CM2_0_LC_12_14_1 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNIM2CM2_0_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNIM2CM2_0_LC_12_14_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \b2v_inst6.curr_state_RNIM2CM2_0_LC_12_14_1  (
            .in0(N__35899),
            .in1(N__36146),
            .in2(N__36133),
            .in3(N__36820),
            .lcout(\b2v_inst6.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_0_LC_12_14_2 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_0_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_0_LC_12_14_2 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \b2v_inst6.curr_state_0_LC_12_14_2  (
            .in0(N__36802),
            .in1(N__35631),
            .in2(N__36790),
            .in3(N__35655),
            .lcout(\b2v_inst6.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36660),
            .ce(N__36366),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI6AE43_1_LC_12_14_3 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI6AE43_1_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI6AE43_1_LC_12_14_3 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \b2v_inst6.curr_state_RNI6AE43_1_LC_12_14_3  (
            .in0(N__35900),
            .in1(N__36670),
            .in2(N__36700),
            .in3(N__36706),
            .lcout(\b2v_inst6.curr_stateZ0Z_1 ),
            .ltout(\b2v_inst6.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_12_14_4 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m4_0_LC_12_14_4 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m4_0_LC_12_14_4  (
            .in0(N__36787),
            .in1(N__35656),
            .in2(N__35635),
            .in3(N__35630),
            .lcout(\b2v_inst6.curr_state_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_RNI_1_LC_12_14_5 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_RNI_1_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_RNI_1_LC_12_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \b2v_inst6.curr_state_RNI_1_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36800),
            .lcout(\b2v_inst6.N_2937_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_12_14_6 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_12_14_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \b2v_inst6.curr_state_7_1_0__m6_i_a3_LC_12_14_6  (
            .in0(N__36801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36783),
            .lcout(\b2v_inst6.m6_i_a3 ),
            .ltout(\b2v_inst6.m6_i_a3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b2v_inst6.curr_state_1_LC_12_14_7 .C_ON=1'b0;
    defparam \b2v_inst6.curr_state_1_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \b2v_inst6.curr_state_1_LC_12_14_7 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \b2v_inst6.curr_state_1_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__36692),
            .in2(N__36673),
            .in3(_gnd_net_),
            .lcout(\b2v_inst6.curr_state_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36660),
            .ce(N__36366),
            .sr(_gnd_net_));
endmodule // TOP
